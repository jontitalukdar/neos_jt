module sha1(clk_i, rst_i, text_i, text_o, cmd_i, cmd_w_i, cmd_o, d_out_1, q_in_1, qn_in_1, d_out_2, q_in_2, qn_in_2, d_out_3, q_in_3, qn_in_3, d_out_4, q_in_4, qn_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, q_in_7, d_out_8, q_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, qn_in_11, d_out_12, q_in_12, d_out_13, q_in_13, d_out_14, q_in_14, d_out_15, q_in_15, d_out_16, q_in_16, qn_in_16, d_out_17, q_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, q_in_20, d_out_21, q_in_21, d_out_22, q_in_22, d_out_23, q_in_23, d_out_24, q_in_24, d_out_25, q_in_25, d_out_26, q_in_26, d_out_27, q_in_27, qn_in_27, d_out_28, q_in_28, d_out_29, q_in_29, d_out_30, q_in_30, d_out_31, q_in_31, d_out_32, q_in_32, qn_in_32, d_out_33, q_in_33, d_out_34, q_in_34, d_out_35, q_in_35, d_out_36, q_in_36, d_out_37, q_in_37, d_out_38, q_in_38, d_out_39, q_in_39, d_out_40, q_in_40, d_out_41, q_in_41, d_out_42, q_in_42, d_out_43, q_in_43, qn_in_43, d_out_44, q_in_44, d_out_45, q_in_45, d_out_46, q_in_46, d_out_47, q_in_47, d_out_48, q_in_48, qn_in_48, d_out_49, q_in_49, d_out_50, q_in_50, d_out_51, q_in_51, d_out_52, q_in_52, d_out_53, q_in_53, d_out_54, q_in_54, d_out_55, q_in_55, d_out_56, q_in_56, d_out_57, q_in_57, d_out_58, q_in_58, d_out_59, q_in_59, qn_in_59, d_out_60, q_in_60, d_out_61, q_in_61, d_out_62, q_in_62, d_out_63, q_in_63, d_out_64, q_in_64, qn_in_64, d_out_65, q_in_65, d_out_66, q_in_66, d_out_67, q_in_67, d_out_68, q_in_68, d_out_69, q_in_69, d_out_70, q_in_70, d_out_71, q_in_71, d_out_72, q_in_72, d_out_73, q_in_73, d_out_74, q_in_74, d_out_75, q_in_75, qn_in_75, d_out_76, q_in_76, d_out_77, q_in_77, d_out_78, q_in_78, d_out_79, q_in_79, d_out_80, q_in_80, qn_in_80, d_out_81, q_in_81, d_out_82, q_in_82, d_out_83, q_in_83, d_out_84, q_in_84, d_out_85, q_in_85, d_out_86, q_in_86, d_out_87, q_in_87, d_out_88, q_in_88, d_out_89, q_in_89, d_out_90, q_in_90, d_out_91, q_in_91, qn_in_91, d_out_92, q_in_92, d_out_93, q_in_93, d_out_94, q_in_94, d_out_95, q_in_95, d_out_96, q_in_96, qn_in_96, d_out_97, q_in_97, d_out_98, q_in_98, d_out_99, q_in_99, d_out_100, q_in_100, d_out_101, q_in_101, d_out_102, q_in_102, d_out_103, q_in_103, d_out_104, q_in_104, d_out_105, q_in_105, d_out_106, q_in_106, d_out_107, q_in_107, qn_in_107, d_out_108, q_in_108, d_out_109, q_in_109, d_out_110, q_in_110, d_out_111, q_in_111, d_out_112, q_in_112, qn_in_112, d_out_113, q_in_113, d_out_114, q_in_114, d_out_115, q_in_115, d_out_116, q_in_116, d_out_117, q_in_117, d_out_118, q_in_118, d_out_119, q_in_119, d_out_120, q_in_120, d_out_121, q_in_121, d_out_122, q_in_122, d_out_123, q_in_123, qn_in_123, d_out_124, q_in_124, d_out_125, q_in_125, d_out_126, q_in_126, d_out_127, q_in_127, d_out_128, q_in_128, qn_in_128, d_out_129, q_in_129, d_out_130, q_in_130, d_out_131, q_in_131, d_out_132, q_in_132, d_out_133, q_in_133, d_out_134, q_in_134, d_out_135, q_in_135, d_out_136, q_in_136, d_out_137, q_in_137, d_out_138, q_in_138, d_out_139, q_in_139, qn_in_139, d_out_140, q_in_140, d_out_141, q_in_141, d_out_142, q_in_142, d_out_143, q_in_143, d_out_144, q_in_144, qn_in_144, d_out_145, q_in_145, d_out_146, q_in_146, d_out_147, q_in_147, d_out_148, q_in_148, d_out_149, q_in_149, d_out_150, q_in_150, d_out_151, q_in_151, d_out_152, q_in_152, d_out_153, q_in_153, d_out_154, q_in_154, d_out_155, q_in_155, qn_in_155, d_out_156, q_in_156, d_out_157, q_in_157, d_out_158, q_in_158, d_out_159, q_in_159, d_out_160, q_in_160, qn_in_160, d_out_161, q_in_161, d_out_162, q_in_162, d_out_163, q_in_163, d_out_164, q_in_164, d_out_165, q_in_165, d_out_166, q_in_166, d_out_167, q_in_167, d_out_168, q_in_168, d_out_169, q_in_169, d_out_170, q_in_170, d_out_171, q_in_171, qn_in_171, d_out_172, q_in_172, d_out_173, q_in_173, d_out_174, q_in_174, d_out_175, q_in_175, d_out_176, q_in_176, qn_in_176, d_out_177, q_in_177, d_out_178, q_in_178, d_out_179, q_in_179, d_out_180, q_in_180, d_out_181, q_in_181, d_out_182, q_in_182, d_out_183, q_in_183, d_out_184, q_in_184, d_out_185, q_in_185, d_out_186, q_in_186, d_out_187, q_in_187, qn_in_187, d_out_188, q_in_188, d_out_189, q_in_189, d_out_190, q_in_190, d_out_191, q_in_191, d_out_192, q_in_192, qn_in_192, d_out_193, q_in_193, d_out_194, q_in_194, d_out_195, q_in_195, d_out_196, q_in_196, d_out_197, q_in_197, d_out_198, q_in_198, d_out_199, q_in_199, d_out_200, q_in_200, d_out_201, q_in_201, d_out_202, q_in_202, d_out_203, q_in_203, qn_in_203, d_out_204, q_in_204, d_out_205, q_in_205, d_out_206, q_in_206, d_out_207, q_in_207, d_out_208, q_in_208, qn_in_208, d_out_209, q_in_209, d_out_210, q_in_210, d_out_211, q_in_211, d_out_212, q_in_212, d_out_213, q_in_213, d_out_214, q_in_214, d_out_215, q_in_215, d_out_216, q_in_216, d_out_217, q_in_217, d_out_218, q_in_218, d_out_219, q_in_219, qn_in_219, d_out_220, q_in_220, d_out_221, q_in_221, d_out_222, q_in_222, d_out_223, q_in_223, d_out_224, q_in_224, qn_in_224, d_out_225, q_in_225, d_out_226, q_in_226, d_out_227, q_in_227, d_out_228, q_in_228, d_out_229, q_in_229, d_out_230, q_in_230, d_out_231, q_in_231, d_out_232, q_in_232, d_out_233, q_in_233, d_out_234, q_in_234, d_out_235, q_in_235, qn_in_235, d_out_236, q_in_236, d_out_237, q_in_237, d_out_238, q_in_238, d_out_239, q_in_239, d_out_240, q_in_240, qn_in_240, d_out_241, q_in_241, d_out_242, q_in_242, d_out_243, q_in_243, d_out_244, q_in_244, d_out_245, q_in_245, d_out_246, q_in_246, d_out_247, q_in_247, d_out_248, q_in_248, d_out_249, q_in_249, d_out_250, q_in_250, d_out_251, q_in_251, qn_in_251, d_out_252, q_in_252, d_out_253, q_in_253, d_out_254, q_in_254, d_out_255, q_in_255, d_out_256, q_in_256, qn_in_256, d_out_257, q_in_257, d_out_258, q_in_258, d_out_259, q_in_259, d_out_260, q_in_260, d_out_261, q_in_261, d_out_262, q_in_262, d_out_263, q_in_263, d_out_264, q_in_264, d_out_265, q_in_265, d_out_266, q_in_266, d_out_267, q_in_267, qn_in_267, d_out_268, q_in_268, d_out_269, q_in_269, d_out_270, q_in_270, d_out_271, q_in_271, d_out_272, q_in_272, qn_in_272, d_out_273, q_in_273, d_out_274, q_in_274, d_out_275, q_in_275, d_out_276, q_in_276, d_out_277, q_in_277, d_out_278, q_in_278, d_out_279, q_in_279, d_out_280, q_in_280, d_out_281, q_in_281, d_out_282, q_in_282, d_out_283, q_in_283, qn_in_283, d_out_284, q_in_284, d_out_285, q_in_285, d_out_286, q_in_286, d_out_287, q_in_287, d_out_288, q_in_288, qn_in_288, d_out_289, q_in_289, d_out_290, q_in_290, d_out_291, q_in_291, d_out_292, q_in_292, d_out_293, q_in_293, d_out_294, q_in_294, d_out_295, q_in_295, d_out_296, q_in_296, d_out_297, q_in_297, d_out_298, q_in_298, d_out_299, q_in_299, qn_in_299, d_out_300, q_in_300, d_out_301, q_in_301, d_out_302, q_in_302, d_out_303, q_in_303, d_out_304, q_in_304, qn_in_304, d_out_305, q_in_305, d_out_306, q_in_306, d_out_307, q_in_307, d_out_308, q_in_308, d_out_309, q_in_309, d_out_310, q_in_310, d_out_311, q_in_311, d_out_312, q_in_312, d_out_313, q_in_313, d_out_314, q_in_314, d_out_315, q_in_315, qn_in_315, d_out_316, q_in_316, d_out_317, q_in_317, d_out_318, q_in_318, d_out_319, q_in_319, d_out_320, q_in_320, qn_in_320, d_out_321, q_in_321, d_out_322, q_in_322, d_out_323, q_in_323, d_out_324, q_in_324, d_out_325, q_in_325, d_out_326, q_in_326, d_out_327, q_in_327, d_out_328, q_in_328, d_out_329, q_in_329, d_out_330, q_in_330, d_out_331, q_in_331, qn_in_331, d_out_332, q_in_332, d_out_333, q_in_333, d_out_334, q_in_334, d_out_335, q_in_335, d_out_336, q_in_336, qn_in_336, d_out_337, q_in_337, d_out_338, q_in_338, d_out_339, q_in_339, d_out_340, q_in_340, d_out_341, q_in_341, d_out_342, q_in_342, d_out_343, q_in_343, d_out_344, q_in_344, d_out_345, q_in_345, d_out_346, q_in_346, d_out_347, q_in_347, qn_in_347, d_out_348, q_in_348, d_out_349, q_in_349, d_out_350, q_in_350, d_out_351, q_in_351, d_out_352, q_in_352, qn_in_352, d_out_353, q_in_353, d_out_354, q_in_354, d_out_355, q_in_355, d_out_356, q_in_356, d_out_357, q_in_357, d_out_358, q_in_358, d_out_359, q_in_359, d_out_360, q_in_360, d_out_361, q_in_361, d_out_362, q_in_362, d_out_363, q_in_363, qn_in_363, d_out_364, q_in_364, d_out_365, q_in_365, d_out_366, q_in_366, d_out_367, q_in_367, d_out_368, q_in_368, qn_in_368, d_out_369, q_in_369, d_out_370, q_in_370, d_out_371, q_in_371, d_out_372, q_in_372, d_out_373, q_in_373, d_out_374, q_in_374, d_out_375, q_in_375, d_out_376, q_in_376, d_out_377, q_in_377, d_out_378, q_in_378, d_out_379, q_in_379, qn_in_379, d_out_380, q_in_380, d_out_381, q_in_381, d_out_382, q_in_382, d_out_383, q_in_383, d_out_384, q_in_384, qn_in_384, d_out_385, q_in_385, d_out_386, q_in_386, d_out_387, q_in_387, d_out_388, q_in_388, d_out_389, q_in_389, d_out_390, q_in_390, d_out_391, q_in_391, d_out_392, q_in_392, d_out_393, q_in_393, d_out_394, q_in_394, d_out_395, q_in_395, qn_in_395, d_out_396, q_in_396, d_out_397, q_in_397, d_out_398, q_in_398, d_out_399, q_in_399, d_out_400, q_in_400, qn_in_400, d_out_401, q_in_401, d_out_402, q_in_402, d_out_403, q_in_403, d_out_404, q_in_404, d_out_405, q_in_405, d_out_406, q_in_406, d_out_407, q_in_407, d_out_408, q_in_408, d_out_409, q_in_409, d_out_410, q_in_410, d_out_411, q_in_411, qn_in_411, d_out_412, q_in_412, d_out_413, q_in_413, d_out_414, q_in_414, d_out_415, q_in_415, d_out_416, q_in_416, qn_in_416, d_out_417, q_in_417, d_out_418, q_in_418, d_out_419, q_in_419, d_out_420, q_in_420, d_out_421, q_in_421, d_out_422, q_in_422, d_out_423, q_in_423, d_out_424, q_in_424, d_out_425, q_in_425, d_out_426, q_in_426, d_out_427, q_in_427, qn_in_427, d_out_428, q_in_428, d_out_429, q_in_429, d_out_430, q_in_430, d_out_431, q_in_431, d_out_432, q_in_432, qn_in_432, d_out_433, q_in_433, d_out_434, q_in_434, d_out_435, q_in_435, d_out_436, q_in_436, d_out_437, q_in_437, d_out_438, q_in_438, d_out_439, q_in_439, d_out_440, q_in_440, d_out_441, q_in_441, d_out_442, q_in_442, d_out_443, q_in_443, qn_in_443, d_out_444, q_in_444, d_out_445, q_in_445, d_out_446, q_in_446, d_out_447, q_in_447, d_out_448, q_in_448, qn_in_448, d_out_449, q_in_449, d_out_450, q_in_450, d_out_451, q_in_451, d_out_452, q_in_452, d_out_453, q_in_453, d_out_454, q_in_454, d_out_455, q_in_455, d_out_456, q_in_456, d_out_457, q_in_457, d_out_458, q_in_458, d_out_459, q_in_459, qn_in_459, d_out_460, q_in_460, d_out_461, q_in_461, d_out_462, q_in_462, d_out_463, q_in_463, d_out_464, q_in_464, qn_in_464, d_out_465, q_in_465, d_out_466, q_in_466, d_out_467, q_in_467, d_out_468, q_in_468, d_out_469, q_in_469, d_out_470, q_in_470, d_out_471, q_in_471, d_out_472, q_in_472, d_out_473, q_in_473, d_out_474, q_in_474, d_out_475, q_in_475, qn_in_475, d_out_476, q_in_476, d_out_477, q_in_477, d_out_478, q_in_478, d_out_479, q_in_479, d_out_480, q_in_480, qn_in_480, d_out_481, q_in_481, d_out_482, q_in_482, d_out_483, q_in_483, d_out_484, q_in_484, d_out_485, q_in_485, d_out_486, q_in_486, d_out_487, q_in_487, d_out_488, q_in_488, d_out_489, q_in_489, d_out_490, q_in_490, d_out_491, q_in_491, qn_in_491, d_out_492, q_in_492, d_out_493, q_in_493, d_out_494, q_in_494, d_out_495, q_in_495, d_out_496, q_in_496, qn_in_496, d_out_497, q_in_497, d_out_498, q_in_498, d_out_499, q_in_499, d_out_500, q_in_500, d_out_501, q_in_501, d_out_502, q_in_502, d_out_503, q_in_503, d_out_504, q_in_504, d_out_505, q_in_505, d_out_506, q_in_506, d_out_507, q_in_507, qn_in_507, d_out_508, q_in_508, d_out_509, q_in_509, d_out_510, q_in_510, d_out_511, q_in_511, d_out_512, q_in_512, qn_in_512, d_out_513, q_in_513, d_out_514, q_in_514, d_out_515, q_in_515, d_out_516, q_in_516, d_out_517, q_in_517, d_out_518, q_in_518, qn_in_518, d_out_519, q_in_519, qn_in_519, d_out_520, q_in_520, d_out_521, q_in_521, qn_in_521, d_out_522, q_in_522, d_out_523, q_in_523, qn_in_523, d_out_524, q_in_524, d_out_525, q_in_525, qn_in_525, d_out_526, q_in_526, d_out_527, q_in_527, qn_in_527, d_out_528, q_in_528, d_out_529, q_in_529, qn_in_529, d_out_530, q_in_530, d_out_531, q_in_531, qn_in_531, d_out_532, q_in_532, d_out_533, q_in_533, qn_in_533, d_out_534, q_in_534, d_out_535, q_in_535, d_out_536, q_in_536, qn_in_536, d_out_537, q_in_537, d_out_538, q_in_538, d_out_539, q_in_539, d_out_540, q_in_540, d_out_541, q_in_541, d_out_542, q_in_542, d_out_543, q_in_543, d_out_544, q_in_544, d_out_545, q_in_545, d_out_546, q_in_546, d_out_547, q_in_547, qn_in_547, d_out_548, q_in_548, d_out_549, q_in_549, d_out_550, q_in_550, d_out_551, q_in_551, d_out_552, q_in_552, d_out_553, q_in_553, d_out_554, q_in_554, d_out_555, q_in_555, d_out_556, q_in_556, d_out_557, q_in_557, d_out_558, q_in_558, qn_in_558, d_out_559, q_in_559, d_out_560, q_in_560, qn_in_560, d_out_561, q_in_561, d_out_562, q_in_562, d_out_563, q_in_563, qn_in_563, d_out_564, q_in_564, d_out_565, q_in_565, d_out_566, q_in_566, qn_in_566, d_out_567, q_in_567, d_out_568, q_in_568, d_out_569, q_in_569, qn_in_569, d_out_570, q_in_570, d_out_571, q_in_571, qn_in_571, d_out_572, q_in_572, d_out_573, q_in_573, qn_in_573, d_out_574, q_in_574, d_out_575, q_in_575, qn_in_575, d_out_576, q_in_576, d_out_577, q_in_577, qn_in_577, d_out_578, q_in_578, d_out_579, q_in_579, qn_in_579, d_out_580, q_in_580, d_out_581, q_in_581, qn_in_581, d_out_582, q_in_582, d_out_583, q_in_583, qn_in_583, d_out_584, q_in_584, d_out_585, q_in_585, qn_in_585, d_out_586, q_in_586, d_out_587, q_in_587, qn_in_587, d_out_588, q_in_588, d_out_589, q_in_589, qn_in_589, d_out_590, q_in_590, d_out_591, q_in_591, qn_in_591, d_out_592, q_in_592, d_out_593, q_in_593, qn_in_593, d_out_594, q_in_594, d_out_595, q_in_595, d_out_596, q_in_596, qn_in_596, d_out_597, q_in_597, d_out_598, q_in_598, qn_in_598, d_out_599, q_in_599, d_out_600, q_in_600, qn_in_600, d_out_601, q_in_601, d_out_602, q_in_602, d_out_603, q_in_603, qn_in_603, d_out_604, q_in_604, d_out_605, q_in_605, qn_in_605, d_out_606, q_in_606, d_out_607, q_in_607, qn_in_607, d_out_608, q_in_608, d_out_609, q_in_609, qn_in_609, d_out_610, q_in_610, d_out_611, q_in_611, qn_in_611, d_out_612, q_in_612, d_out_613, q_in_613, qn_in_613, d_out_614, q_in_614, d_out_615, q_in_615, qn_in_615, d_out_616, q_in_616, d_out_617, q_in_617, qn_in_617, d_out_618, q_in_618, d_out_619, q_in_619, qn_in_619, d_out_620, q_in_620, d_out_621, q_in_621, qn_in_621, d_out_622, q_in_622, qn_in_622, d_out_623, q_in_623, qn_in_623, d_out_624, q_in_624, qn_in_624, d_out_625, q_in_625, d_out_626, q_in_626, qn_in_626, d_out_627, q_in_627, qn_in_627, d_out_628, q_in_628, d_out_629, q_in_629, qn_in_629, d_out_630, q_in_630, d_out_631, q_in_631, qn_in_631, d_out_632, q_in_632, qn_in_632, d_out_633, q_in_633, qn_in_633, d_out_634, q_in_634, d_out_635, q_in_635, qn_in_635, d_out_636, q_in_636, d_out_637, q_in_637, qn_in_637, d_out_638, q_in_638, d_out_639, q_in_639, qn_in_639, d_out_640, q_in_640, d_out_641, q_in_641, qn_in_641, d_out_642, q_in_642, d_out_643, q_in_643, qn_in_643, d_out_644, q_in_644, d_out_645, q_in_645, qn_in_645, d_out_646, q_in_646, d_out_647, q_in_647, qn_in_647, d_out_648, q_in_648, d_out_649, q_in_649, qn_in_649, d_out_650, q_in_650, d_out_651, q_in_651, qn_in_651, d_out_652, q_in_652, d_out_653, q_in_653, qn_in_653, d_out_654, q_in_654, d_out_655, q_in_655, qn_in_655, d_out_656, q_in_656, d_out_657, q_in_657, qn_in_657, d_out_658, q_in_658, d_out_659, q_in_659, qn_in_659, d_out_660, q_in_660, d_out_661, q_in_661, qn_in_661, d_out_662, q_in_662, d_out_663, q_in_663, qn_in_663, d_out_664, q_in_664, d_out_665, q_in_665, qn_in_665, d_out_666, q_in_666, d_out_667, q_in_667, qn_in_667, d_out_668, q_in_668, d_out_669, q_in_669, qn_in_669, d_out_670, q_in_670, d_out_671, q_in_671, d_out_672, q_in_672, qn_in_672, d_out_673, q_in_673, qn_in_673, d_out_674, q_in_674, d_out_675, q_in_675, d_out_676, q_in_676, qn_in_676, d_out_677, q_in_677, d_out_678, q_in_678, qn_in_678, d_out_679, q_in_679, qn_in_679, d_out_680, q_in_680, d_out_681, q_in_681, d_out_682, q_in_682, d_out_683, q_in_683, d_out_684, q_in_684, qn_in_684, d_out_685, q_in_685, d_out_686, q_in_686, d_out_687, q_in_687, d_out_688, q_in_688, d_out_689, q_in_689, d_out_690, q_in_690, d_out_691, q_in_691, d_out_692, q_in_692, d_out_693, q_in_693, d_out_694, q_in_694, d_out_695, q_in_695, d_out_696, q_in_696, d_out_697, q_in_697, d_out_698, q_in_698, d_out_699, q_in_699, d_out_700, q_in_700, qn_in_700, d_out_701, q_in_701, qn_in_701, d_out_702, q_in_702, d_out_703, q_in_703, d_out_704, q_in_704, d_out_705, q_in_705, d_out_706, q_in_706, d_out_707, q_in_707, d_out_708, q_in_708, d_out_709, q_in_709, d_out_710, q_in_710, d_out_711, q_in_711, d_out_712, q_in_712, d_out_713, q_in_713, d_out_714, q_in_714, d_out_715, q_in_715, d_out_716, q_in_716, d_out_717, q_in_717, d_out_718, q_in_718, qn_in_718, d_out_719, q_in_719, d_out_720, q_in_720, d_out_721, q_in_721, d_out_722, q_in_722, d_out_723, q_in_723, d_out_724, q_in_724, d_out_725, q_in_725, d_out_726, q_in_726, d_out_727, q_in_727, d_out_728, q_in_728, d_out_729, q_in_729, d_out_730, q_in_730, d_out_731, q_in_731, d_out_732, q_in_732, d_out_733, q_in_733, d_out_734, q_in_734, d_out_735, q_in_735, d_out_736, q_in_736, d_out_737, q_in_737, d_out_738, q_in_738, d_out_739, q_in_739, d_out_740, q_in_740, d_out_741, q_in_741, d_out_742, q_in_742, d_out_743, q_in_743, d_out_744, q_in_744, d_out_745, q_in_745, d_out_746, q_in_746, d_out_747, q_in_747, d_out_748, q_in_748, d_out_749, q_in_749, d_out_750, q_in_750, d_out_751, q_in_751, d_out_752, q_in_752, d_out_753, q_in_753, d_out_754, q_in_754, d_out_755, q_in_755, d_out_756, q_in_756, d_out_757, q_in_757, d_out_758, q_in_758, d_out_759, q_in_759, d_out_760, q_in_760, d_out_761, q_in_761, d_out_762, q_in_762, d_out_763, q_in_763, d_out_764, q_in_764, d_out_765, q_in_765, d_out_766, q_in_766, d_out_767, q_in_767, d_out_768, q_in_768, d_out_769, q_in_769, d_out_770, q_in_770, d_out_771, q_in_771, d_out_772, q_in_772, d_out_773, q_in_773, d_out_774, q_in_774, d_out_775, q_in_775, d_out_776, q_in_776, d_out_777, q_in_777, d_out_778, q_in_778, d_out_779, q_in_779, d_out_780, q_in_780, qn_in_780, d_out_781, q_in_781, qn_in_781, d_out_782, q_in_782, qn_in_782, d_out_783, q_in_783, qn_in_783, d_out_784, q_in_784, qn_in_784, d_out_785, q_in_785, qn_in_785, d_out_786, q_in_786, qn_in_786, d_out_787, q_in_787, qn_in_787, d_out_788, q_in_788, qn_in_788, d_out_789, q_in_789, qn_in_789, d_out_790, q_in_790, qn_in_790, d_out_791, q_in_791, qn_in_791, d_out_792, q_in_792, qn_in_792, d_out_793, q_in_793, qn_in_793, d_out_794, q_in_794, qn_in_794, d_out_795, q_in_795, qn_in_795, d_out_796, q_in_796, qn_in_796, d_out_797, q_in_797, qn_in_797, d_out_798, q_in_798, qn_in_798, d_out_799, q_in_799, qn_in_799, d_out_800, q_in_800, qn_in_800, d_out_801, q_in_801, qn_in_801, d_out_802, q_in_802, qn_in_802, d_out_803, q_in_803, qn_in_803, d_out_804, q_in_804, qn_in_804, d_out_805, q_in_805, qn_in_805, d_out_806, q_in_806, qn_in_806, d_out_807, q_in_807, qn_in_807, d_out_808, q_in_808, qn_in_808, d_out_809, q_in_809, qn_in_809, d_out_810, q_in_810, qn_in_810, d_out_811, q_in_811, qn_in_811, d_out_812, q_in_812, qn_in_812, d_out_813, q_in_813, qn_in_813, d_out_814, q_in_814, qn_in_814, d_out_815, q_in_815, qn_in_815, d_out_816, q_in_816, qn_in_816, d_out_817, q_in_817, qn_in_817, d_out_818, q_in_818, qn_in_818, d_out_819, q_in_819, qn_in_819, d_out_820, q_in_820, qn_in_820, d_out_821, q_in_821, qn_in_821, d_out_822, q_in_822, qn_in_822, d_out_823, q_in_823, qn_in_823, d_out_824, q_in_824, qn_in_824, d_out_825, q_in_825, qn_in_825, d_out_826, q_in_826, qn_in_826, d_out_827, q_in_827, qn_in_827, d_out_828, q_in_828, qn_in_828, d_out_829, q_in_829, d_out_830, q_in_830, d_out_831, q_in_831, d_out_832, q_in_832, d_out_833, q_in_833, d_out_834, q_in_834, d_out_835, q_in_835, d_out_836, q_in_836, qn_in_836, d_out_837, q_in_837, d_out_838, q_in_838, d_out_839, q_in_839, d_out_840, q_in_840, d_out_841, q_in_841, d_out_842, q_in_842, d_out_843, q_in_843, d_out_844, q_in_844, d_out_845, q_in_845, d_out_846, q_in_846, d_out_847, q_in_847, d_out_848, q_in_848, d_out_849, q_in_849, d_out_850, q_in_850, d_out_851, q_in_851, d_out_852, q_in_852, d_out_853, q_in_853, d_out_854, q_in_854, d_out_855, q_in_855, d_out_856, q_in_856, d_out_857, q_in_857, d_out_858, q_in_858, d_out_859, q_in_859, d_out_860, q_in_860, d_out_861, q_in_861, d_out_862, q_in_862, d_out_863, q_in_863, d_out_864, q_in_864, d_out_865, q_in_865, d_out_866, q_in_866, d_out_867, q_in_867, d_out_868, q_in_868, d_out_869, q_in_869, d_out_870, q_in_870, d_out_871, q_in_871, d_out_872, q_in_872, d_out_873, q_in_873, d_out_874, q_in_874, d_out_875, q_in_875, d_out_876, q_in_876, d_out_877, q_in_877, d_out_878, q_in_878, d_out_879, q_in_879, d_out_880, q_in_880, d_out_881, q_in_881, d_out_882, q_in_882, d_out_883, q_in_883, d_out_884, q_in_884, d_out_885, q_in_885, d_out_886, q_in_886, d_out_887, q_in_887, d_out_888, q_in_888, d_out_889, q_in_889, d_out_890, q_in_890, d_out_891, q_in_891, d_out_892, q_in_892, d_out_893, q_in_893, qn_in_893, d_out_894, q_in_894, qn_in_894, d_out_895, q_in_895, d_out_896, q_in_896, qn_in_896, d_out_897, q_in_897, qn_in_897, d_out_898, q_in_898, qn_in_898, d_out_899, q_in_899, qn_in_899, d_out_900, q_in_900, qn_in_900, d_out_901, q_in_901, qn_in_901, d_out_902, q_in_902, qn_in_902, d_out_903, q_in_903, qn_in_903, d_out_904, q_in_904, qn_in_904, d_out_905, q_in_905, qn_in_905, d_out_906, q_in_906, qn_in_906, d_out_907, q_in_907, qn_in_907, d_out_908, q_in_908, qn_in_908, d_out_909, q_in_909, qn_in_909, d_out_910, q_in_910, qn_in_910);
input qn_in_491;
input qn_in_836;
input qn_in_480;
input qn_in_560;
input qn_in_475;
input qn_in_464;
input qn_in_459;
input qn_in_818;
input qn_in_59;
input qn_in_448;
input qn_in_443;
input qn_in_432;
input qn_in_910;
input qn_in_427;
input qn_in_908;
input qn_in_907;
input qn_in_906;
input qn_in_905;
input qn_in_904;
input qn_in_903;
input qn_in_902;
input qn_in_901;
input qn_in_651;
input qn_in_899;
input qn_in_416;
input qn_in_897;
input qn_in_896;
input qn_in_894;
input qn_in_411;
input qn_in_400;
input qn_in_395;
input qn_in_384;
input qn_in_795;
input qn_in_379;
input qn_in_368;
input qn_in_363;
input qn_in_811;
input qn_in_624;
input qn_in_352;
input qn_in_347;
input qn_in_828;
input qn_in_827;
input qn_in_826;
input qn_in_825;
input qn_in_824;
input qn_in_823;
input qn_in_822;
input qn_in_821;
input qn_in_820;
input qn_in_819;
input qn_in_336;
input qn_in_817;
input qn_in_816;
input qn_in_815;
input qn_in_814;
input qn_in_331;
input qn_in_812;
input qn_in_635;
input qn_in_320;
input qn_in_315;
input qn_in_813;
input qn_in_304;
input qn_in_299;
input qn_in_810;
input qn_in_809;
input qn_in_808;
input qn_in_807;
input qn_in_806;
input qn_in_805;
input qn_in_804;
input qn_in_803;
input qn_in_802;
input qn_in_801;
input qn_in_288;
input qn_in_799;
input qn_in_798;
input qn_in_797;
input qn_in_796;
input qn_in_283;
input qn_in_794;
input qn_in_793;
input qn_in_792;
input qn_in_791;
input qn_in_790;
input qn_in_789;
input qn_in_788;
input qn_in_787;
input qn_in_786;
input qn_in_785;
input qn_in_272;
input qn_in_783;
input qn_in_782;
input qn_in_781;
input qn_in_780;
input qn_in_267;
input qn_in_672;
input qn_in_256;
input qn_in_251;
input qn_in_240;
input qn_in_898;
input qn_in_235;
input qn_in_619;
input qn_in_224;
input qn_in_219;
input qn_in_208;
input qn_in_718;
input qn_in_203;
input qn_in_192;
input qn_in_701;
input qn_in_700;
input qn_in_187;
input qn_in_176;
input qn_in_684;
input qn_in_171;
input qn_in_679;
input qn_in_678;
input qn_in_676;
input qn_in_523;
input qn_in_673;
input qn_in_160;
input qn_in_669;
input qn_in_155;
input qn_in_665;
input qn_in_663;
input qn_in_661;
input qn_in_893;
input qn_in_659;
input qn_in_657;
input qn_in_144;
input qn_in_655;
input qn_in_653;
input qn_in_139;
input qn_in_649;
input qn_in_647;
input qn_in_645;
input qn_in_643;
input qn_in_603;
input qn_in_641;
input qn_in_128;
input qn_in_639;
input qn_in_637;
input qn_in_123;
input qn_in_633;
input qn_in_632;
input qn_in_631;
input qn_in_629;
input qn_in_627;
input qn_in_626;
input qn_in_112;
input qn_in_623;
input qn_in_622;
input qn_in_621;
input qn_in_667;
input qn_in_107;
input qn_in_617;
input qn_in_615;
input qn_in_613;
input qn_in_800;
input qn_in_611;
input qn_in_909;
input qn_in_609;
input qn_in_96;
input qn_in_607;
input qn_in_605;
input qn_in_91;
input qn_in_600;
input qn_in_598;
input qn_in_596;
input qn_in_593;
input qn_in_80;
input qn_in_591;
input qn_in_589;
input qn_in_75;
input qn_in_585;
input qn_in_583;
input qn_in_581;
input qn_in_579;
input qn_in_577;
input qn_in_64;
input qn_in_575;
input qn_in_573;
input qn_in_571;
input qn_in_569;
input qn_in_566;
input qn_in_563;
input qn_in_48;
input qn_in_558;
input qn_in_900;
input qn_in_43;
input qn_in_784;
input qn_in_547;
input qn_in_587;
input qn_in_32;
input qn_in_27;
input qn_in_536;
input qn_in_533;
input qn_in_531;
input qn_in_529;
input qn_in_16;
input qn_in_527;
input qn_in_525;
input qn_in_11;
input qn_in_521;
input qn_in_519;
input qn_in_518;
input qn_in_4;
input qn_in_3;
input qn_in_2;
input qn_in_1;
input qn_in_512;
input qn_in_507;
input qn_in_496;
input q_in_910;
input q_in_909;
input q_in_908;
input q_in_907;
input q_in_906;
input q_in_905;
input q_in_904;
input q_in_903;
input q_in_902;
input q_in_901;
input q_in_900;
input q_in_899;
input q_in_898;
input q_in_897;
input q_in_896;
input q_in_895;
input q_in_894;
input q_in_893;
input q_in_892;
input q_in_891;
input q_in_890;
input q_in_889;
input q_in_888;
input q_in_887;
input q_in_886;
input q_in_885;
input q_in_884;
input q_in_883;
input q_in_882;
input q_in_881;
input q_in_880;
input q_in_879;
input q_in_878;
input q_in_877;
input q_in_876;
input q_in_875;
input q_in_874;
input q_in_873;
input q_in_872;
input q_in_871;
input q_in_870;
input q_in_869;
input q_in_868;
input q_in_867;
input q_in_866;
input q_in_865;
input q_in_864;
input q_in_863;
input q_in_862;
input q_in_861;
input q_in_860;
input q_in_859;
input q_in_858;
input q_in_857;
input q_in_856;
input q_in_855;
input q_in_854;
input q_in_853;
input q_in_852;
input q_in_851;
input q_in_850;
input q_in_849;
input q_in_848;
input q_in_847;
input q_in_846;
input q_in_845;
input q_in_844;
input q_in_843;
input q_in_842;
input q_in_841;
input q_in_840;
input q_in_839;
input q_in_838;
input q_in_837;
input q_in_836;
input q_in_835;
input q_in_834;
input q_in_833;
input q_in_832;
input q_in_831;
input q_in_830;
input q_in_829;
input q_in_828;
input q_in_827;
input q_in_826;
input q_in_825;
input q_in_824;
input q_in_823;
input q_in_822;
input q_in_821;
input q_in_820;
input q_in_819;
input q_in_818;
input q_in_817;
input q_in_816;
input q_in_815;
input q_in_814;
input q_in_813;
input q_in_812;
input q_in_811;
input q_in_810;
input q_in_809;
input q_in_808;
input q_in_807;
input q_in_806;
input q_in_805;
input q_in_804;
input q_in_803;
input q_in_802;
input q_in_801;
input q_in_800;
input q_in_799;
input q_in_798;
input q_in_797;
input q_in_796;
input q_in_795;
input q_in_794;
input q_in_793;
input q_in_792;
input q_in_791;
input q_in_790;
input q_in_789;
input q_in_788;
input q_in_787;
input q_in_786;
input q_in_785;
input q_in_784;
input q_in_783;
input q_in_782;
input q_in_781;
input q_in_780;
input q_in_779;
input q_in_778;
input q_in_777;
input q_in_776;
input q_in_775;
input q_in_774;
input q_in_773;
input q_in_772;
input q_in_771;
input q_in_770;
input q_in_769;
input q_in_768;
input q_in_767;
input q_in_766;
input q_in_765;
input q_in_764;
input q_in_763;
input q_in_762;
input q_in_761;
input q_in_760;
input q_in_759;
input q_in_758;
input q_in_757;
input q_in_756;
input q_in_755;
input q_in_754;
input q_in_753;
input q_in_752;
input q_in_751;
input q_in_750;
input q_in_749;
input q_in_748;
input q_in_747;
input q_in_746;
input q_in_745;
input q_in_744;
input q_in_743;
input q_in_742;
input q_in_741;
input q_in_740;
input q_in_739;
input q_in_738;
input q_in_737;
input q_in_736;
input q_in_735;
input q_in_734;
input q_in_733;
input q_in_732;
input q_in_731;
input q_in_730;
input q_in_729;
input q_in_728;
input q_in_727;
input q_in_726;
input q_in_725;
input q_in_724;
input q_in_723;
input q_in_722;
input q_in_721;
input q_in_720;
input q_in_719;
input q_in_718;
input q_in_717;
input q_in_716;
input q_in_715;
input q_in_714;
input q_in_713;
input q_in_712;
input q_in_711;
input q_in_710;
input q_in_709;
input q_in_708;
input q_in_707;
input q_in_706;
input q_in_705;
input q_in_704;
input q_in_703;
input q_in_702;
input q_in_701;
input q_in_700;
input q_in_699;
input q_in_698;
input q_in_697;
input q_in_696;
input q_in_695;
input q_in_694;
input q_in_693;
input q_in_692;
input q_in_691;
input q_in_690;
input q_in_689;
input q_in_688;
input q_in_687;
input q_in_686;
input q_in_685;
input q_in_684;
input q_in_683;
input q_in_682;
input q_in_681;
input q_in_680;
input q_in_679;
input q_in_678;
input q_in_677;
input q_in_676;
input q_in_675;
input q_in_674;
input q_in_673;
input q_in_672;
input q_in_671;
input q_in_670;
input q_in_669;
input q_in_668;
input q_in_667;
input q_in_666;
input q_in_665;
input q_in_664;
input q_in_663;
input q_in_662;
input q_in_661;
input q_in_660;
input q_in_659;
input q_in_658;
input q_in_657;
input q_in_656;
input q_in_655;
input q_in_654;
input q_in_653;
input q_in_652;
input q_in_651;
input q_in_650;
input q_in_649;
input q_in_648;
input q_in_647;
input q_in_646;
input q_in_645;
input q_in_644;
input q_in_643;
input q_in_642;
input q_in_641;
input q_in_640;
input q_in_639;
input q_in_638;
input q_in_637;
input q_in_636;
input q_in_635;
input q_in_634;
input q_in_633;
input q_in_632;
input q_in_631;
input q_in_630;
input q_in_629;
input q_in_628;
input q_in_627;
input q_in_626;
input q_in_625;
input q_in_624;
input q_in_623;
input q_in_622;
input q_in_621;
input q_in_620;
input q_in_619;
input q_in_618;
input q_in_617;
input q_in_616;
input q_in_615;
input q_in_614;
input q_in_613;
input q_in_612;
input q_in_611;
input q_in_610;
input q_in_609;
input q_in_608;
input q_in_607;
input q_in_606;
input q_in_605;
input q_in_604;
input q_in_603;
input q_in_602;
input q_in_601;
input q_in_600;
input q_in_599;
input q_in_598;
input q_in_597;
input q_in_596;
input q_in_595;
input q_in_594;
input q_in_593;
input q_in_592;
input q_in_591;
input q_in_590;
input q_in_589;
input q_in_588;
input q_in_587;
input q_in_586;
input q_in_585;
input q_in_584;
input q_in_583;
input q_in_582;
input q_in_581;
input q_in_580;
input q_in_579;
input q_in_578;
input q_in_577;
input q_in_576;
input q_in_575;
input q_in_574;
input q_in_573;
input q_in_572;
input q_in_571;
input q_in_570;
input q_in_569;
input q_in_568;
input q_in_567;
input q_in_566;
input q_in_565;
input q_in_564;
input q_in_563;
input q_in_562;
input q_in_561;
input q_in_560;
input q_in_559;
input q_in_558;
input q_in_557;
input q_in_556;
input q_in_555;
input q_in_554;
input q_in_553;
input q_in_552;
input q_in_551;
input q_in_550;
input q_in_549;
input q_in_548;
input q_in_547;
input q_in_546;
input q_in_545;
input q_in_544;
input q_in_543;
input q_in_542;
input q_in_541;
input q_in_540;
input q_in_539;
input q_in_538;
input q_in_537;
input q_in_536;
input q_in_535;
input q_in_534;
input q_in_533;
input q_in_532;
input q_in_531;
input q_in_530;
input q_in_529;
input q_in_528;
input q_in_527;
input q_in_526;
input q_in_525;
input q_in_524;
input q_in_523;
input q_in_522;
input q_in_521;
input q_in_520;
input q_in_519;
input q_in_518;
input q_in_517;
input q_in_516;
input q_in_515;
input q_in_514;
input q_in_513;
input q_in_512;
input q_in_511;
input q_in_510;
input q_in_509;
input q_in_508;
input q_in_507;
input q_in_506;
input q_in_505;
input q_in_504;
input q_in_503;
input q_in_502;
input q_in_501;
input q_in_500;
input q_in_499;
input q_in_498;
input q_in_497;
input q_in_496;
input q_in_495;
input q_in_494;
input q_in_493;
input q_in_492;
input q_in_491;
input q_in_490;
input q_in_489;
input q_in_488;
input q_in_487;
input q_in_486;
input q_in_485;
input q_in_484;
input q_in_483;
input q_in_482;
input q_in_481;
input q_in_480;
input q_in_479;
input q_in_478;
input q_in_477;
input q_in_476;
input q_in_475;
input q_in_474;
input q_in_473;
input q_in_472;
input q_in_471;
input q_in_470;
input q_in_469;
input q_in_468;
input q_in_467;
input q_in_466;
input q_in_465;
input q_in_464;
input q_in_463;
input q_in_462;
input q_in_461;
input q_in_460;
input q_in_459;
input q_in_458;
input q_in_457;
input q_in_456;
input q_in_455;
input q_in_454;
input q_in_453;
input q_in_452;
input q_in_451;
input q_in_450;
input q_in_449;
input q_in_448;
input q_in_447;
input q_in_446;
input q_in_445;
input q_in_444;
input q_in_443;
input q_in_442;
input q_in_441;
input q_in_440;
input q_in_439;
input q_in_438;
input q_in_437;
input q_in_436;
input q_in_435;
input q_in_434;
input q_in_433;
input q_in_432;
input q_in_431;
input q_in_430;
input q_in_429;
input q_in_428;
input q_in_427;
input q_in_426;
input q_in_425;
input q_in_424;
input q_in_423;
input q_in_422;
input q_in_421;
input q_in_420;
input q_in_419;
input q_in_418;
input q_in_417;
input q_in_416;
input q_in_415;
input q_in_414;
input q_in_413;
input q_in_412;
input q_in_411;
input q_in_410;
input q_in_409;
input q_in_408;
input q_in_407;
input q_in_406;
input q_in_405;
input q_in_404;
input q_in_403;
input q_in_402;
input q_in_401;
input q_in_400;
input q_in_399;
input q_in_398;
input q_in_397;
input q_in_396;
input q_in_395;
input q_in_394;
input q_in_393;
input q_in_392;
input q_in_391;
input q_in_390;
input q_in_389;
input q_in_388;
input q_in_387;
input q_in_386;
input q_in_385;
input q_in_384;
input q_in_383;
input q_in_382;
input q_in_381;
input q_in_380;
input q_in_379;
input q_in_378;
input q_in_377;
input q_in_376;
input q_in_375;
input q_in_374;
input q_in_373;
input q_in_372;
input q_in_371;
input q_in_370;
input q_in_369;
input q_in_368;
input q_in_367;
input q_in_366;
input q_in_365;
input q_in_364;
input q_in_363;
input q_in_362;
input q_in_361;
input q_in_360;
input q_in_359;
input q_in_358;
input q_in_357;
input q_in_356;
input q_in_355;
input q_in_354;
input q_in_353;
input q_in_352;
input q_in_351;
input q_in_350;
input q_in_349;
input q_in_348;
input q_in_347;
input q_in_346;
input q_in_345;
input q_in_344;
input q_in_343;
input q_in_342;
input q_in_341;
input q_in_340;
input q_in_339;
input q_in_338;
input q_in_337;
input q_in_336;
input q_in_335;
input q_in_334;
input q_in_333;
input q_in_332;
input q_in_331;
input q_in_330;
input q_in_329;
input q_in_328;
input q_in_327;
input q_in_326;
input q_in_325;
input q_in_324;
input q_in_323;
input q_in_322;
input q_in_321;
input q_in_320;
input q_in_319;
input q_in_318;
input q_in_317;
input q_in_316;
input q_in_315;
input q_in_314;
input q_in_313;
input q_in_312;
input q_in_311;
input q_in_310;
input q_in_309;
input q_in_308;
input q_in_307;
input q_in_306;
input q_in_305;
input q_in_304;
input q_in_303;
input q_in_302;
input q_in_301;
input q_in_300;
input q_in_299;
input q_in_298;
input q_in_297;
input q_in_296;
input q_in_295;
input q_in_294;
input q_in_293;
input q_in_292;
input q_in_291;
input q_in_290;
input q_in_289;
input q_in_288;
input q_in_287;
input q_in_286;
input q_in_285;
input q_in_284;
input q_in_283;
input q_in_282;
input q_in_281;
input q_in_280;
input q_in_279;
input q_in_278;
input q_in_277;
input q_in_276;
input q_in_275;
input q_in_274;
input q_in_273;
input q_in_272;
input q_in_271;
input q_in_270;
input q_in_269;
input q_in_268;
input q_in_267;
input q_in_266;
input q_in_265;
input q_in_264;
input q_in_263;
input q_in_262;
input q_in_261;
input q_in_260;
input q_in_259;
input q_in_258;
input q_in_257;
input q_in_256;
input q_in_255;
input q_in_254;
input q_in_253;
input q_in_252;
input q_in_251;
input q_in_250;
input q_in_249;
input q_in_248;
input q_in_247;
input q_in_246;
input q_in_245;
input q_in_244;
input q_in_243;
input q_in_242;
input q_in_241;
input q_in_240;
input q_in_239;
input q_in_238;
input q_in_237;
input q_in_236;
input q_in_235;
input q_in_234;
input q_in_233;
input q_in_232;
input q_in_231;
input q_in_230;
input q_in_229;
input q_in_228;
input q_in_227;
input q_in_226;
input q_in_225;
input q_in_224;
input q_in_223;
input q_in_222;
input q_in_221;
input q_in_220;
input q_in_219;
input q_in_218;
input q_in_217;
input q_in_216;
input q_in_215;
input q_in_214;
input q_in_213;
input q_in_212;
input q_in_211;
input q_in_210;
input q_in_209;
input q_in_208;
input q_in_207;
input q_in_206;
input q_in_205;
input q_in_204;
input q_in_203;
input q_in_202;
input q_in_201;
input q_in_200;
input q_in_199;
input q_in_198;
input q_in_197;
input q_in_196;
input q_in_195;
input q_in_194;
input q_in_193;
input q_in_192;
input q_in_191;
input q_in_190;
input q_in_189;
input q_in_188;
input q_in_187;
input q_in_186;
input q_in_185;
input q_in_184;
input q_in_183;
input q_in_182;
input q_in_181;
input q_in_180;
input q_in_179;
input q_in_178;
input q_in_177;
input q_in_176;
input q_in_175;
input q_in_174;
input q_in_173;
input q_in_172;
input q_in_171;
input q_in_170;
input q_in_169;
input q_in_168;
input q_in_167;
input q_in_166;
input q_in_165;
input q_in_164;
input q_in_163;
input q_in_162;
input q_in_161;
input q_in_160;
input q_in_159;
input q_in_158;
input q_in_157;
input q_in_156;
input q_in_155;
input q_in_154;
input q_in_153;
input q_in_152;
input q_in_151;
input q_in_150;
input q_in_149;
input q_in_148;
input q_in_147;
input q_in_146;
input q_in_145;
input q_in_144;
input q_in_143;
input q_in_142;
input q_in_141;
input q_in_140;
input q_in_139;
input q_in_138;
input q_in_137;
input q_in_136;
input q_in_135;
input q_in_134;
input q_in_133;
input q_in_132;
input q_in_131;
input q_in_130;
input q_in_129;
input q_in_128;
input q_in_127;
input q_in_126;
input q_in_125;
input q_in_124;
input q_in_123;
input q_in_122;
input q_in_121;
input q_in_120;
input q_in_119;
input q_in_118;
input q_in_117;
input q_in_116;
input q_in_115;
input q_in_114;
input q_in_113;
input q_in_112;
input q_in_111;
input q_in_110;
input q_in_109;
input q_in_108;
input q_in_107;
input q_in_106;
input q_in_105;
input q_in_104;
input q_in_103;
input q_in_102;
input q_in_101;
input q_in_100;
input q_in_99;
input q_in_98;
input q_in_97;
input q_in_96;
input q_in_95;
input q_in_94;
input q_in_93;
input q_in_92;
input q_in_91;
input q_in_90;
input q_in_89;
input q_in_88;
input q_in_87;
input q_in_86;
input q_in_85;
input q_in_84;
input q_in_83;
input q_in_82;
input q_in_81;
input q_in_80;
input q_in_79;
input q_in_78;
input q_in_77;
input q_in_76;
input q_in_75;
input q_in_74;
input q_in_73;
input q_in_72;
input q_in_71;
input q_in_70;
input q_in_69;
input q_in_68;
input q_in_67;
input q_in_66;
input q_in_65;
input q_in_64;
input q_in_63;
input q_in_62;
input q_in_61;
input q_in_60;
input q_in_59;
input q_in_58;
input q_in_57;
input q_in_56;
input q_in_55;
input q_in_54;
input q_in_53;
input q_in_52;
input q_in_51;
input q_in_50;
input q_in_49;
input q_in_48;
input q_in_47;
input q_in_46;
input q_in_45;
input q_in_44;
input q_in_43;
input q_in_42;
input q_in_41;
input q_in_40;
input q_in_39;
input q_in_38;
input q_in_37;
input q_in_36;
input q_in_35;
input q_in_34;
input q_in_33;
input q_in_32;
input q_in_31;
input q_in_30;
input q_in_29;
input q_in_28;
input q_in_27;
input q_in_26;
input q_in_25;
input q_in_24;
input q_in_23;
input q_in_22;
input q_in_21;
input q_in_20;
input q_in_19;
input q_in_18;
input q_in_17;
input q_in_16;
input q_in_15;
input q_in_14;
input q_in_13;
input q_in_12;
input q_in_11;
input q_in_10;
input q_in_9;
input q_in_8;
input q_in_7;
input q_in_6;
input q_in_5;
input q_in_4;
input q_in_3;
input q_in_2;
input q_in_1;
input clk_i, rst_i, cmd_w_i;
input [2:0] cmd_i;
input [31:0] text_i;
output d_out_910;
output d_out_909;
output d_out_908;
output d_out_907;
output d_out_906;
output d_out_905;
output d_out_904;
output d_out_903;
output d_out_902;
output d_out_901;
output d_out_900;
output d_out_899;
output d_out_898;
output d_out_897;
output d_out_896;
output d_out_895;
output d_out_894;
output d_out_893;
output d_out_892;
output d_out_891;
output d_out_890;
output d_out_889;
output d_out_888;
output d_out_887;
output d_out_886;
output d_out_885;
output d_out_884;
output d_out_883;
output d_out_882;
output d_out_881;
output d_out_880;
output d_out_879;
output d_out_878;
output d_out_877;
output d_out_876;
output d_out_875;
output d_out_874;
output d_out_873;
output d_out_872;
output d_out_871;
output d_out_870;
output d_out_869;
output d_out_868;
output d_out_867;
output d_out_866;
output d_out_865;
output d_out_864;
output d_out_863;
output d_out_862;
output d_out_861;
output d_out_860;
output d_out_859;
output d_out_858;
output d_out_857;
output d_out_856;
output d_out_855;
output d_out_854;
output d_out_853;
output d_out_852;
output d_out_851;
output d_out_850;
output d_out_849;
output d_out_848;
output d_out_847;
output d_out_846;
output d_out_845;
output d_out_844;
output d_out_843;
output d_out_842;
output d_out_841;
output d_out_840;
output d_out_839;
output d_out_838;
output d_out_837;
output d_out_836;
output d_out_835;
output d_out_834;
output d_out_833;
output d_out_832;
output d_out_831;
output d_out_830;
output d_out_829;
output d_out_828;
output d_out_827;
output d_out_826;
output d_out_825;
output d_out_824;
output d_out_823;
output d_out_822;
output d_out_821;
output d_out_820;
output d_out_819;
output d_out_818;
output d_out_817;
output d_out_816;
output d_out_815;
output d_out_814;
output d_out_813;
output d_out_812;
output d_out_811;
output d_out_810;
output d_out_809;
output d_out_808;
output d_out_807;
output d_out_806;
output d_out_805;
output d_out_804;
output d_out_803;
output d_out_802;
output d_out_801;
output d_out_800;
output d_out_799;
output d_out_798;
output d_out_797;
output d_out_796;
output d_out_795;
output d_out_794;
output d_out_793;
output d_out_792;
output d_out_791;
output d_out_790;
output d_out_789;
output d_out_788;
output d_out_787;
output d_out_786;
output d_out_785;
output d_out_784;
output d_out_783;
output d_out_782;
output d_out_781;
output d_out_780;
output d_out_779;
output d_out_778;
output d_out_777;
output d_out_776;
output d_out_775;
output d_out_774;
output d_out_773;
output d_out_772;
output d_out_771;
output d_out_770;
output d_out_769;
output d_out_768;
output d_out_767;
output d_out_766;
output d_out_765;
output d_out_764;
output d_out_763;
output d_out_762;
output d_out_761;
output d_out_760;
output d_out_759;
output d_out_758;
output d_out_757;
output d_out_756;
output d_out_755;
output d_out_754;
output d_out_753;
output d_out_752;
output d_out_751;
output d_out_750;
output d_out_749;
output d_out_748;
output d_out_747;
output d_out_746;
output d_out_745;
output d_out_744;
output d_out_743;
output d_out_742;
output d_out_741;
output d_out_740;
output d_out_739;
output d_out_738;
output d_out_737;
output d_out_736;
output d_out_735;
output d_out_734;
output d_out_733;
output d_out_732;
output d_out_731;
output d_out_730;
output d_out_729;
output d_out_728;
output d_out_727;
output d_out_726;
output d_out_725;
output d_out_724;
output d_out_723;
output d_out_722;
output d_out_721;
output d_out_720;
output d_out_719;
output d_out_718;
output d_out_717;
output d_out_716;
output d_out_715;
output d_out_714;
output d_out_713;
output d_out_712;
output d_out_711;
output d_out_710;
output d_out_709;
output d_out_708;
output d_out_707;
output d_out_706;
output d_out_705;
output d_out_704;
output d_out_703;
output d_out_702;
output d_out_701;
output d_out_700;
output d_out_699;
output d_out_698;
output d_out_697;
output d_out_696;
output d_out_695;
output d_out_694;
output d_out_693;
output d_out_692;
output d_out_691;
output d_out_690;
output d_out_689;
output d_out_688;
output d_out_687;
output d_out_686;
output d_out_685;
output d_out_684;
output d_out_683;
output d_out_682;
output d_out_681;
output d_out_680;
output d_out_679;
output d_out_678;
output d_out_677;
output d_out_676;
output d_out_675;
output d_out_674;
output d_out_673;
output d_out_672;
output d_out_671;
output d_out_670;
output d_out_669;
output d_out_668;
output d_out_667;
output d_out_666;
output d_out_665;
output d_out_664;
output d_out_663;
output d_out_662;
output d_out_661;
output d_out_660;
output d_out_659;
output d_out_658;
output d_out_657;
output d_out_656;
output d_out_655;
output d_out_654;
output d_out_653;
output d_out_652;
output d_out_651;
output d_out_650;
output d_out_649;
output d_out_648;
output d_out_647;
output d_out_646;
output d_out_645;
output d_out_644;
output d_out_643;
output d_out_642;
output d_out_641;
output d_out_640;
output d_out_639;
output d_out_638;
output d_out_637;
output d_out_636;
output d_out_635;
output d_out_634;
output d_out_633;
output d_out_632;
output d_out_631;
output d_out_630;
output d_out_629;
output d_out_628;
output d_out_627;
output d_out_626;
output d_out_625;
output d_out_624;
output d_out_623;
output d_out_622;
output d_out_621;
output d_out_620;
output d_out_619;
output d_out_618;
output d_out_617;
output d_out_616;
output d_out_615;
output d_out_614;
output d_out_613;
output d_out_612;
output d_out_611;
output d_out_610;
output d_out_609;
output d_out_608;
output d_out_607;
output d_out_606;
output d_out_605;
output d_out_604;
output d_out_603;
output d_out_602;
output d_out_601;
output d_out_600;
output d_out_599;
output d_out_598;
output d_out_597;
output d_out_596;
output d_out_595;
output d_out_594;
output d_out_593;
output d_out_592;
output d_out_591;
output d_out_590;
output d_out_589;
output d_out_588;
output d_out_587;
output d_out_586;
output d_out_585;
output d_out_584;
output d_out_583;
output d_out_582;
output d_out_581;
output d_out_580;
output d_out_579;
output d_out_578;
output d_out_577;
output d_out_576;
output d_out_575;
output d_out_574;
output d_out_573;
output d_out_572;
output d_out_571;
output d_out_570;
output d_out_569;
output d_out_568;
output d_out_567;
output d_out_566;
output d_out_565;
output d_out_564;
output d_out_563;
output d_out_562;
output d_out_561;
output d_out_560;
output d_out_559;
output d_out_558;
output d_out_557;
output d_out_556;
output d_out_555;
output d_out_554;
output d_out_553;
output d_out_552;
output d_out_551;
output d_out_550;
output d_out_549;
output d_out_548;
output d_out_547;
output d_out_546;
output d_out_545;
output d_out_544;
output d_out_543;
output d_out_542;
output d_out_541;
output d_out_540;
output d_out_539;
output d_out_538;
output d_out_537;
output d_out_536;
output d_out_535;
output d_out_534;
output d_out_533;
output d_out_532;
output d_out_531;
output d_out_530;
output d_out_529;
output d_out_528;
output d_out_527;
output d_out_526;
output d_out_525;
output d_out_524;
output d_out_523;
output d_out_522;
output d_out_521;
output d_out_520;
output d_out_519;
output d_out_518;
output d_out_517;
output d_out_516;
output d_out_515;
output d_out_514;
output d_out_513;
output d_out_512;
output d_out_511;
output d_out_510;
output d_out_509;
output d_out_508;
output d_out_507;
output d_out_506;
output d_out_505;
output d_out_504;
output d_out_503;
output d_out_502;
output d_out_501;
output d_out_500;
output d_out_499;
output d_out_498;
output d_out_497;
output d_out_496;
output d_out_495;
output d_out_494;
output d_out_493;
output d_out_492;
output d_out_491;
output d_out_490;
output d_out_489;
output d_out_488;
output d_out_487;
output d_out_486;
output d_out_485;
output d_out_484;
output d_out_483;
output d_out_482;
output d_out_481;
output d_out_480;
output d_out_479;
output d_out_478;
output d_out_477;
output d_out_476;
output d_out_475;
output d_out_474;
output d_out_473;
output d_out_472;
output d_out_471;
output d_out_470;
output d_out_469;
output d_out_468;
output d_out_467;
output d_out_466;
output d_out_465;
output d_out_464;
output d_out_463;
output d_out_462;
output d_out_461;
output d_out_460;
output d_out_459;
output d_out_458;
output d_out_457;
output d_out_456;
output d_out_455;
output d_out_454;
output d_out_453;
output d_out_452;
output d_out_451;
output d_out_450;
output d_out_449;
output d_out_448;
output d_out_447;
output d_out_446;
output d_out_445;
output d_out_444;
output d_out_443;
output d_out_442;
output d_out_441;
output d_out_440;
output d_out_439;
output d_out_438;
output d_out_437;
output d_out_436;
output d_out_435;
output d_out_434;
output d_out_433;
output d_out_432;
output d_out_431;
output d_out_430;
output d_out_429;
output d_out_428;
output d_out_427;
output d_out_426;
output d_out_425;
output d_out_424;
output d_out_423;
output d_out_422;
output d_out_421;
output d_out_420;
output d_out_419;
output d_out_418;
output d_out_417;
output d_out_416;
output d_out_415;
output d_out_414;
output d_out_413;
output d_out_412;
output d_out_411;
output d_out_410;
output d_out_409;
output d_out_408;
output d_out_407;
output d_out_406;
output d_out_405;
output d_out_404;
output d_out_403;
output d_out_402;
output d_out_401;
output d_out_400;
output d_out_399;
output d_out_398;
output d_out_397;
output d_out_396;
output d_out_395;
output d_out_394;
output d_out_393;
output d_out_392;
output d_out_391;
output d_out_390;
output d_out_389;
output d_out_388;
output d_out_387;
output d_out_386;
output d_out_385;
output d_out_384;
output d_out_383;
output d_out_382;
output d_out_381;
output d_out_380;
output d_out_379;
output d_out_378;
output d_out_377;
output d_out_376;
output d_out_375;
output d_out_374;
output d_out_373;
output d_out_372;
output d_out_371;
output d_out_370;
output d_out_369;
output d_out_368;
output d_out_367;
output d_out_366;
output d_out_365;
output d_out_364;
output d_out_363;
output d_out_362;
output d_out_361;
output d_out_360;
output d_out_359;
output d_out_358;
output d_out_357;
output d_out_356;
output d_out_355;
output d_out_354;
output d_out_353;
output d_out_352;
output d_out_351;
output d_out_350;
output d_out_349;
output d_out_348;
output d_out_347;
output d_out_346;
output d_out_345;
output d_out_344;
output d_out_343;
output d_out_342;
output d_out_341;
output d_out_340;
output d_out_339;
output d_out_338;
output d_out_337;
output d_out_336;
output d_out_335;
output d_out_334;
output d_out_333;
output d_out_332;
output d_out_331;
output d_out_330;
output d_out_329;
output d_out_328;
output d_out_327;
output d_out_326;
output d_out_325;
output d_out_324;
output d_out_323;
output d_out_322;
output d_out_321;
output d_out_320;
output d_out_319;
output d_out_318;
output d_out_317;
output d_out_316;
output d_out_315;
output d_out_314;
output d_out_313;
output d_out_312;
output d_out_311;
output d_out_310;
output d_out_309;
output d_out_308;
output d_out_307;
output d_out_306;
output d_out_305;
output d_out_304;
output d_out_303;
output d_out_302;
output d_out_301;
output d_out_300;
output d_out_299;
output d_out_298;
output d_out_297;
output d_out_296;
output d_out_295;
output d_out_294;
output d_out_293;
output d_out_292;
output d_out_291;
output d_out_290;
output d_out_289;
output d_out_288;
output d_out_287;
output d_out_286;
output d_out_285;
output d_out_284;
output d_out_283;
output d_out_282;
output d_out_281;
output d_out_280;
output d_out_279;
output d_out_278;
output d_out_277;
output d_out_276;
output d_out_275;
output d_out_274;
output d_out_273;
output d_out_272;
output d_out_271;
output d_out_270;
output d_out_269;
output d_out_268;
output d_out_267;
output d_out_266;
output d_out_265;
output d_out_264;
output d_out_263;
output d_out_262;
output d_out_261;
output d_out_260;
output d_out_259;
output d_out_258;
output d_out_257;
output d_out_256;
output d_out_255;
output d_out_254;
output d_out_253;
output d_out_252;
output d_out_251;
output d_out_250;
output d_out_249;
output d_out_248;
output d_out_247;
output d_out_246;
output d_out_245;
output d_out_244;
output d_out_243;
output d_out_242;
output d_out_241;
output d_out_240;
output d_out_239;
output d_out_238;
output d_out_237;
output d_out_236;
output d_out_235;
output d_out_234;
output d_out_233;
output d_out_232;
output d_out_231;
output d_out_230;
output d_out_229;
output d_out_228;
output d_out_227;
output d_out_226;
output d_out_225;
output d_out_224;
output d_out_223;
output d_out_222;
output d_out_221;
output d_out_220;
output d_out_219;
output d_out_218;
output d_out_217;
output d_out_216;
output d_out_215;
output d_out_214;
output d_out_213;
output d_out_212;
output d_out_211;
output d_out_210;
output d_out_209;
output d_out_208;
output d_out_207;
output d_out_206;
output d_out_205;
output d_out_204;
output d_out_203;
output d_out_202;
output d_out_201;
output d_out_200;
output d_out_199;
output d_out_198;
output d_out_197;
output d_out_196;
output d_out_195;
output d_out_194;
output d_out_193;
output d_out_192;
output d_out_191;
output d_out_190;
output d_out_189;
output d_out_188;
output d_out_187;
output d_out_186;
output d_out_185;
output d_out_184;
output d_out_183;
output d_out_182;
output d_out_181;
output d_out_180;
output d_out_179;
output d_out_178;
output d_out_177;
output d_out_176;
output d_out_175;
output d_out_174;
output d_out_173;
output d_out_172;
output d_out_171;
output d_out_170;
output d_out_169;
output d_out_168;
output d_out_167;
output d_out_166;
output d_out_165;
output d_out_164;
output d_out_163;
output d_out_162;
output d_out_161;
output d_out_160;
output d_out_159;
output d_out_158;
output d_out_157;
output d_out_156;
output d_out_155;
output d_out_154;
output d_out_153;
output d_out_152;
output d_out_151;
output d_out_150;
output d_out_149;
output d_out_148;
output d_out_147;
output d_out_146;
output d_out_145;
output d_out_144;
output d_out_143;
output d_out_142;
output d_out_141;
output d_out_140;
output d_out_139;
output d_out_138;
output d_out_137;
output d_out_136;
output d_out_135;
output d_out_134;
output d_out_133;
output d_out_132;
output d_out_131;
output d_out_130;
output d_out_129;
output d_out_128;
output d_out_127;
output d_out_126;
output d_out_125;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_121;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_116;
output d_out_115;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_111;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_83;
output d_out_82;
output d_out_81;
output d_out_80;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_76;
output d_out_75;
output d_out_74;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_64;
output d_out_63;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_50;
output d_out_49;
output d_out_48;
output d_out_47;
output d_out_46;
output d_out_45;
output d_out_44;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_30;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_5;
output d_out_4;
output d_out_3;
output d_out_2;
output d_out_1;
output [3:0] cmd_o;
output [31:0] text_o;
wire [2:0] read_counter;
wire [31:0] H4;
wire [31:0] H3;
wire [31:0] H2;
wire [31:0] H1;
wire [31:0] H0;
wire [95:0] SHA1_result;
wire [31:0] next_C;
wire [31:0] next_A;
wire [31:0] Wt;
wire [31:0] Kt;
wire [31:0] SHA1_ft_BCD;
wire [5:0] round;
wire SHA1_result_151, SHA1_result_148, SHA1_result_136, SHA1_result_135, SHA1_result_134, SHA1_result_133, SHA1_result_132, SHA1_result_131, SHA1_result_130, SHA1_result_129, SHA1_result_128, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, 
  N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, 
  N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, 
  N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1715, N1716, N1717, N1718, N1719, N1720, N2583, N2585, N2587, N2589, N2590, N2592, N2595, n341, n345, n347, n412, n422, n423, n433, n437, n438, n440, n442, n443, n444, n445, n446, n447, n448, 
  n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n470, n471, n472, n473, n474, n475, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, 
  n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, 
  n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, 
  n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, 
  n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, 
  n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, 
  n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, 
  n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, 
  n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, 
  n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, 
  n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, 
  n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, 
  n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, 
  n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, 
  n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, 
  n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, 
  n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, 
  n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n8262, n8264, 
  n8266, n8268, n8270, n8272, n8274, n8276, n8278, n8280, n8282, n8284, n8286, n8288, n8290, n8292, n8294, n8296, n8298, n8300, n8302, n8304, n8306, n8308, n8310, n8312, n8314, n8316, n8318, n8320, n8322, n8323, n8326, n8328, n8330, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, 
  N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
  N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, n9299, n9300, n9301, n9302, n9303, n9304, n9308, n9309, n9310, n9311, n9313, n9314, n9315, n9316, n9317, n9325, n9326, n9327, n9332, n9333, n9334, 
  n9338, n9339, n9340, n9344, n9345, n9346, n9350, n9351, n9352, n9356, n9357, n9358, n9362, n9363, n9364, n9368, n9369, n9370, n9374, n9375, n9376, n9380, n9381, n9382, n9386, n9387, n9388, n9392, n9393, n9394, n9398, n9399, n9400, n9404, n9405, n9406, n9410, n9411, n9412, n9416, n9417, n9418, n9422, n9423, n9424, n9428, n9429, n9430, n9431, n9432, 
  n9434, n9435, n9436, n9437, n9438, n9440, n9441, n9442, n9443, n9444, n9446, n9447, n9448, n9449, n9450, n9452, n9453, n9454, n9455, n9456, n9458, n9459, n9460, n9461, n9462, n9464, n9465, n9466, n9467, n9468, n9470, n9471, n9472, n9473, n9474, n9476, n9477, n9478, n9479, n9480, n9482, n9483, n9484, n9485, n9486, n9488, n9489, n9490, n9491, n9492, 
  n9494, n9495, n9496, n9497, n9498, n9500, n9501, n9502, n9503, n9504, n9506, n9507, n9508, n9509, n9510, n9512, n9513, n9514, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, 
  n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9621, n9622, n9623, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, 
  n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, 
  n9713, n9714, n9715, n9716, n9717, n9718, n9721, n9722, n9723, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, 
  n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, 
  n9817, n9818, n9820, n9821, n9822, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, 
  n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9921, n9922, 
  n9923, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, 
  n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10025, n10026, 
  n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, 
  n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, 
  n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, 
  n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, 
  n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, 
  n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10313, n10314, n10315, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, 
  n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, 
  n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, 
  n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, 
  n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, 
  n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, 
  n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, 
  n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, 
  n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10711, n10712, n10713, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, 
  n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, 
  n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10810, n10811, n10812, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, 
  n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, 
  n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10909, n10910, n10911, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, 
  n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, 
  n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11114, n11835, n11836, n11837, n11838, n11839, n11840, n11843, n11844, n11845, n11846, n11853, n11865, n11872, n11879, n11886, n11893, n11900, n11907, n11914, n11921, n11928, n11935, n11942, n11949, n11956, n11963, n11970, n11977, n11984, n11991, n11998, n11999, n12000, n12001, n12002, n12005, n12006, n12007, n12008, n12009, n12010, n12011, 
  n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12047, n12048, n12049, n12050, n12051, n12054, n12055, n12056, n12057, n12058, n12061, n12062, n12063, n12064, n12065, n12068, n12069, 
  n12070, n12071, n12072, n12075, n12076, n12077, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, 
  n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12916, n12918, n12920, n12922, n12924, n12926, n12928, n12930, n12932, n12934, n12936, n12938, n12940, n12942, n12944, n12946, n12948, n12950, n12952, n12954, n12956, n12958, n12960, n12962, n12964, n12966, n12968, n12970, n12972, n12974, 
  n12976, n12978, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, 
  n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, 
  n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, 
  n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, 
  n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, 
  n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, 
  n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, 
  n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, 
  n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, 
  n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, 
  n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, 
  n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, 
  n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, 
  n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, 
  n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, 
  n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, 
  n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, 
  n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, 
  n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, 
  n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, 
  n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, 
  n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, 
  n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, 
  n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, 
  n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, 
  n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, 
  n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, 
  n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, 
  n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, 
  n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, 
  n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, 
  n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, 
  n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, 
  n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, 
  n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, 
  n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, 
  n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, 
  n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, 
  n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, 
  n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, 
  n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, 
  n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, 
  n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, 
  n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, 
  n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, 
  n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, 
  n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, 
  n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, 
  n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, _add_3_root_add_136_4_n403, 
  _add_3_root_add_136_4_n402, _add_3_root_add_136_4_n401, _add_3_root_add_136_4_n400, _add_3_root_add_136_4_n399, _add_3_root_add_136_4_n398, _add_3_root_add_136_4_n397, _add_3_root_add_136_4_n396, _add_3_root_add_136_4_n395, _add_3_root_add_136_4_n394, _add_3_root_add_136_4_n393, _add_3_root_add_136_4_n392, _add_3_root_add_136_4_n391, _add_3_root_add_136_4_n390, _add_3_root_add_136_4_n389, _add_3_root_add_136_4_n388, _add_3_root_add_136_4_n387, _add_3_root_add_136_4_n386, _add_3_root_add_136_4_n385, _add_3_root_add_136_4_n384, _add_3_root_add_136_4_n383, _add_3_root_add_136_4_n382, _add_3_root_add_136_4_n381, _add_3_root_add_136_4_n380, _add_3_root_add_136_4_n379, _add_3_root_add_136_4_n378, _add_3_root_add_136_4_n377, _add_3_root_add_136_4_n376, _add_3_root_add_136_4_n375, _add_3_root_add_136_4_n374, _add_3_root_add_136_4_n373, _add_3_root_add_136_4_n372, _add_3_root_add_136_4_n371, _add_3_root_add_136_4_n370, _add_3_root_add_136_4_n369, _add_3_root_add_136_4_n368, _add_3_root_add_136_4_n367, _add_3_root_add_136_4_n366, _add_3_root_add_136_4_n365, _add_3_root_add_136_4_n364, _add_3_root_add_136_4_n363, _add_3_root_add_136_4_n362, _add_3_root_add_136_4_n361, _add_3_root_add_136_4_n360, _add_3_root_add_136_4_n359, _add_3_root_add_136_4_n358, _add_3_root_add_136_4_n357, _add_3_root_add_136_4_n356, _add_3_root_add_136_4_n355, _add_3_root_add_136_4_n354, _add_3_root_add_136_4_n353, 
  _add_3_root_add_136_4_n352, _add_3_root_add_136_4_n351, _add_3_root_add_136_4_n350, _add_3_root_add_136_4_n349, _add_3_root_add_136_4_n348, _add_3_root_add_136_4_n347, _add_3_root_add_136_4_n346, _add_3_root_add_136_4_n345, _add_3_root_add_136_4_n344, _add_3_root_add_136_4_n343, _add_3_root_add_136_4_n342, _add_3_root_add_136_4_n341, _add_3_root_add_136_4_n340, _add_3_root_add_136_4_n339, _add_3_root_add_136_4_n338, _add_3_root_add_136_4_n337, _add_3_root_add_136_4_n336, _add_3_root_add_136_4_n335, _add_3_root_add_136_4_n334, _add_3_root_add_136_4_n333, _add_3_root_add_136_4_n332, _add_3_root_add_136_4_n331, _add_3_root_add_136_4_n330, _add_3_root_add_136_4_n329, _add_3_root_add_136_4_n328, _add_3_root_add_136_4_n327, _add_3_root_add_136_4_n326, _add_3_root_add_136_4_n325, _add_3_root_add_136_4_n324, _add_3_root_add_136_4_n323, _add_3_root_add_136_4_n322, _add_3_root_add_136_4_n321, _add_3_root_add_136_4_n320, _add_3_root_add_136_4_n319, _add_3_root_add_136_4_n318, _add_3_root_add_136_4_n317, _add_3_root_add_136_4_n316, _add_3_root_add_136_4_n315, _add_3_root_add_136_4_n314, _add_3_root_add_136_4_n313, _add_3_root_add_136_4_n312, _add_3_root_add_136_4_n311, _add_3_root_add_136_4_n310, _add_3_root_add_136_4_n309, _add_3_root_add_136_4_n308, _add_3_root_add_136_4_n307, _add_3_root_add_136_4_n306, _add_3_root_add_136_4_n305, _add_3_root_add_136_4_n304, _add_3_root_add_136_4_n303, 
  _add_3_root_add_136_4_n302, _add_3_root_add_136_4_n301, _add_3_root_add_136_4_n300, _add_3_root_add_136_4_n299, _add_3_root_add_136_4_n298, _add_3_root_add_136_4_n297, _add_3_root_add_136_4_n296, _add_3_root_add_136_4_n295, _add_3_root_add_136_4_n294, _add_3_root_add_136_4_n293, _add_3_root_add_136_4_n292, _add_3_root_add_136_4_n291, _add_3_root_add_136_4_n290, _add_3_root_add_136_4_n289, _add_3_root_add_136_4_n288, _add_3_root_add_136_4_n287, _add_3_root_add_136_4_n286, _add_3_root_add_136_4_n285, _add_3_root_add_136_4_n284, _add_3_root_add_136_4_n283, _add_3_root_add_136_4_n282, _add_3_root_add_136_4_n281, _add_3_root_add_136_4_n280, _add_3_root_add_136_4_n279, _add_3_root_add_136_4_n278, _add_3_root_add_136_4_n277, _add_3_root_add_136_4_n276, _add_3_root_add_136_4_n275, _add_3_root_add_136_4_n274, _add_3_root_add_136_4_n273, _add_3_root_add_136_4_n272, _add_3_root_add_136_4_n271, _add_3_root_add_136_4_n270, _add_3_root_add_136_4_n269, _add_3_root_add_136_4_n268, _add_3_root_add_136_4_n267, _add_3_root_add_136_4_n266, _add_3_root_add_136_4_n265, _add_3_root_add_136_4_n264, _add_3_root_add_136_4_n263, _add_3_root_add_136_4_n262, _add_3_root_add_136_4_n261, _add_3_root_add_136_4_n260, _add_3_root_add_136_4_n259, _add_3_root_add_136_4_n258, _add_3_root_add_136_4_n257, _add_3_root_add_136_4_n256, _add_3_root_add_136_4_n255, _add_3_root_add_136_4_n254, _add_3_root_add_136_4_n253, 
  _add_3_root_add_136_4_n252, _add_3_root_add_136_4_n251, _add_3_root_add_136_4_n250, _add_3_root_add_136_4_n249, _add_3_root_add_136_4_n248, _add_3_root_add_136_4_n247, _add_3_root_add_136_4_n246, _add_3_root_add_136_4_n245, _add_3_root_add_136_4_n244, _add_3_root_add_136_4_n243, _add_3_root_add_136_4_n242, _add_3_root_add_136_4_n241, _add_3_root_add_136_4_n240, _add_3_root_add_136_4_n239, _add_3_root_add_136_4_n238, _add_3_root_add_136_4_n237, _add_3_root_add_136_4_n236, _add_3_root_add_136_4_n235, _add_3_root_add_136_4_n234, _add_3_root_add_136_4_n233, _add_3_root_add_136_4_n232, _add_3_root_add_136_4_n231, _add_3_root_add_136_4_n230, _add_3_root_add_136_4_n229, _add_3_root_add_136_4_n228, _add_3_root_add_136_4_n227, _add_3_root_add_136_4_n226, _add_3_root_add_136_4_n225, _add_3_root_add_136_4_n224, _add_3_root_add_136_4_n223, _add_3_root_add_136_4_n222, _add_3_root_add_136_4_n221, _add_3_root_add_136_4_n220, _add_3_root_add_136_4_n219, _add_3_root_add_136_4_n218, _add_3_root_add_136_4_n217, _add_3_root_add_136_4_n216, _add_3_root_add_136_4_n215, _add_3_root_add_136_4_n214, _add_3_root_add_136_4_n213, _add_3_root_add_136_4_n212, _add_3_root_add_136_4_n211, _add_3_root_add_136_4_n210, _add_3_root_add_136_4_n209, _add_3_root_add_136_4_n208, _add_3_root_add_136_4_n207, _add_3_root_add_136_4_n206, _add_3_root_add_136_4_n205, _add_3_root_add_136_4_n204, _add_3_root_add_136_4_n203, 
  _add_3_root_add_136_4_n202, _add_3_root_add_136_4_n201, _add_3_root_add_136_4_n200, _add_3_root_add_136_4_n199, _add_3_root_add_136_4_n198, _add_3_root_add_136_4_n197, _add_3_root_add_136_4_n196, _add_3_root_add_136_4_n195, _add_3_root_add_136_4_n194, _add_3_root_add_136_4_n193, _add_3_root_add_136_4_n192, _add_3_root_add_136_4_n191, _add_3_root_add_136_4_n190, _add_3_root_add_136_4_n189, _add_3_root_add_136_4_n188, _add_3_root_add_136_4_n187, _add_3_root_add_136_4_n186, _add_3_root_add_136_4_n185, _add_3_root_add_136_4_n184, _add_3_root_add_136_4_n183, _add_3_root_add_136_4_n182, _add_3_root_add_136_4_n181, _add_3_root_add_136_4_n180, _add_3_root_add_136_4_n179, _add_3_root_add_136_4_n178, _add_3_root_add_136_4_n177, _add_3_root_add_136_4_n176, _add_3_root_add_136_4_n175, _add_3_root_add_136_4_n174, _add_3_root_add_136_4_n173, _add_3_root_add_136_4_n172, _add_3_root_add_136_4_n171, _add_3_root_add_136_4_n170, _add_3_root_add_136_4_n169, _add_3_root_add_136_4_n168, _add_3_root_add_136_4_n167, _add_3_root_add_136_4_n166, _add_3_root_add_136_4_n165, _add_3_root_add_136_4_n164, _add_3_root_add_136_4_n163, _add_3_root_add_136_4_n162, _add_3_root_add_136_4_n161, _add_3_root_add_136_4_n160, _add_3_root_add_136_4_n159, _add_3_root_add_136_4_n158, _add_3_root_add_136_4_n157, _add_3_root_add_136_4_n156, _add_3_root_add_136_4_n155, _add_3_root_add_136_4_n154, _add_3_root_add_136_4_n153, 
  _add_3_root_add_136_4_n152, _add_3_root_add_136_4_n151, _add_3_root_add_136_4_n150, _add_3_root_add_136_4_n149, _add_3_root_add_136_4_n148, _add_3_root_add_136_4_n147, _add_3_root_add_136_4_n146, _add_3_root_add_136_4_n145, _add_3_root_add_136_4_n144, _add_3_root_add_136_4_n143, _add_3_root_add_136_4_n142, _add_3_root_add_136_4_n141, _add_3_root_add_136_4_n140, _add_3_root_add_136_4_n139, _add_3_root_add_136_4_n138, _add_3_root_add_136_4_n137, _add_3_root_add_136_4_n136, _add_3_root_add_136_4_n135, _add_3_root_add_136_4_n134, _add_3_root_add_136_4_n133, _add_3_root_add_136_4_n132, _add_3_root_add_136_4_n131, _add_3_root_add_136_4_n130, _add_3_root_add_136_4_n129, _add_3_root_add_136_4_n128, _add_3_root_add_136_4_n127, _add_3_root_add_136_4_n126, _add_3_root_add_136_4_n125, _add_3_root_add_136_4_n124, _add_3_root_add_136_4_n123, _add_3_root_add_136_4_n122, _add_3_root_add_136_4_n121, _add_3_root_add_136_4_n120, _add_3_root_add_136_4_n119, _add_3_root_add_136_4_n118, _add_3_root_add_136_4_n117, _add_3_root_add_136_4_n116, _add_3_root_add_136_4_n115, _add_3_root_add_136_4_n114, _add_3_root_add_136_4_n113, _add_3_root_add_136_4_n112, _add_3_root_add_136_4_n111, _add_3_root_add_136_4_n110, _add_3_root_add_136_4_n109, _add_3_root_add_136_4_n108, _add_3_root_add_136_4_n107, _add_3_root_add_136_4_n106, _add_3_root_add_136_4_n105, _add_3_root_add_136_4_n104, _add_3_root_add_136_4_n103, 
  _add_3_root_add_136_4_n102, _add_3_root_add_136_4_n101, _add_3_root_add_136_4_n100, _add_3_root_add_136_4_n99, _add_3_root_add_136_4_n98, _add_3_root_add_136_4_n97, _add_3_root_add_136_4_n96, _add_3_root_add_136_4_n95, _add_3_root_add_136_4_n94, _add_3_root_add_136_4_n93, _add_3_root_add_136_4_n92, _add_3_root_add_136_4_n91, _add_3_root_add_136_4_n90, _add_3_root_add_136_4_n89, _add_3_root_add_136_4_n87, _add_3_root_add_136_4_n86, _add_3_root_add_136_4_n85, _add_3_root_add_136_4_n84, _add_3_root_add_136_4_n83, _add_3_root_add_136_4_n81, _add_3_root_add_136_4_n80, _add_3_root_add_136_4_n79, _add_3_root_add_136_4_n78, _add_3_root_add_136_4_n76, _add_3_root_add_136_4_n73, _add_3_root_add_136_4_n72, _add_3_root_add_136_4_n71, _add_3_root_add_136_4_n70, _add_3_root_add_136_4_n69, _add_3_root_add_136_4_n68, _add_3_root_add_136_4_n67, _add_3_root_add_136_4_n66, _add_3_root_add_136_4_n65, _add_3_root_add_136_4_n64, _add_3_root_add_136_4_n63, _add_3_root_add_136_4_n62, _add_3_root_add_136_4_n61, _add_3_root_add_136_4_n60, _add_3_root_add_136_4_n59, _add_3_root_add_136_4_n58, _add_3_root_add_136_4_n57, _add_3_root_add_136_4_n56, _add_3_root_add_136_4_n55, _add_3_root_add_136_4_n54, _add_3_root_add_136_4_n53, _add_3_root_add_136_4_n52, _add_3_root_add_136_4_n50, _add_3_root_add_136_4_n48, _add_3_root_add_136_4_n47, _add_3_root_add_136_4_n46, 
  _add_3_root_add_136_4_n45, _add_3_root_add_136_4_n44, _add_3_root_add_136_4_n43, _add_3_root_add_136_4_n42, _add_3_root_add_136_4_n41, _add_3_root_add_136_4_n40, _add_3_root_add_136_4_n39, _add_3_root_add_136_4_n38, _add_3_root_add_136_4_n37, _add_3_root_add_136_4_n36, _add_3_root_add_136_4_n35, _add_3_root_add_136_4_n34, _add_3_root_add_136_4_n33, _add_3_root_add_136_4_n32, _add_3_root_add_136_4_n31, _add_3_root_add_136_4_n30, _add_3_root_add_136_4_n29, _add_3_root_add_136_4_n28, _add_3_root_add_136_4_n27, _add_3_root_add_136_4_n26, _add_3_root_add_136_4_n25, _add_3_root_add_136_4_n24, _add_3_root_add_136_4_n23, _add_3_root_add_136_4_n22, _add_3_root_add_136_4_n21, _add_3_root_add_136_4_n20, _add_3_root_add_136_4_n19, _add_3_root_add_136_4_n18, _add_3_root_add_136_4_n17, _add_3_root_add_136_4_n16, _add_3_root_add_136_4_n15, _add_3_root_add_136_4_n14, _add_3_root_add_136_4_n12, _add_3_root_add_136_4_n11, _add_3_root_add_136_4_n10, _add_3_root_add_136_4_n9, _add_3_root_add_136_4_n8, _add_3_root_add_136_4_n7, _add_3_root_add_136_4_n6, _add_3_root_add_136_4_n5, _add_3_root_add_136_4_n4, _add_3_root_add_136_4_n3, _add_3_root_add_136_4_n2, _add_2_root_add_136_4_n437, _add_2_root_add_136_4_n436, _add_2_root_add_136_4_n435, _add_2_root_add_136_4_n434, _add_2_root_add_136_4_n433, _add_2_root_add_136_4_n432, _add_2_root_add_136_4_n431, 
  _add_2_root_add_136_4_n430, _add_2_root_add_136_4_n429, _add_2_root_add_136_4_n428, _add_2_root_add_136_4_n427, _add_2_root_add_136_4_n426, _add_2_root_add_136_4_n425, _add_2_root_add_136_4_n424, _add_2_root_add_136_4_n423, _add_2_root_add_136_4_n422, _add_2_root_add_136_4_n421, _add_2_root_add_136_4_n420, _add_2_root_add_136_4_n419, _add_2_root_add_136_4_n418, _add_2_root_add_136_4_n417, _add_2_root_add_136_4_n416, _add_2_root_add_136_4_n415, _add_2_root_add_136_4_n414, _add_2_root_add_136_4_n413, _add_2_root_add_136_4_n412, _add_2_root_add_136_4_n411, _add_2_root_add_136_4_n410, _add_2_root_add_136_4_n409, _add_2_root_add_136_4_n408, _add_2_root_add_136_4_n407, _add_2_root_add_136_4_n406, _add_2_root_add_136_4_n405, _add_2_root_add_136_4_n404, _add_2_root_add_136_4_n403, _add_2_root_add_136_4_n402, _add_2_root_add_136_4_n401, _add_2_root_add_136_4_n400, _add_2_root_add_136_4_n399, _add_2_root_add_136_4_n398, _add_2_root_add_136_4_n397, _add_2_root_add_136_4_n396, _add_2_root_add_136_4_n395, _add_2_root_add_136_4_n394, _add_2_root_add_136_4_n393, _add_2_root_add_136_4_n392, _add_2_root_add_136_4_n391, _add_2_root_add_136_4_n390, _add_2_root_add_136_4_n389, _add_2_root_add_136_4_n388, _add_2_root_add_136_4_n387, _add_2_root_add_136_4_n386, _add_2_root_add_136_4_n385, _add_2_root_add_136_4_n384, _add_2_root_add_136_4_n383, _add_2_root_add_136_4_n382, _add_2_root_add_136_4_n381, 
  _add_2_root_add_136_4_n380, _add_2_root_add_136_4_n379, _add_2_root_add_136_4_n378, _add_2_root_add_136_4_n377, _add_2_root_add_136_4_n376, _add_2_root_add_136_4_n375, _add_2_root_add_136_4_n374, _add_2_root_add_136_4_n373, _add_2_root_add_136_4_n372, _add_2_root_add_136_4_n371, _add_2_root_add_136_4_n370, _add_2_root_add_136_4_n369, _add_2_root_add_136_4_n368, _add_2_root_add_136_4_n367, _add_2_root_add_136_4_n366, _add_2_root_add_136_4_n365, _add_2_root_add_136_4_n364, _add_2_root_add_136_4_n363, _add_2_root_add_136_4_n362, _add_2_root_add_136_4_n361, _add_2_root_add_136_4_n360, _add_2_root_add_136_4_n359, _add_2_root_add_136_4_n358, _add_2_root_add_136_4_n357, _add_2_root_add_136_4_n356, _add_2_root_add_136_4_n355, _add_2_root_add_136_4_n354, _add_2_root_add_136_4_n353, _add_2_root_add_136_4_n352, _add_2_root_add_136_4_n351, _add_2_root_add_136_4_n350, _add_2_root_add_136_4_n349, _add_2_root_add_136_4_n348, _add_2_root_add_136_4_n347, _add_2_root_add_136_4_n346, _add_2_root_add_136_4_n345, _add_2_root_add_136_4_n344, _add_2_root_add_136_4_n343, _add_2_root_add_136_4_n342, _add_2_root_add_136_4_n341, _add_2_root_add_136_4_n340, _add_2_root_add_136_4_n339, _add_2_root_add_136_4_n338, _add_2_root_add_136_4_n337, _add_2_root_add_136_4_n336, _add_2_root_add_136_4_n335, _add_2_root_add_136_4_n334, _add_2_root_add_136_4_n333, _add_2_root_add_136_4_n332, _add_2_root_add_136_4_n331, 
  _add_2_root_add_136_4_n330, _add_2_root_add_136_4_n329, _add_2_root_add_136_4_n328, _add_2_root_add_136_4_n327, _add_2_root_add_136_4_n326, _add_2_root_add_136_4_n325, _add_2_root_add_136_4_n324, _add_2_root_add_136_4_n323, _add_2_root_add_136_4_n322, _add_2_root_add_136_4_n321, _add_2_root_add_136_4_n320, _add_2_root_add_136_4_n319, _add_2_root_add_136_4_n318, _add_2_root_add_136_4_n317, _add_2_root_add_136_4_n316, _add_2_root_add_136_4_n315, _add_2_root_add_136_4_n314, _add_2_root_add_136_4_n313, _add_2_root_add_136_4_n312, _add_2_root_add_136_4_n311, _add_2_root_add_136_4_n310, _add_2_root_add_136_4_n309, _add_2_root_add_136_4_n308, _add_2_root_add_136_4_n307, _add_2_root_add_136_4_n306, _add_2_root_add_136_4_n305, _add_2_root_add_136_4_n304, _add_2_root_add_136_4_n303, _add_2_root_add_136_4_n302, _add_2_root_add_136_4_n301, _add_2_root_add_136_4_n300, _add_2_root_add_136_4_n299, _add_2_root_add_136_4_n298, _add_2_root_add_136_4_n297, _add_2_root_add_136_4_n296, _add_2_root_add_136_4_n295, _add_2_root_add_136_4_n294, _add_2_root_add_136_4_n293, _add_2_root_add_136_4_n292, _add_2_root_add_136_4_n291, _add_2_root_add_136_4_n290, _add_2_root_add_136_4_n289, _add_2_root_add_136_4_n288, _add_2_root_add_136_4_n287, _add_2_root_add_136_4_n286, _add_2_root_add_136_4_n285, _add_2_root_add_136_4_n284, _add_2_root_add_136_4_n283, _add_2_root_add_136_4_n282, _add_2_root_add_136_4_n281, 
  _add_2_root_add_136_4_n280, _add_2_root_add_136_4_n279, _add_2_root_add_136_4_n278, _add_2_root_add_136_4_n277, _add_2_root_add_136_4_n276, _add_2_root_add_136_4_n275, _add_2_root_add_136_4_n274, _add_2_root_add_136_4_n273, _add_2_root_add_136_4_n272, _add_2_root_add_136_4_n271, _add_2_root_add_136_4_n270, _add_2_root_add_136_4_n269, _add_2_root_add_136_4_n268, _add_2_root_add_136_4_n267, _add_2_root_add_136_4_n266, _add_2_root_add_136_4_n265, _add_2_root_add_136_4_n264, _add_2_root_add_136_4_n263, _add_2_root_add_136_4_n262, _add_2_root_add_136_4_n261, _add_2_root_add_136_4_n260, _add_2_root_add_136_4_n259, _add_2_root_add_136_4_n258, _add_2_root_add_136_4_n257, _add_2_root_add_136_4_n256, _add_2_root_add_136_4_n255, _add_2_root_add_136_4_n254, _add_2_root_add_136_4_n253, _add_2_root_add_136_4_n252, _add_2_root_add_136_4_n251, _add_2_root_add_136_4_n250, _add_2_root_add_136_4_n249, _add_2_root_add_136_4_n248, _add_2_root_add_136_4_n247, _add_2_root_add_136_4_n246, _add_2_root_add_136_4_n245, _add_2_root_add_136_4_n244, _add_2_root_add_136_4_n243, _add_2_root_add_136_4_n242, _add_2_root_add_136_4_n241, _add_2_root_add_136_4_n240, _add_2_root_add_136_4_n239, _add_2_root_add_136_4_n238, _add_2_root_add_136_4_n237, _add_2_root_add_136_4_n236, _add_2_root_add_136_4_n235, _add_2_root_add_136_4_n234, _add_2_root_add_136_4_n233, _add_2_root_add_136_4_n232, _add_2_root_add_136_4_n231, 
  _add_2_root_add_136_4_n230, _add_2_root_add_136_4_n229, _add_2_root_add_136_4_n228, _add_2_root_add_136_4_n227, _add_2_root_add_136_4_n226, _add_2_root_add_136_4_n225, _add_2_root_add_136_4_n224, _add_2_root_add_136_4_n223, _add_2_root_add_136_4_n222, _add_2_root_add_136_4_n221, _add_2_root_add_136_4_n220, _add_2_root_add_136_4_n219, _add_2_root_add_136_4_n218, _add_2_root_add_136_4_n217, _add_2_root_add_136_4_n216, _add_2_root_add_136_4_n215, _add_2_root_add_136_4_n214, _add_2_root_add_136_4_n213, _add_2_root_add_136_4_n212, _add_2_root_add_136_4_n211, _add_2_root_add_136_4_n210, _add_2_root_add_136_4_n209, _add_2_root_add_136_4_n208, _add_2_root_add_136_4_n207, _add_2_root_add_136_4_n206, _add_2_root_add_136_4_n205, _add_2_root_add_136_4_n204, _add_2_root_add_136_4_n203, _add_2_root_add_136_4_n202, _add_2_root_add_136_4_n201, _add_2_root_add_136_4_n200, _add_2_root_add_136_4_n199, _add_2_root_add_136_4_n198, _add_2_root_add_136_4_n197, _add_2_root_add_136_4_n196, _add_2_root_add_136_4_n195, _add_2_root_add_136_4_n194, _add_2_root_add_136_4_n193, _add_2_root_add_136_4_n192, _add_2_root_add_136_4_n191, _add_2_root_add_136_4_n190, _add_2_root_add_136_4_n189, _add_2_root_add_136_4_n188, _add_2_root_add_136_4_n187, _add_2_root_add_136_4_n186, _add_2_root_add_136_4_n185, _add_2_root_add_136_4_n184, _add_2_root_add_136_4_n183, _add_2_root_add_136_4_n182, _add_2_root_add_136_4_n181, 
  _add_2_root_add_136_4_n180, _add_2_root_add_136_4_n179, _add_2_root_add_136_4_n178, _add_2_root_add_136_4_n177, _add_2_root_add_136_4_n176, _add_2_root_add_136_4_n175, _add_2_root_add_136_4_n174, _add_2_root_add_136_4_n173, _add_2_root_add_136_4_n172, _add_2_root_add_136_4_n171, _add_2_root_add_136_4_n170, _add_2_root_add_136_4_n169, _add_2_root_add_136_4_n168, _add_2_root_add_136_4_n167, _add_2_root_add_136_4_n166, _add_2_root_add_136_4_n165, _add_2_root_add_136_4_n164, _add_2_root_add_136_4_n163, _add_2_root_add_136_4_n162, _add_2_root_add_136_4_n161, _add_2_root_add_136_4_n160, _add_2_root_add_136_4_n159, _add_2_root_add_136_4_n158, _add_2_root_add_136_4_n157, _add_2_root_add_136_4_n156, _add_2_root_add_136_4_n155, _add_2_root_add_136_4_n154, _add_2_root_add_136_4_n153, _add_2_root_add_136_4_n152, _add_2_root_add_136_4_n151, _add_2_root_add_136_4_n150, _add_2_root_add_136_4_n149, _add_2_root_add_136_4_n148, _add_2_root_add_136_4_n147, _add_2_root_add_136_4_n146, _add_2_root_add_136_4_n145, _add_2_root_add_136_4_n144, _add_2_root_add_136_4_n143, _add_2_root_add_136_4_n142, _add_2_root_add_136_4_n141, _add_2_root_add_136_4_n140, _add_2_root_add_136_4_n139, _add_2_root_add_136_4_n138, _add_2_root_add_136_4_n137, _add_2_root_add_136_4_n136, _add_2_root_add_136_4_n135, _add_2_root_add_136_4_n134, _add_2_root_add_136_4_n133, _add_2_root_add_136_4_n132, _add_2_root_add_136_4_n131, 
  _add_2_root_add_136_4_n130, _add_2_root_add_136_4_n129, _add_2_root_add_136_4_n128, _add_2_root_add_136_4_n127, _add_2_root_add_136_4_n126, _add_2_root_add_136_4_n125, _add_2_root_add_136_4_n124, _add_2_root_add_136_4_n123, _add_2_root_add_136_4_n122, _add_2_root_add_136_4_n121, _add_2_root_add_136_4_n120, _add_2_root_add_136_4_n119, _add_2_root_add_136_4_n118, _add_2_root_add_136_4_n117, _add_2_root_add_136_4_n116, _add_2_root_add_136_4_n115, _add_2_root_add_136_4_n114, _add_2_root_add_136_4_n113, _add_2_root_add_136_4_n112, _add_2_root_add_136_4_n111, _add_2_root_add_136_4_n110, _add_2_root_add_136_4_n109, _add_2_root_add_136_4_n108, _add_2_root_add_136_4_n107, _add_2_root_add_136_4_n106, _add_2_root_add_136_4_n105, _add_2_root_add_136_4_n104, _add_2_root_add_136_4_n103, _add_2_root_add_136_4_n102, _add_2_root_add_136_4_n101, _add_2_root_add_136_4_n100, _add_2_root_add_136_4_n99, _add_2_root_add_136_4_n98, _add_2_root_add_136_4_n97, _add_2_root_add_136_4_n96, _add_2_root_add_136_4_n95, _add_2_root_add_136_4_n94, _add_2_root_add_136_4_n93, _add_2_root_add_136_4_n92, _add_2_root_add_136_4_n91, _add_2_root_add_136_4_n90, _add_2_root_add_136_4_n89, _add_2_root_add_136_4_n88, _add_2_root_add_136_4_n87, _add_2_root_add_136_4_n86, _add_2_root_add_136_4_n85, _add_2_root_add_136_4_n84, _add_2_root_add_136_4_n83, _add_2_root_add_136_4_n82, _add_2_root_add_136_4_n81, 
  _add_2_root_add_136_4_n80, _add_2_root_add_136_4_n79, _add_2_root_add_136_4_n78, _add_2_root_add_136_4_n77, _add_2_root_add_136_4_n76, _add_2_root_add_136_4_n75, _add_2_root_add_136_4_n74, _add_2_root_add_136_4_n73, _add_2_root_add_136_4_n72, _add_2_root_add_136_4_n71, _add_2_root_add_136_4_n70, _add_2_root_add_136_4_n69, _add_2_root_add_136_4_n68, _add_2_root_add_136_4_n67, _add_2_root_add_136_4_n66, _add_2_root_add_136_4_n65, _add_2_root_add_136_4_n64, _add_2_root_add_136_4_n63, _add_2_root_add_136_4_n62, _add_2_root_add_136_4_n61, _add_2_root_add_136_4_n60, _add_2_root_add_136_4_n59, _add_2_root_add_136_4_n58, _add_2_root_add_136_4_n57, _add_2_root_add_136_4_n56, _add_2_root_add_136_4_n55, _add_2_root_add_136_4_n54, _add_2_root_add_136_4_n53, _add_2_root_add_136_4_n52, _add_2_root_add_136_4_n51, _add_2_root_add_136_4_n50, _add_2_root_add_136_4_n49, _add_2_root_add_136_4_n48, _add_2_root_add_136_4_n47, _add_2_root_add_136_4_n46, _add_2_root_add_136_4_n45, _add_2_root_add_136_4_n44, _add_2_root_add_136_4_n43, _add_2_root_add_136_4_n42, _add_2_root_add_136_4_n41, _add_2_root_add_136_4_n40, _add_2_root_add_136_4_n39, _add_2_root_add_136_4_n38, _add_2_root_add_136_4_n37, _add_2_root_add_136_4_n36, _add_2_root_add_136_4_n35, _add_2_root_add_136_4_n34, _add_2_root_add_136_4_n33, _add_2_root_add_136_4_n32, _add_2_root_add_136_4_n31, 
  _add_2_root_add_136_4_n30, _add_2_root_add_136_4_n29, _add_2_root_add_136_4_n28, _add_2_root_add_136_4_n26, _add_2_root_add_136_4_n25, _add_2_root_add_136_4_n24, _add_2_root_add_136_4_n23, _add_2_root_add_136_4_n22, _add_2_root_add_136_4_n21, _add_2_root_add_136_4_n20, _add_2_root_add_136_4_n19, _add_2_root_add_136_4_n18, _add_2_root_add_136_4_n17, _add_2_root_add_136_4_n16, _add_2_root_add_136_4_n15, _add_2_root_add_136_4_n14, _add_2_root_add_136_4_n13, _add_2_root_add_136_4_n11, _add_2_root_add_136_4_n10, _add_2_root_add_136_4_n9, _add_2_root_add_136_4_n8, _add_2_root_add_136_4_n7, _add_2_root_add_136_4_n6, _add_2_root_add_136_4_n5, _add_2_root_add_136_4_n4, _add_2_root_add_136_4_n3, _add_2_root_add_136_4_n2, _add_2_root_add_136_4_n1, _add_514_n377, _add_514_n376, _add_514_n375, _add_514_n374, _add_514_n373, _add_514_n372, _add_514_n371, _add_514_n370, _add_514_n369, _add_514_n368, _add_514_n367, _add_514_n366, _add_514_n365, _add_514_n364, _add_514_n363, _add_514_n362, _add_514_n361, _add_514_n360, _add_514_n359, _add_514_n358, _add_514_n357, _add_514_n356, 
  _add_514_n355, _add_514_n354, _add_514_n353, _add_514_n352, _add_514_n351, _add_514_n350, _add_514_n349, _add_514_n348, _add_514_n347, _add_514_n346, _add_514_n345, _add_514_n344, _add_514_n343, _add_514_n342, _add_514_n341, _add_514_n340, _add_514_n339, _add_514_n338, _add_514_n337, _add_514_n336, _add_514_n335, _add_514_n334, _add_514_n333, _add_514_n332, _add_514_n331, _add_514_n330, _add_514_n329, _add_514_n328, _add_514_n327, _add_514_n326, _add_514_n325, _add_514_n324, _add_514_n323, _add_514_n322, _add_514_n321, _add_514_n320, _add_514_n319, _add_514_n318, _add_514_n317, _add_514_n316, _add_514_n315, _add_514_n314, _add_514_n313, _add_514_n312, _add_514_n311, _add_514_n310, _add_514_n309, _add_514_n308, _add_514_n307, _add_514_n306, 
  _add_514_n305, _add_514_n304, _add_514_n303, _add_514_n302, _add_514_n301, _add_514_n300, _add_514_n299, _add_514_n298, _add_514_n297, _add_514_n296, _add_514_n295, _add_514_n294, _add_514_n293, _add_514_n292, _add_514_n291, _add_514_n290, _add_514_n289, _add_514_n288, _add_514_n287, _add_514_n286, _add_514_n285, _add_514_n284, _add_514_n283, _add_514_n282, _add_514_n281, _add_514_n280, _add_514_n279, _add_514_n278, _add_514_n277, _add_514_n276, _add_514_n275, _add_514_n274, _add_514_n273, _add_514_n272, _add_514_n271, _add_514_n270, _add_514_n269, _add_514_n268, _add_514_n267, _add_514_n266, _add_514_n265, _add_514_n264, _add_514_n263, _add_514_n262, _add_514_n261, _add_514_n260, _add_514_n259, _add_514_n258, _add_514_n257, _add_514_n256, 
  _add_514_n255, _add_514_n254, _add_514_n253, _add_514_n252, _add_514_n251, _add_514_n250, _add_514_n249, _add_514_n248, _add_514_n247, _add_514_n246, _add_514_n245, _add_514_n244, _add_514_n243, _add_514_n242, _add_514_n241, _add_514_n240, _add_514_n239, _add_514_n238, _add_514_n237, _add_514_n236, _add_514_n235, _add_514_n234, _add_514_n233, _add_514_n232, _add_514_n231, _add_514_n230, _add_514_n229, _add_514_n228, _add_514_n227, _add_514_n226, _add_514_n225, _add_514_n224, _add_514_n223, _add_514_n222, _add_514_n221, _add_514_n220, _add_514_n219, _add_514_n218, _add_514_n217, _add_514_n216, _add_514_n215, _add_514_n214, _add_514_n213, _add_514_n212, _add_514_n211, _add_514_n210, _add_514_n209, _add_514_n208, _add_514_n207, _add_514_n206, 
  _add_514_n205, _add_514_n204, _add_514_n203, _add_514_n202, _add_514_n201, _add_514_n200, _add_514_n199, _add_514_n198, _add_514_n197, _add_514_n196, _add_514_n195, _add_514_n194, _add_514_n193, _add_514_n192, _add_514_n191, _add_514_n190, _add_514_n189, _add_514_n188, _add_514_n187, _add_514_n186, _add_514_n185, _add_514_n184, _add_514_n183, _add_514_n182, _add_514_n181, _add_514_n180, _add_514_n179, _add_514_n178, _add_514_n177, _add_514_n176, _add_514_n175, _add_514_n174, _add_514_n173, _add_514_n172, _add_514_n171, _add_514_n170, _add_514_n169, _add_514_n168, _add_514_n167, _add_514_n166, _add_514_n165, _add_514_n164, _add_514_n163, _add_514_n162, _add_514_n161, _add_514_n160, _add_514_n159, _add_514_n158, _add_514_n157, _add_514_n156, 
  _add_514_n155, _add_514_n154, _add_514_n153, _add_514_n152, _add_514_n151, _add_514_n150, _add_514_n149, _add_514_n148, _add_514_n147, _add_514_n146, _add_514_n145, _add_514_n144, _add_514_n143, _add_514_n142, _add_514_n141, _add_514_n140, _add_514_n139, _add_514_n138, _add_514_n137, _add_514_n136, _add_514_n135, _add_514_n134, _add_514_n133, _add_514_n132, _add_514_n131, _add_514_n130, _add_514_n129, _add_514_n128, _add_514_n127, _add_514_n126, _add_514_n125, _add_514_n124, _add_514_n123, _add_514_n122, _add_514_n121, _add_514_n120, _add_514_n119, _add_514_n118, _add_514_n117, _add_514_n116, _add_514_n115, _add_514_n114, _add_514_n113, _add_514_n112, _add_514_n111, _add_514_n110, _add_514_n109, _add_514_n108, _add_514_n107, _add_514_n106, 
  _add_514_n105, _add_514_n104, _add_514_n103, _add_514_n102, _add_514_n101, _add_514_n100, _add_514_n99, _add_514_n98, _add_514_n97, _add_514_n96, _add_514_n95, _add_514_n94, _add_514_n93, _add_514_n92, _add_514_n91, _add_514_n90, _add_514_n89, _add_514_n88, _add_514_n87, _add_514_n86, _add_514_n85, _add_514_n84, _add_514_n83, _add_514_n82, _add_514_n81, _add_514_n80, _add_514_n79, _add_514_n78, _add_514_n77, _add_514_n76, _add_514_n75, _add_514_n74, _add_514_n73, _add_514_n72, _add_514_n71, _add_514_n70, _add_514_n69, _add_514_n68, _add_514_n67, _add_514_n66, _add_514_n65, _add_514_n64, _add_514_n63, _add_514_n62, _add_514_n61, _add_514_n60, _add_514_n59, _add_514_n58, _add_514_n57, _add_514_n56, 
  _add_514_n55, _add_514_n54, _add_514_n53, _add_514_n52, _add_514_n51, _add_514_n50, _add_514_n49, _add_514_n48, _add_514_n47, _add_514_n46, _add_514_n45, _add_514_n44, _add_514_n43, _add_514_n42, _add_514_n41, _add_514_n40, _add_514_n39, _add_514_n38, _add_514_n37, _add_514_n36, _add_514_n35, _add_514_n34, _add_514_n33, _add_514_n32, _add_514_n31, _add_514_n30, _add_514_n29, _add_514_n28, _add_514_n27, _add_514_n26, _add_514_n25, _add_514_n24, _add_514_n23, _add_514_n22, _add_514_n21, _add_514_n20, _add_514_n19, _add_514_n18, _add_514_n17, _add_514_n16, _add_514_n15, _add_514_n14, _add_514_n12, _add_514_n11, _add_514_n10, _add_514_n9, _add_514_n8, _add_514_n7, _add_514_n6, _add_514_n5, 
  _add_514_n4, _add_514_n3, _add_514_n2, _add_514_n1, _add_513_n377, _add_513_n376, _add_513_n375, _add_513_n374, _add_513_n373, _add_513_n372, _add_513_n371, _add_513_n370, _add_513_n369, _add_513_n368, _add_513_n367, _add_513_n366, _add_513_n365, _add_513_n364, _add_513_n363, _add_513_n362, _add_513_n361, _add_513_n360, _add_513_n359, _add_513_n358, _add_513_n357, _add_513_n356, _add_513_n355, _add_513_n354, _add_513_n353, _add_513_n352, _add_513_n351, _add_513_n350, _add_513_n349, _add_513_n348, _add_513_n347, _add_513_n346, _add_513_n345, _add_513_n344, _add_513_n343, _add_513_n342, _add_513_n341, _add_513_n340, _add_513_n339, _add_513_n338, _add_513_n337, _add_513_n336, _add_513_n335, _add_513_n334, _add_513_n333, _add_513_n332, 
  _add_513_n331, _add_513_n330, _add_513_n329, _add_513_n328, _add_513_n327, _add_513_n326, _add_513_n325, _add_513_n324, _add_513_n323, _add_513_n322, _add_513_n321, _add_513_n320, _add_513_n319, _add_513_n318, _add_513_n317, _add_513_n316, _add_513_n315, _add_513_n314, _add_513_n313, _add_513_n312, _add_513_n311, _add_513_n310, _add_513_n309, _add_513_n308, _add_513_n307, _add_513_n306, _add_513_n305, _add_513_n304, _add_513_n303, _add_513_n302, _add_513_n301, _add_513_n300, _add_513_n299, _add_513_n298, _add_513_n297, _add_513_n296, _add_513_n295, _add_513_n294, _add_513_n293, _add_513_n292, _add_513_n291, _add_513_n290, _add_513_n289, _add_513_n288, _add_513_n287, _add_513_n286, _add_513_n285, _add_513_n284, _add_513_n283, _add_513_n282, 
  _add_513_n281, _add_513_n280, _add_513_n279, _add_513_n278, _add_513_n277, _add_513_n276, _add_513_n275, _add_513_n274, _add_513_n273, _add_513_n272, _add_513_n271, _add_513_n270, _add_513_n269, _add_513_n268, _add_513_n267, _add_513_n266, _add_513_n265, _add_513_n264, _add_513_n263, _add_513_n262, _add_513_n261, _add_513_n260, _add_513_n259, _add_513_n258, _add_513_n257, _add_513_n256, _add_513_n255, _add_513_n254, _add_513_n253, _add_513_n252, _add_513_n251, _add_513_n250, _add_513_n249, _add_513_n248, _add_513_n247, _add_513_n246, _add_513_n245, _add_513_n244, _add_513_n243, _add_513_n242, _add_513_n241, _add_513_n240, _add_513_n239, _add_513_n238, _add_513_n237, _add_513_n236, _add_513_n235, _add_513_n234, _add_513_n233, _add_513_n232, 
  _add_513_n231, _add_513_n230, _add_513_n229, _add_513_n228, _add_513_n227, _add_513_n226, _add_513_n225, _add_513_n224, _add_513_n223, _add_513_n222, _add_513_n221, _add_513_n220, _add_513_n219, _add_513_n218, _add_513_n217, _add_513_n216, _add_513_n215, _add_513_n214, _add_513_n213, _add_513_n212, _add_513_n211, _add_513_n210, _add_513_n209, _add_513_n208, _add_513_n207, _add_513_n206, _add_513_n205, _add_513_n204, _add_513_n203, _add_513_n202, _add_513_n201, _add_513_n200, _add_513_n199, _add_513_n198, _add_513_n197, _add_513_n196, _add_513_n195, _add_513_n194, _add_513_n193, _add_513_n192, _add_513_n191, _add_513_n190, _add_513_n189, _add_513_n188, _add_513_n187, _add_513_n186, _add_513_n185, _add_513_n184, _add_513_n183, _add_513_n182, 
  _add_513_n181, _add_513_n180, _add_513_n179, _add_513_n178, _add_513_n177, _add_513_n176, _add_513_n175, _add_513_n174, _add_513_n173, _add_513_n172, _add_513_n171, _add_513_n170, _add_513_n169, _add_513_n168, _add_513_n167, _add_513_n166, _add_513_n165, _add_513_n164, _add_513_n163, _add_513_n162, _add_513_n161, _add_513_n160, _add_513_n159, _add_513_n158, _add_513_n157, _add_513_n156, _add_513_n155, _add_513_n154, _add_513_n153, _add_513_n152, _add_513_n151, _add_513_n150, _add_513_n149, _add_513_n148, _add_513_n147, _add_513_n146, _add_513_n145, _add_513_n144, _add_513_n143, _add_513_n142, _add_513_n141, _add_513_n140, _add_513_n139, _add_513_n138, _add_513_n137, _add_513_n136, _add_513_n135, _add_513_n134, _add_513_n133, _add_513_n132, 
  _add_513_n131, _add_513_n130, _add_513_n129, _add_513_n128, _add_513_n127, _add_513_n126, _add_513_n125, _add_513_n124, _add_513_n123, _add_513_n122, _add_513_n121, _add_513_n120, _add_513_n119, _add_513_n118, _add_513_n117, _add_513_n116, _add_513_n115, _add_513_n114, _add_513_n113, _add_513_n112, _add_513_n111, _add_513_n110, _add_513_n109, _add_513_n108, _add_513_n107, _add_513_n106, _add_513_n105, _add_513_n104, _add_513_n103, _add_513_n102, _add_513_n101, _add_513_n100, _add_513_n99, _add_513_n98, _add_513_n97, _add_513_n96, _add_513_n95, _add_513_n94, _add_513_n93, _add_513_n92, _add_513_n91, _add_513_n90, _add_513_n89, _add_513_n88, _add_513_n87, _add_513_n86, _add_513_n85, _add_513_n84, _add_513_n83, _add_513_n82, 
  _add_513_n81, _add_513_n80, _add_513_n79, _add_513_n78, _add_513_n77, _add_513_n76, _add_513_n75, _add_513_n74, _add_513_n73, _add_513_n72, _add_513_n71, _add_513_n70, _add_513_n69, _add_513_n68, _add_513_n67, _add_513_n66, _add_513_n65, _add_513_n64, _add_513_n63, _add_513_n62, _add_513_n61, _add_513_n60, _add_513_n59, _add_513_n58, _add_513_n57, _add_513_n56, _add_513_n55, _add_513_n54, _add_513_n53, _add_513_n52, _add_513_n51, _add_513_n50, _add_513_n49, _add_513_n48, _add_513_n47, _add_513_n46, _add_513_n45, _add_513_n44, _add_513_n43, _add_513_n42, _add_513_n41, _add_513_n40, _add_513_n39, _add_513_n38, _add_513_n37, _add_513_n36, _add_513_n35, _add_513_n34, _add_513_n33, _add_513_n32, 
  _add_513_n31, _add_513_n30, _add_513_n29, _add_513_n28, _add_513_n27, _add_513_n26, _add_513_n25, _add_513_n24, _add_513_n23, _add_513_n22, _add_513_n21, _add_513_n20, _add_513_n19, _add_513_n18, _add_513_n17, _add_513_n16, _add_513_n15, _add_513_n14, _add_513_n13, _add_513_n12, _add_513_n11, _add_513_n10, _add_513_n8, _add_513_n7, _add_513_n6, _add_513_n5, _add_513_n4, _add_513_n3, _add_513_n2, _add_513_n1, _add_516_n390, _add_516_n389, _add_516_n388, _add_516_n387, _add_516_n386, _add_516_n385, _add_516_n384, _add_516_n383, _add_516_n382, _add_516_n381, _add_516_n380, _add_516_n379, _add_516_n378, _add_516_n377, _add_516_n376, _add_516_n375, _add_516_n374, _add_516_n373, _add_516_n372, _add_516_n371, 
  _add_516_n370, _add_516_n369, _add_516_n368, _add_516_n367, _add_516_n366, _add_516_n365, _add_516_n364, _add_516_n363, _add_516_n362, _add_516_n361, _add_516_n360, _add_516_n359, _add_516_n358, _add_516_n357, _add_516_n356, _add_516_n355, _add_516_n354, _add_516_n353, _add_516_n352, _add_516_n351, _add_516_n350, _add_516_n349, _add_516_n348, _add_516_n347, _add_516_n346, _add_516_n345, _add_516_n344, _add_516_n343, _add_516_n342, _add_516_n341, _add_516_n340, _add_516_n339, _add_516_n338, _add_516_n337, _add_516_n336, _add_516_n335, _add_516_n334, _add_516_n333, _add_516_n332, _add_516_n331, _add_516_n330, _add_516_n329, _add_516_n328, _add_516_n327, _add_516_n326, _add_516_n325, _add_516_n324, _add_516_n323, _add_516_n322, _add_516_n321, 
  _add_516_n320, _add_516_n319, _add_516_n318, _add_516_n317, _add_516_n316, _add_516_n315, _add_516_n314, _add_516_n313, _add_516_n312, _add_516_n311, _add_516_n310, _add_516_n309, _add_516_n308, _add_516_n307, _add_516_n306, _add_516_n305, _add_516_n304, _add_516_n303, _add_516_n302, _add_516_n301, _add_516_n300, _add_516_n299, _add_516_n298, _add_516_n297, _add_516_n296, _add_516_n295, _add_516_n294, _add_516_n293, _add_516_n292, _add_516_n291, _add_516_n290, _add_516_n289, _add_516_n288, _add_516_n287, _add_516_n286, _add_516_n285, _add_516_n284, _add_516_n283, _add_516_n282, _add_516_n281, _add_516_n280, _add_516_n279, _add_516_n278, _add_516_n277, _add_516_n276, _add_516_n275, _add_516_n274, _add_516_n273, _add_516_n272, _add_516_n271, 
  _add_516_n270, _add_516_n269, _add_516_n268, _add_516_n267, _add_516_n266, _add_516_n265, _add_516_n264, _add_516_n263, _add_516_n262, _add_516_n261, _add_516_n260, _add_516_n259, _add_516_n258, _add_516_n257, _add_516_n256, _add_516_n255, _add_516_n254, _add_516_n253, _add_516_n252, _add_516_n251, _add_516_n250, _add_516_n249, _add_516_n248, _add_516_n247, _add_516_n246, _add_516_n245, _add_516_n244, _add_516_n243, _add_516_n242, _add_516_n241, _add_516_n240, _add_516_n239, _add_516_n238, _add_516_n237, _add_516_n236, _add_516_n235, _add_516_n234, _add_516_n233, _add_516_n232, _add_516_n231, _add_516_n230, _add_516_n229, _add_516_n228, _add_516_n227, _add_516_n226, _add_516_n225, _add_516_n224, _add_516_n223, _add_516_n222, _add_516_n221, 
  _add_516_n220, _add_516_n219, _add_516_n218, _add_516_n217, _add_516_n216, _add_516_n215, _add_516_n214, _add_516_n213, _add_516_n212, _add_516_n211, _add_516_n210, _add_516_n209, _add_516_n208, _add_516_n207, _add_516_n206, _add_516_n205, _add_516_n204, _add_516_n203, _add_516_n202, _add_516_n201, _add_516_n200, _add_516_n199, _add_516_n198, _add_516_n197, _add_516_n196, _add_516_n195, _add_516_n194, _add_516_n193, _add_516_n192, _add_516_n191, _add_516_n190, _add_516_n189, _add_516_n188, _add_516_n187, _add_516_n186, _add_516_n185, _add_516_n184, _add_516_n183, _add_516_n182, _add_516_n181, _add_516_n180, _add_516_n179, _add_516_n178, _add_516_n177, _add_516_n176, _add_516_n175, _add_516_n174, _add_516_n173, _add_516_n172, _add_516_n171, 
  _add_516_n170, _add_516_n169, _add_516_n168, _add_516_n167, _add_516_n166, _add_516_n165, _add_516_n164, _add_516_n163, _add_516_n162, _add_516_n161, _add_516_n160, _add_516_n159, _add_516_n158, _add_516_n157, _add_516_n156, _add_516_n155, _add_516_n154, _add_516_n153, _add_516_n152, _add_516_n151, _add_516_n150, _add_516_n149, _add_516_n148, _add_516_n147, _add_516_n146, _add_516_n145, _add_516_n144, _add_516_n143, _add_516_n142, _add_516_n141, _add_516_n140, _add_516_n139, _add_516_n138, _add_516_n137, _add_516_n136, _add_516_n135, _add_516_n134, _add_516_n133, _add_516_n132, _add_516_n131, _add_516_n130, _add_516_n129, _add_516_n128, _add_516_n127, _add_516_n126, _add_516_n125, _add_516_n124, _add_516_n123, _add_516_n122, _add_516_n121, 
  _add_516_n120, _add_516_n119, _add_516_n118, _add_516_n117, _add_516_n116, _add_516_n115, _add_516_n114, _add_516_n113, _add_516_n112, _add_516_n111, _add_516_n110, _add_516_n109, _add_516_n108, _add_516_n107, _add_516_n106, _add_516_n105, _add_516_n104, _add_516_n103, _add_516_n102, _add_516_n101, _add_516_n100, _add_516_n99, _add_516_n98, _add_516_n97, _add_516_n96, _add_516_n95, _add_516_n94, _add_516_n93, _add_516_n92, _add_516_n91, _add_516_n90, _add_516_n89, _add_516_n88, _add_516_n87, _add_516_n86, _add_516_n85, _add_516_n84, _add_516_n83, _add_516_n82, _add_516_n81, _add_516_n80, _add_516_n79, _add_516_n78, _add_516_n77, _add_516_n76, _add_516_n75, _add_516_n74, _add_516_n73, _add_516_n72, _add_516_n71, 
  _add_516_n70, _add_516_n69, _add_516_n68, _add_516_n67, _add_516_n66, _add_516_n65, _add_516_n64, _add_516_n63, _add_516_n62, _add_516_n61, _add_516_n60, _add_516_n59, _add_516_n58, _add_516_n57, _add_516_n56, _add_516_n55, _add_516_n54, _add_516_n53, _add_516_n52, _add_516_n51, _add_516_n50, _add_516_n49, _add_516_n48, _add_516_n47, _add_516_n46, _add_516_n45, _add_516_n44, _add_516_n43, _add_516_n42, _add_516_n41, _add_516_n40, _add_516_n39, _add_516_n38, _add_516_n37, _add_516_n36, _add_516_n35, _add_516_n34, _add_516_n33, _add_516_n32, _add_516_n31, _add_516_n30, _add_516_n29, _add_516_n28, _add_516_n27, _add_516_n26, _add_516_n25, _add_516_n24, _add_516_n23, _add_516_n22, _add_516_n21, 
  _add_516_n20, _add_516_n19, _add_516_n18, _add_516_n17, _add_516_n16, _add_516_n15, _add_516_n14, _add_516_n13, _add_516_n12, _add_516_n11, _add_516_n10, _add_516_n9, _add_516_n8, _add_516_n7, _add_516_n6, _add_516_n5, _add_516_n4, _add_516_n3, _add_516_n2, _add_516_n1, _add_515_n375, _add_515_n374, _add_515_n373, _add_515_n372, _add_515_n371, _add_515_n370, _add_515_n369, _add_515_n368, _add_515_n367, _add_515_n366, _add_515_n365, _add_515_n364, _add_515_n363, _add_515_n362, _add_515_n361, _add_515_n360, _add_515_n359, _add_515_n358, _add_515_n357, _add_515_n356, _add_515_n355, _add_515_n354, _add_515_n353, _add_515_n352, _add_515_n351, _add_515_n350, _add_515_n349, _add_515_n348, _add_515_n347, _add_515_n346, 
  _add_515_n345, _add_515_n344, _add_515_n343, _add_515_n342, _add_515_n341, _add_515_n340, _add_515_n339, _add_515_n338, _add_515_n337, _add_515_n336, _add_515_n335, _add_515_n334, _add_515_n333, _add_515_n332, _add_515_n331, _add_515_n330, _add_515_n329, _add_515_n328, _add_515_n327, _add_515_n326, _add_515_n325, _add_515_n324, _add_515_n323, _add_515_n322, _add_515_n321, _add_515_n320, _add_515_n319, _add_515_n318, _add_515_n317, _add_515_n316, _add_515_n315, _add_515_n314, _add_515_n313, _add_515_n312, _add_515_n311, _add_515_n310, _add_515_n309, _add_515_n308, _add_515_n307, _add_515_n306, _add_515_n305, _add_515_n304, _add_515_n303, _add_515_n302, _add_515_n301, _add_515_n300, _add_515_n299, _add_515_n298, _add_515_n297, _add_515_n296, 
  _add_515_n295, _add_515_n294, _add_515_n293, _add_515_n292, _add_515_n291, _add_515_n290, _add_515_n289, _add_515_n288, _add_515_n287, _add_515_n286, _add_515_n285, _add_515_n284, _add_515_n283, _add_515_n282, _add_515_n281, _add_515_n280, _add_515_n279, _add_515_n278, _add_515_n277, _add_515_n276, _add_515_n275, _add_515_n274, _add_515_n273, _add_515_n272, _add_515_n271, _add_515_n270, _add_515_n269, _add_515_n268, _add_515_n267, _add_515_n266, _add_515_n265, _add_515_n264, _add_515_n263, _add_515_n262, _add_515_n261, _add_515_n260, _add_515_n259, _add_515_n258, _add_515_n257, _add_515_n256, _add_515_n255, _add_515_n254, _add_515_n253, _add_515_n252, _add_515_n251, _add_515_n250, _add_515_n249, _add_515_n248, _add_515_n247, _add_515_n246, 
  _add_515_n245, _add_515_n244, _add_515_n243, _add_515_n242, _add_515_n241, _add_515_n240, _add_515_n239, _add_515_n238, _add_515_n237, _add_515_n236, _add_515_n235, _add_515_n234, _add_515_n233, _add_515_n232, _add_515_n231, _add_515_n230, _add_515_n229, _add_515_n228, _add_515_n227, _add_515_n226, _add_515_n225, _add_515_n224, _add_515_n223, _add_515_n222, _add_515_n221, _add_515_n220, _add_515_n219, _add_515_n218, _add_515_n217, _add_515_n216, _add_515_n215, _add_515_n214, _add_515_n213, _add_515_n212, _add_515_n211, _add_515_n210, _add_515_n209, _add_515_n208, _add_515_n207, _add_515_n206, _add_515_n205, _add_515_n204, _add_515_n203, _add_515_n202, _add_515_n201, _add_515_n200, _add_515_n199, _add_515_n198, _add_515_n197, _add_515_n196, 
  _add_515_n195, _add_515_n194, _add_515_n193, _add_515_n192, _add_515_n191, _add_515_n190, _add_515_n189, _add_515_n188, _add_515_n187, _add_515_n186, _add_515_n185, _add_515_n184, _add_515_n183, _add_515_n182, _add_515_n181, _add_515_n180, _add_515_n179, _add_515_n178, _add_515_n177, _add_515_n176, _add_515_n175, _add_515_n174, _add_515_n173, _add_515_n172, _add_515_n171, _add_515_n170, _add_515_n169, _add_515_n168, _add_515_n167, _add_515_n166, _add_515_n165, _add_515_n164, _add_515_n163, _add_515_n162, _add_515_n161, _add_515_n160, _add_515_n159, _add_515_n158, _add_515_n157, _add_515_n156, _add_515_n155, _add_515_n154, _add_515_n153, _add_515_n152, _add_515_n151, _add_515_n150, _add_515_n149, _add_515_n148, _add_515_n147, _add_515_n146, 
  _add_515_n145, _add_515_n144, _add_515_n143, _add_515_n142, _add_515_n141, _add_515_n140, _add_515_n139, _add_515_n138, _add_515_n137, _add_515_n136, _add_515_n135, _add_515_n134, _add_515_n133, _add_515_n132, _add_515_n131, _add_515_n130, _add_515_n129, _add_515_n128, _add_515_n127, _add_515_n126, _add_515_n125, _add_515_n124, _add_515_n123, _add_515_n122, _add_515_n121, _add_515_n120, _add_515_n119, _add_515_n118, _add_515_n117, _add_515_n116, _add_515_n115, _add_515_n114, _add_515_n113, _add_515_n112, _add_515_n111, _add_515_n110, _add_515_n109, _add_515_n108, _add_515_n107, _add_515_n106, _add_515_n105, _add_515_n104, _add_515_n103, _add_515_n102, _add_515_n101, _add_515_n100, _add_515_n99, _add_515_n98, _add_515_n97, _add_515_n96, 
  _add_515_n95, _add_515_n94, _add_515_n93, _add_515_n92, _add_515_n91, _add_515_n90, _add_515_n89, _add_515_n88, _add_515_n87, _add_515_n86, _add_515_n85, _add_515_n84, _add_515_n83, _add_515_n82, _add_515_n81, _add_515_n80, _add_515_n79, _add_515_n78, _add_515_n77, _add_515_n76, _add_515_n75, _add_515_n74, _add_515_n73, _add_515_n72, _add_515_n71, _add_515_n70, _add_515_n69, _add_515_n68, _add_515_n67, _add_515_n66, _add_515_n65, _add_515_n64, _add_515_n63, _add_515_n62, _add_515_n61, _add_515_n60, _add_515_n59, _add_515_n58, _add_515_n57, _add_515_n56, _add_515_n55, _add_515_n54, _add_515_n53, _add_515_n52, _add_515_n51, _add_515_n50, _add_515_n49, _add_515_n48, _add_515_n47, _add_515_n46, 
  _add_515_n45, _add_515_n44, _add_515_n43, _add_515_n42, _add_515_n41, _add_515_n40, _add_515_n39, _add_515_n38, _add_515_n37, _add_515_n36, _add_515_n35, _add_515_n34, _add_515_n33, _add_515_n32, _add_515_n31, _add_515_n30, _add_515_n29, _add_515_n28, _add_515_n27, _add_515_n26, _add_515_n25, _add_515_n24, _add_515_n23, _add_515_n22, _add_515_n21, _add_515_n20, _add_515_n19, _add_515_n18, _add_515_n17, _add_515_n16, _add_515_n14, _add_515_n13, _add_515_n12, _add_515_n11, _add_515_n10, _add_515_n9, _add_515_n8, _add_515_n7, _add_515_n6, _add_515_n5, _add_515_n4, _add_515_n3, _add_515_n2, _add_515_n1, _add_1_root_add_136_4_n411, _add_1_root_add_136_4_n410, _add_1_root_add_136_4_n409, _add_1_root_add_136_4_n408, _add_1_root_add_136_4_n407, _add_1_root_add_136_4_n406, 
  _add_1_root_add_136_4_n405, _add_1_root_add_136_4_n404, _add_1_root_add_136_4_n403, _add_1_root_add_136_4_n402, _add_1_root_add_136_4_n401, _add_1_root_add_136_4_n400, _add_1_root_add_136_4_n399, _add_1_root_add_136_4_n398, _add_1_root_add_136_4_n397, _add_1_root_add_136_4_n396, _add_1_root_add_136_4_n395, _add_1_root_add_136_4_n394, _add_1_root_add_136_4_n393, _add_1_root_add_136_4_n392, _add_1_root_add_136_4_n391, _add_1_root_add_136_4_n390, _add_1_root_add_136_4_n389, _add_1_root_add_136_4_n388, _add_1_root_add_136_4_n387, _add_1_root_add_136_4_n386, _add_1_root_add_136_4_n385, _add_1_root_add_136_4_n384, _add_1_root_add_136_4_n383, _add_1_root_add_136_4_n382, _add_1_root_add_136_4_n381, _add_1_root_add_136_4_n380, _add_1_root_add_136_4_n379, _add_1_root_add_136_4_n378, _add_1_root_add_136_4_n377, _add_1_root_add_136_4_n376, _add_1_root_add_136_4_n375, _add_1_root_add_136_4_n374, _add_1_root_add_136_4_n373, _add_1_root_add_136_4_n372, _add_1_root_add_136_4_n371, _add_1_root_add_136_4_n370, _add_1_root_add_136_4_n369, _add_1_root_add_136_4_n368, _add_1_root_add_136_4_n367, _add_1_root_add_136_4_n366, _add_1_root_add_136_4_n365, _add_1_root_add_136_4_n364, _add_1_root_add_136_4_n363, _add_1_root_add_136_4_n362, _add_1_root_add_136_4_n361, _add_1_root_add_136_4_n360, _add_1_root_add_136_4_n359, _add_1_root_add_136_4_n358, _add_1_root_add_136_4_n357, _add_1_root_add_136_4_n356, 
  _add_1_root_add_136_4_n355, _add_1_root_add_136_4_n354, _add_1_root_add_136_4_n353, _add_1_root_add_136_4_n352, _add_1_root_add_136_4_n351, _add_1_root_add_136_4_n350, _add_1_root_add_136_4_n349, _add_1_root_add_136_4_n348, _add_1_root_add_136_4_n347, _add_1_root_add_136_4_n346, _add_1_root_add_136_4_n345, _add_1_root_add_136_4_n344, _add_1_root_add_136_4_n343, _add_1_root_add_136_4_n342, _add_1_root_add_136_4_n341, _add_1_root_add_136_4_n340, _add_1_root_add_136_4_n339, _add_1_root_add_136_4_n338, _add_1_root_add_136_4_n337, _add_1_root_add_136_4_n336, _add_1_root_add_136_4_n335, _add_1_root_add_136_4_n334, _add_1_root_add_136_4_n333, _add_1_root_add_136_4_n332, _add_1_root_add_136_4_n331, _add_1_root_add_136_4_n330, _add_1_root_add_136_4_n329, _add_1_root_add_136_4_n328, _add_1_root_add_136_4_n327, _add_1_root_add_136_4_n326, _add_1_root_add_136_4_n325, _add_1_root_add_136_4_n324, _add_1_root_add_136_4_n323, _add_1_root_add_136_4_n322, _add_1_root_add_136_4_n321, _add_1_root_add_136_4_n320, _add_1_root_add_136_4_n319, _add_1_root_add_136_4_n318, _add_1_root_add_136_4_n317, _add_1_root_add_136_4_n316, _add_1_root_add_136_4_n315, _add_1_root_add_136_4_n314, _add_1_root_add_136_4_n313, _add_1_root_add_136_4_n312, _add_1_root_add_136_4_n311, _add_1_root_add_136_4_n310, _add_1_root_add_136_4_n309, _add_1_root_add_136_4_n308, _add_1_root_add_136_4_n307, _add_1_root_add_136_4_n306, 
  _add_1_root_add_136_4_n305, _add_1_root_add_136_4_n304, _add_1_root_add_136_4_n303, _add_1_root_add_136_4_n302, _add_1_root_add_136_4_n301, _add_1_root_add_136_4_n300, _add_1_root_add_136_4_n299, _add_1_root_add_136_4_n298, _add_1_root_add_136_4_n297, _add_1_root_add_136_4_n296, _add_1_root_add_136_4_n295, _add_1_root_add_136_4_n294, _add_1_root_add_136_4_n293, _add_1_root_add_136_4_n292, _add_1_root_add_136_4_n291, _add_1_root_add_136_4_n290, _add_1_root_add_136_4_n289, _add_1_root_add_136_4_n288, _add_1_root_add_136_4_n287, _add_1_root_add_136_4_n286, _add_1_root_add_136_4_n285, _add_1_root_add_136_4_n284, _add_1_root_add_136_4_n283, _add_1_root_add_136_4_n282, _add_1_root_add_136_4_n281, _add_1_root_add_136_4_n280, _add_1_root_add_136_4_n279, _add_1_root_add_136_4_n278, _add_1_root_add_136_4_n277, _add_1_root_add_136_4_n276, _add_1_root_add_136_4_n275, _add_1_root_add_136_4_n274, _add_1_root_add_136_4_n273, _add_1_root_add_136_4_n272, _add_1_root_add_136_4_n271, _add_1_root_add_136_4_n270, _add_1_root_add_136_4_n269, _add_1_root_add_136_4_n268, _add_1_root_add_136_4_n267, _add_1_root_add_136_4_n266, _add_1_root_add_136_4_n265, _add_1_root_add_136_4_n264, _add_1_root_add_136_4_n263, _add_1_root_add_136_4_n262, _add_1_root_add_136_4_n261, _add_1_root_add_136_4_n260, _add_1_root_add_136_4_n259, _add_1_root_add_136_4_n258, _add_1_root_add_136_4_n257, _add_1_root_add_136_4_n256, 
  _add_1_root_add_136_4_n255, _add_1_root_add_136_4_n254, _add_1_root_add_136_4_n253, _add_1_root_add_136_4_n252, _add_1_root_add_136_4_n251, _add_1_root_add_136_4_n250, _add_1_root_add_136_4_n249, _add_1_root_add_136_4_n248, _add_1_root_add_136_4_n247, _add_1_root_add_136_4_n246, _add_1_root_add_136_4_n245, _add_1_root_add_136_4_n244, _add_1_root_add_136_4_n243, _add_1_root_add_136_4_n242, _add_1_root_add_136_4_n241, _add_1_root_add_136_4_n240, _add_1_root_add_136_4_n239, _add_1_root_add_136_4_n238, _add_1_root_add_136_4_n237, _add_1_root_add_136_4_n236, _add_1_root_add_136_4_n235, _add_1_root_add_136_4_n234, _add_1_root_add_136_4_n233, _add_1_root_add_136_4_n232, _add_1_root_add_136_4_n231, _add_1_root_add_136_4_n230, _add_1_root_add_136_4_n229, _add_1_root_add_136_4_n228, _add_1_root_add_136_4_n227, _add_1_root_add_136_4_n226, _add_1_root_add_136_4_n225, _add_1_root_add_136_4_n224, _add_1_root_add_136_4_n223, _add_1_root_add_136_4_n222, _add_1_root_add_136_4_n221, _add_1_root_add_136_4_n220, _add_1_root_add_136_4_n219, _add_1_root_add_136_4_n218, _add_1_root_add_136_4_n217, _add_1_root_add_136_4_n216, _add_1_root_add_136_4_n215, _add_1_root_add_136_4_n214, _add_1_root_add_136_4_n213, _add_1_root_add_136_4_n212, _add_1_root_add_136_4_n211, _add_1_root_add_136_4_n210, _add_1_root_add_136_4_n209, _add_1_root_add_136_4_n208, _add_1_root_add_136_4_n207, _add_1_root_add_136_4_n206, 
  _add_1_root_add_136_4_n205, _add_1_root_add_136_4_n204, _add_1_root_add_136_4_n203, _add_1_root_add_136_4_n202, _add_1_root_add_136_4_n201, _add_1_root_add_136_4_n200, _add_1_root_add_136_4_n199, _add_1_root_add_136_4_n198, _add_1_root_add_136_4_n197, _add_1_root_add_136_4_n196, _add_1_root_add_136_4_n195, _add_1_root_add_136_4_n194, _add_1_root_add_136_4_n193, _add_1_root_add_136_4_n192, _add_1_root_add_136_4_n191, _add_1_root_add_136_4_n190, _add_1_root_add_136_4_n189, _add_1_root_add_136_4_n188, _add_1_root_add_136_4_n187, _add_1_root_add_136_4_n186, _add_1_root_add_136_4_n185, _add_1_root_add_136_4_n184, _add_1_root_add_136_4_n183, _add_1_root_add_136_4_n182, _add_1_root_add_136_4_n181, _add_1_root_add_136_4_n180, _add_1_root_add_136_4_n179, _add_1_root_add_136_4_n178, _add_1_root_add_136_4_n177, _add_1_root_add_136_4_n176, _add_1_root_add_136_4_n175, _add_1_root_add_136_4_n174, _add_1_root_add_136_4_n173, _add_1_root_add_136_4_n172, _add_1_root_add_136_4_n171, _add_1_root_add_136_4_n170, _add_1_root_add_136_4_n169, _add_1_root_add_136_4_n168, _add_1_root_add_136_4_n167, _add_1_root_add_136_4_n166, _add_1_root_add_136_4_n165, _add_1_root_add_136_4_n164, _add_1_root_add_136_4_n163, _add_1_root_add_136_4_n162, _add_1_root_add_136_4_n161, _add_1_root_add_136_4_n160, _add_1_root_add_136_4_n159, _add_1_root_add_136_4_n158, _add_1_root_add_136_4_n157, _add_1_root_add_136_4_n156, 
  _add_1_root_add_136_4_n155, _add_1_root_add_136_4_n154, _add_1_root_add_136_4_n153, _add_1_root_add_136_4_n152, _add_1_root_add_136_4_n151, _add_1_root_add_136_4_n150, _add_1_root_add_136_4_n149, _add_1_root_add_136_4_n148, _add_1_root_add_136_4_n147, _add_1_root_add_136_4_n146, _add_1_root_add_136_4_n145, _add_1_root_add_136_4_n144, _add_1_root_add_136_4_n143, _add_1_root_add_136_4_n142, _add_1_root_add_136_4_n141, _add_1_root_add_136_4_n140, _add_1_root_add_136_4_n139, _add_1_root_add_136_4_n138, _add_1_root_add_136_4_n137, _add_1_root_add_136_4_n136, _add_1_root_add_136_4_n135, _add_1_root_add_136_4_n134, _add_1_root_add_136_4_n133, _add_1_root_add_136_4_n132, _add_1_root_add_136_4_n131, _add_1_root_add_136_4_n130, _add_1_root_add_136_4_n129, _add_1_root_add_136_4_n128, _add_1_root_add_136_4_n127, _add_1_root_add_136_4_n126, _add_1_root_add_136_4_n125, _add_1_root_add_136_4_n124, _add_1_root_add_136_4_n123, _add_1_root_add_136_4_n122, _add_1_root_add_136_4_n121, _add_1_root_add_136_4_n120, _add_1_root_add_136_4_n119, _add_1_root_add_136_4_n118, _add_1_root_add_136_4_n117, _add_1_root_add_136_4_n116, _add_1_root_add_136_4_n115, _add_1_root_add_136_4_n114, _add_1_root_add_136_4_n113, _add_1_root_add_136_4_n112, _add_1_root_add_136_4_n111, _add_1_root_add_136_4_n110, _add_1_root_add_136_4_n109, _add_1_root_add_136_4_n108, _add_1_root_add_136_4_n107, _add_1_root_add_136_4_n106, 
  _add_1_root_add_136_4_n105, _add_1_root_add_136_4_n104, _add_1_root_add_136_4_n103, _add_1_root_add_136_4_n102, _add_1_root_add_136_4_n101, _add_1_root_add_136_4_n100, _add_1_root_add_136_4_n99, _add_1_root_add_136_4_n98, _add_1_root_add_136_4_n97, _add_1_root_add_136_4_n96, _add_1_root_add_136_4_n95, _add_1_root_add_136_4_n94, _add_1_root_add_136_4_n93, _add_1_root_add_136_4_n92, _add_1_root_add_136_4_n91, _add_1_root_add_136_4_n90, _add_1_root_add_136_4_n89, _add_1_root_add_136_4_n88, _add_1_root_add_136_4_n87, _add_1_root_add_136_4_n86, _add_1_root_add_136_4_n85, _add_1_root_add_136_4_n84, _add_1_root_add_136_4_n83, _add_1_root_add_136_4_n82, _add_1_root_add_136_4_n81, _add_1_root_add_136_4_n80, _add_1_root_add_136_4_n79, _add_1_root_add_136_4_n78, _add_1_root_add_136_4_n77, _add_1_root_add_136_4_n76, _add_1_root_add_136_4_n75, _add_1_root_add_136_4_n74, _add_1_root_add_136_4_n73, _add_1_root_add_136_4_n72, _add_1_root_add_136_4_n71, _add_1_root_add_136_4_n70, _add_1_root_add_136_4_n69, _add_1_root_add_136_4_n68, _add_1_root_add_136_4_n67, _add_1_root_add_136_4_n66, _add_1_root_add_136_4_n65, _add_1_root_add_136_4_n64, _add_1_root_add_136_4_n62, _add_1_root_add_136_4_n60, _add_1_root_add_136_4_n59, _add_1_root_add_136_4_n58, _add_1_root_add_136_4_n57, _add_1_root_add_136_4_n56, _add_1_root_add_136_4_n54, _add_1_root_add_136_4_n53, 
  _add_1_root_add_136_4_n52, _add_1_root_add_136_4_n51, _add_1_root_add_136_4_n50, _add_1_root_add_136_4_n49, _add_1_root_add_136_4_n48, _add_1_root_add_136_4_n47, _add_1_root_add_136_4_n46, _add_1_root_add_136_4_n45, _add_1_root_add_136_4_n44, _add_1_root_add_136_4_n43, _add_1_root_add_136_4_n42, _add_1_root_add_136_4_n41, _add_1_root_add_136_4_n40, _add_1_root_add_136_4_n39, _add_1_root_add_136_4_n38, _add_1_root_add_136_4_n37, _add_1_root_add_136_4_n36, _add_1_root_add_136_4_n35, _add_1_root_add_136_4_n34, _add_1_root_add_136_4_n33, _add_1_root_add_136_4_n32, _add_1_root_add_136_4_n31, _add_1_root_add_136_4_n30, _add_1_root_add_136_4_n29, _add_1_root_add_136_4_n28, _add_1_root_add_136_4_n27, _add_1_root_add_136_4_n26, _add_1_root_add_136_4_n25, _add_1_root_add_136_4_n24, _add_1_root_add_136_4_n23, _add_1_root_add_136_4_n22, _add_1_root_add_136_4_n21, _add_1_root_add_136_4_n20, _add_1_root_add_136_4_n19, _add_1_root_add_136_4_n18, _add_1_root_add_136_4_n17, _add_1_root_add_136_4_n16, _add_1_root_add_136_4_n15, _add_1_root_add_136_4_n14, _add_1_root_add_136_4_n13, _add_1_root_add_136_4_n12, _add_1_root_add_136_4_n11, _add_1_root_add_136_4_n10, _add_1_root_add_136_4_n9, _add_1_root_add_136_4_n8, _add_1_root_add_136_4_n7, _add_1_root_add_136_4_n6, _add_1_root_add_136_4_n5, _add_1_root_add_136_4_n4, _add_1_root_add_136_4_n3, 
  _add_1_root_add_136_4_n2, _add_1_root_add_136_4_n1, _add_512_n426, _add_512_n425, _add_512_n424, _add_512_n423, _add_512_n422, _add_512_n421, _add_512_n420, _add_512_n419, _add_512_n418, _add_512_n417, _add_512_n416, _add_512_n415, _add_512_n414, _add_512_n413, _add_512_n412, _add_512_n411, _add_512_n410, _add_512_n409, _add_512_n408, _add_512_n407, _add_512_n406, _add_512_n405, _add_512_n404, _add_512_n403, _add_512_n402, _add_512_n401, _add_512_n400, _add_512_n399, _add_512_n398, _add_512_n397, _add_512_n396, _add_512_n395, _add_512_n394, _add_512_n393, _add_512_n392, _add_512_n391, _add_512_n390, _add_512_n389, _add_512_n388, _add_512_n387, _add_512_n386, _add_512_n385, _add_512_n384, _add_512_n383, _add_512_n382, _add_512_n381, _add_512_n380, _add_512_n379, 
  _add_512_n378, _add_512_n377, _add_512_n376, _add_512_n375, _add_512_n374, _add_512_n373, _add_512_n372, _add_512_n371, _add_512_n370, _add_512_n369, _add_512_n368, _add_512_n367, _add_512_n366, _add_512_n365, _add_512_n364, _add_512_n363, _add_512_n362, _add_512_n361, _add_512_n360, _add_512_n359, _add_512_n358, _add_512_n357, _add_512_n356, _add_512_n355, _add_512_n354, _add_512_n353, _add_512_n352, _add_512_n351, _add_512_n350, _add_512_n349, _add_512_n348, _add_512_n347, _add_512_n346, _add_512_n345, _add_512_n344, _add_512_n343, _add_512_n342, _add_512_n341, _add_512_n340, _add_512_n339, _add_512_n338, _add_512_n337, _add_512_n336, _add_512_n335, _add_512_n334, _add_512_n333, _add_512_n332, _add_512_n331, _add_512_n330, _add_512_n329, 
  _add_512_n328, _add_512_n327, _add_512_n326, _add_512_n325, _add_512_n324, _add_512_n323, _add_512_n322, _add_512_n321, _add_512_n320, _add_512_n319, _add_512_n318, _add_512_n317, _add_512_n316, _add_512_n315, _add_512_n314, _add_512_n313, _add_512_n312, _add_512_n311, _add_512_n310, _add_512_n309, _add_512_n308, _add_512_n307, _add_512_n306, _add_512_n305, _add_512_n304, _add_512_n303, _add_512_n302, _add_512_n301, _add_512_n300, _add_512_n299, _add_512_n298, _add_512_n297, _add_512_n296, _add_512_n295, _add_512_n294, _add_512_n293, _add_512_n292, _add_512_n291, _add_512_n290, _add_512_n289, _add_512_n288, _add_512_n287, _add_512_n286, _add_512_n285, _add_512_n284, _add_512_n283, _add_512_n282, _add_512_n281, _add_512_n280, _add_512_n279, 
  _add_512_n278, _add_512_n277, _add_512_n276, _add_512_n275, _add_512_n274, _add_512_n273, _add_512_n272, _add_512_n271, _add_512_n270, _add_512_n269, _add_512_n268, _add_512_n267, _add_512_n266, _add_512_n265, _add_512_n264, _add_512_n263, _add_512_n262, _add_512_n261, _add_512_n260, _add_512_n259, _add_512_n258, _add_512_n257, _add_512_n256, _add_512_n255, _add_512_n254, _add_512_n253, _add_512_n252, _add_512_n251, _add_512_n250, _add_512_n249, _add_512_n248, _add_512_n247, _add_512_n246, _add_512_n245, _add_512_n244, _add_512_n243, _add_512_n242, _add_512_n241, _add_512_n240, _add_512_n239, _add_512_n238, _add_512_n237, _add_512_n236, _add_512_n235, _add_512_n234, _add_512_n233, _add_512_n232, _add_512_n231, _add_512_n230, _add_512_n229, 
  _add_512_n228, _add_512_n227, _add_512_n226, _add_512_n225, _add_512_n224, _add_512_n223, _add_512_n222, _add_512_n221, _add_512_n220, _add_512_n219, _add_512_n218, _add_512_n217, _add_512_n216, _add_512_n215, _add_512_n214, _add_512_n213, _add_512_n212, _add_512_n211, _add_512_n210, _add_512_n209, _add_512_n208, _add_512_n207, _add_512_n206, _add_512_n205, _add_512_n204, _add_512_n203, _add_512_n202, _add_512_n201, _add_512_n200, _add_512_n199, _add_512_n198, _add_512_n197, _add_512_n196, _add_512_n195, _add_512_n194, _add_512_n193, _add_512_n192, _add_512_n191, _add_512_n190, _add_512_n189, _add_512_n188, _add_512_n187, _add_512_n186, _add_512_n185, _add_512_n184, _add_512_n183, _add_512_n182, _add_512_n181, _add_512_n180, _add_512_n179, 
  _add_512_n178, _add_512_n177, _add_512_n176, _add_512_n175, _add_512_n174, _add_512_n173, _add_512_n172, _add_512_n171, _add_512_n170, _add_512_n169, _add_512_n168, _add_512_n167, _add_512_n166, _add_512_n165, _add_512_n164, _add_512_n163, _add_512_n162, _add_512_n161, _add_512_n160, _add_512_n159, _add_512_n158, _add_512_n157, _add_512_n156, _add_512_n155, _add_512_n154, _add_512_n153, _add_512_n152, _add_512_n151, _add_512_n150, _add_512_n149, _add_512_n148, _add_512_n147, _add_512_n146, _add_512_n145, _add_512_n144, _add_512_n143, _add_512_n142, _add_512_n141, _add_512_n140, _add_512_n139, _add_512_n138, _add_512_n137, _add_512_n136, _add_512_n135, _add_512_n134, _add_512_n133, _add_512_n132, _add_512_n131, _add_512_n130, _add_512_n129, 
  _add_512_n128, _add_512_n127, _add_512_n126, _add_512_n125, _add_512_n124, _add_512_n123, _add_512_n122, _add_512_n121, _add_512_n120, _add_512_n119, _add_512_n118, _add_512_n117, _add_512_n116, _add_512_n115, _add_512_n114, _add_512_n113, _add_512_n112, _add_512_n111, _add_512_n110, _add_512_n109, _add_512_n108, _add_512_n107, _add_512_n106, _add_512_n105, _add_512_n104, _add_512_n103, _add_512_n102, _add_512_n101, _add_512_n100, _add_512_n99, _add_512_n98, _add_512_n97, _add_512_n96, _add_512_n95, _add_512_n94, _add_512_n93, _add_512_n92, _add_512_n91, _add_512_n90, _add_512_n89, _add_512_n88, _add_512_n87, _add_512_n86, _add_512_n85, _add_512_n84, _add_512_n83, _add_512_n82, _add_512_n81, _add_512_n80, _add_512_n79, 
  _add_512_n78, _add_512_n77, _add_512_n76, _add_512_n75, _add_512_n74, _add_512_n73, _add_512_n72, _add_512_n71, _add_512_n70, _add_512_n69, _add_512_n68, _add_512_n67, _add_512_n66, _add_512_n65, _add_512_n64, _add_512_n63, _add_512_n62, _add_512_n61, _add_512_n60, _add_512_n59, _add_512_n58, _add_512_n57, _add_512_n56, _add_512_n55, _add_512_n54, _add_512_n53, _add_512_n52, _add_512_n51, _add_512_n50, _add_512_n49, _add_512_n48, _add_512_n47, _add_512_n46, _add_512_n45, _add_512_n44, _add_512_n43, _add_512_n42, _add_512_n41, _add_512_n40, _add_512_n39, _add_512_n38, _add_512_n37, _add_512_n36, _add_512_n35, _add_512_n34, _add_512_n33, _add_512_n32, _add_512_n31, _add_512_n30, _add_512_n29, 
  _add_512_n28, _add_512_n27, _add_512_n26, _add_512_n25, _add_512_n24, _add_512_n23, _add_512_n22, _add_512_n21, _add_512_n20, _add_512_n19, _add_512_n18, _add_512_n17, _add_512_n16, _add_512_n15, _add_512_n14, _add_512_n12, _add_512_n11, _add_512_n10, _add_512_n9, _add_512_n8, _add_512_n7, _add_512_n6, _add_512_n5, _add_512_n4, _add_512_n3, _add_512_n2, _add_512_n1, _add_0_root_add_136_4_n435, _add_0_root_add_136_4_n434, _add_0_root_add_136_4_n433, _add_0_root_add_136_4_n432, _add_0_root_add_136_4_n431, _add_0_root_add_136_4_n430, _add_0_root_add_136_4_n429, _add_0_root_add_136_4_n428, _add_0_root_add_136_4_n427, _add_0_root_add_136_4_n426, _add_0_root_add_136_4_n425, _add_0_root_add_136_4_n424, _add_0_root_add_136_4_n423, _add_0_root_add_136_4_n422, _add_0_root_add_136_4_n421, _add_0_root_add_136_4_n420, _add_0_root_add_136_4_n419, _add_0_root_add_136_4_n418, _add_0_root_add_136_4_n417, _add_0_root_add_136_4_n416, _add_0_root_add_136_4_n415, _add_0_root_add_136_4_n414, _add_0_root_add_136_4_n413, 
  _add_0_root_add_136_4_n412, _add_0_root_add_136_4_n411, _add_0_root_add_136_4_n410, _add_0_root_add_136_4_n409, _add_0_root_add_136_4_n408, _add_0_root_add_136_4_n407, _add_0_root_add_136_4_n406, _add_0_root_add_136_4_n405, _add_0_root_add_136_4_n404, _add_0_root_add_136_4_n403, _add_0_root_add_136_4_n402, _add_0_root_add_136_4_n401, _add_0_root_add_136_4_n400, _add_0_root_add_136_4_n399, _add_0_root_add_136_4_n398, _add_0_root_add_136_4_n397, _add_0_root_add_136_4_n396, _add_0_root_add_136_4_n395, _add_0_root_add_136_4_n394, _add_0_root_add_136_4_n393, _add_0_root_add_136_4_n392, _add_0_root_add_136_4_n391, _add_0_root_add_136_4_n390, _add_0_root_add_136_4_n389, _add_0_root_add_136_4_n388, _add_0_root_add_136_4_n387, _add_0_root_add_136_4_n386, _add_0_root_add_136_4_n385, _add_0_root_add_136_4_n384, _add_0_root_add_136_4_n383, _add_0_root_add_136_4_n382, _add_0_root_add_136_4_n381, _add_0_root_add_136_4_n380, _add_0_root_add_136_4_n379, _add_0_root_add_136_4_n378, _add_0_root_add_136_4_n377, _add_0_root_add_136_4_n376, _add_0_root_add_136_4_n375, _add_0_root_add_136_4_n374, _add_0_root_add_136_4_n373, _add_0_root_add_136_4_n372, _add_0_root_add_136_4_n371, _add_0_root_add_136_4_n370, _add_0_root_add_136_4_n369, _add_0_root_add_136_4_n368, _add_0_root_add_136_4_n367, _add_0_root_add_136_4_n366, _add_0_root_add_136_4_n365, _add_0_root_add_136_4_n364, _add_0_root_add_136_4_n363, 
  _add_0_root_add_136_4_n362, _add_0_root_add_136_4_n361, _add_0_root_add_136_4_n360, _add_0_root_add_136_4_n359, _add_0_root_add_136_4_n358, _add_0_root_add_136_4_n357, _add_0_root_add_136_4_n356, _add_0_root_add_136_4_n355, _add_0_root_add_136_4_n354, _add_0_root_add_136_4_n353, _add_0_root_add_136_4_n352, _add_0_root_add_136_4_n351, _add_0_root_add_136_4_n350, _add_0_root_add_136_4_n349, _add_0_root_add_136_4_n348, _add_0_root_add_136_4_n347, _add_0_root_add_136_4_n346, _add_0_root_add_136_4_n345, _add_0_root_add_136_4_n344, _add_0_root_add_136_4_n343, _add_0_root_add_136_4_n342, _add_0_root_add_136_4_n341, _add_0_root_add_136_4_n340, _add_0_root_add_136_4_n339, _add_0_root_add_136_4_n338, _add_0_root_add_136_4_n337, _add_0_root_add_136_4_n336, _add_0_root_add_136_4_n335, _add_0_root_add_136_4_n334, _add_0_root_add_136_4_n333, _add_0_root_add_136_4_n332, _add_0_root_add_136_4_n331, _add_0_root_add_136_4_n330, _add_0_root_add_136_4_n329, _add_0_root_add_136_4_n328, _add_0_root_add_136_4_n327, _add_0_root_add_136_4_n326, _add_0_root_add_136_4_n325, _add_0_root_add_136_4_n324, _add_0_root_add_136_4_n323, _add_0_root_add_136_4_n322, _add_0_root_add_136_4_n321, _add_0_root_add_136_4_n320, _add_0_root_add_136_4_n319, _add_0_root_add_136_4_n318, _add_0_root_add_136_4_n317, _add_0_root_add_136_4_n316, _add_0_root_add_136_4_n315, _add_0_root_add_136_4_n314, _add_0_root_add_136_4_n313, 
  _add_0_root_add_136_4_n312, _add_0_root_add_136_4_n311, _add_0_root_add_136_4_n310, _add_0_root_add_136_4_n309, _add_0_root_add_136_4_n308, _add_0_root_add_136_4_n307, _add_0_root_add_136_4_n306, _add_0_root_add_136_4_n305, _add_0_root_add_136_4_n304, _add_0_root_add_136_4_n303, _add_0_root_add_136_4_n302, _add_0_root_add_136_4_n301, _add_0_root_add_136_4_n300, _add_0_root_add_136_4_n299, _add_0_root_add_136_4_n298, _add_0_root_add_136_4_n297, _add_0_root_add_136_4_n296, _add_0_root_add_136_4_n295, _add_0_root_add_136_4_n294, _add_0_root_add_136_4_n293, _add_0_root_add_136_4_n292, _add_0_root_add_136_4_n291, _add_0_root_add_136_4_n290, _add_0_root_add_136_4_n289, _add_0_root_add_136_4_n288, _add_0_root_add_136_4_n287, _add_0_root_add_136_4_n286, _add_0_root_add_136_4_n285, _add_0_root_add_136_4_n284, _add_0_root_add_136_4_n283, _add_0_root_add_136_4_n282, _add_0_root_add_136_4_n281, _add_0_root_add_136_4_n280, _add_0_root_add_136_4_n279, _add_0_root_add_136_4_n278, _add_0_root_add_136_4_n277, _add_0_root_add_136_4_n276, _add_0_root_add_136_4_n275, _add_0_root_add_136_4_n274, _add_0_root_add_136_4_n273, _add_0_root_add_136_4_n272, _add_0_root_add_136_4_n271, _add_0_root_add_136_4_n270, _add_0_root_add_136_4_n269, _add_0_root_add_136_4_n268, _add_0_root_add_136_4_n267, _add_0_root_add_136_4_n266, _add_0_root_add_136_4_n265, _add_0_root_add_136_4_n264, _add_0_root_add_136_4_n263, 
  _add_0_root_add_136_4_n262, _add_0_root_add_136_4_n261, _add_0_root_add_136_4_n260, _add_0_root_add_136_4_n259, _add_0_root_add_136_4_n258, _add_0_root_add_136_4_n257, _add_0_root_add_136_4_n256, _add_0_root_add_136_4_n255, _add_0_root_add_136_4_n254, _add_0_root_add_136_4_n253, _add_0_root_add_136_4_n252, _add_0_root_add_136_4_n251, _add_0_root_add_136_4_n250, _add_0_root_add_136_4_n249, _add_0_root_add_136_4_n248, _add_0_root_add_136_4_n247, _add_0_root_add_136_4_n246, _add_0_root_add_136_4_n245, _add_0_root_add_136_4_n244, _add_0_root_add_136_4_n243, _add_0_root_add_136_4_n242, _add_0_root_add_136_4_n241, _add_0_root_add_136_4_n240, _add_0_root_add_136_4_n239, _add_0_root_add_136_4_n238, _add_0_root_add_136_4_n237, _add_0_root_add_136_4_n236, _add_0_root_add_136_4_n235, _add_0_root_add_136_4_n234, _add_0_root_add_136_4_n233, _add_0_root_add_136_4_n232, _add_0_root_add_136_4_n231, _add_0_root_add_136_4_n230, _add_0_root_add_136_4_n229, _add_0_root_add_136_4_n228, _add_0_root_add_136_4_n227, _add_0_root_add_136_4_n226, _add_0_root_add_136_4_n225, _add_0_root_add_136_4_n224, _add_0_root_add_136_4_n223, _add_0_root_add_136_4_n222, _add_0_root_add_136_4_n221, _add_0_root_add_136_4_n220, _add_0_root_add_136_4_n219, _add_0_root_add_136_4_n218, _add_0_root_add_136_4_n217, _add_0_root_add_136_4_n216, _add_0_root_add_136_4_n215, _add_0_root_add_136_4_n214, _add_0_root_add_136_4_n213, 
  _add_0_root_add_136_4_n212, _add_0_root_add_136_4_n211, _add_0_root_add_136_4_n210, _add_0_root_add_136_4_n209, _add_0_root_add_136_4_n208, _add_0_root_add_136_4_n207, _add_0_root_add_136_4_n206, _add_0_root_add_136_4_n205, _add_0_root_add_136_4_n204, _add_0_root_add_136_4_n203, _add_0_root_add_136_4_n202, _add_0_root_add_136_4_n201, _add_0_root_add_136_4_n200, _add_0_root_add_136_4_n199, _add_0_root_add_136_4_n198, _add_0_root_add_136_4_n197, _add_0_root_add_136_4_n196, _add_0_root_add_136_4_n195, _add_0_root_add_136_4_n194, _add_0_root_add_136_4_n193, _add_0_root_add_136_4_n192, _add_0_root_add_136_4_n191, _add_0_root_add_136_4_n190, _add_0_root_add_136_4_n189, _add_0_root_add_136_4_n188, _add_0_root_add_136_4_n187, _add_0_root_add_136_4_n186, _add_0_root_add_136_4_n185, _add_0_root_add_136_4_n184, _add_0_root_add_136_4_n183, _add_0_root_add_136_4_n182, _add_0_root_add_136_4_n181, _add_0_root_add_136_4_n180, _add_0_root_add_136_4_n179, _add_0_root_add_136_4_n178, _add_0_root_add_136_4_n177, _add_0_root_add_136_4_n176, _add_0_root_add_136_4_n175, _add_0_root_add_136_4_n174, _add_0_root_add_136_4_n173, _add_0_root_add_136_4_n172, _add_0_root_add_136_4_n171, _add_0_root_add_136_4_n170, _add_0_root_add_136_4_n169, _add_0_root_add_136_4_n168, _add_0_root_add_136_4_n167, _add_0_root_add_136_4_n166, _add_0_root_add_136_4_n165, _add_0_root_add_136_4_n164, _add_0_root_add_136_4_n163, 
  _add_0_root_add_136_4_n162, _add_0_root_add_136_4_n161, _add_0_root_add_136_4_n160, _add_0_root_add_136_4_n159, _add_0_root_add_136_4_n158, _add_0_root_add_136_4_n157, _add_0_root_add_136_4_n156, _add_0_root_add_136_4_n155, _add_0_root_add_136_4_n154, _add_0_root_add_136_4_n153, _add_0_root_add_136_4_n152, _add_0_root_add_136_4_n151, _add_0_root_add_136_4_n150, _add_0_root_add_136_4_n149, _add_0_root_add_136_4_n148, _add_0_root_add_136_4_n147, _add_0_root_add_136_4_n146, _add_0_root_add_136_4_n145, _add_0_root_add_136_4_n144, _add_0_root_add_136_4_n143, _add_0_root_add_136_4_n142, _add_0_root_add_136_4_n141, _add_0_root_add_136_4_n140, _add_0_root_add_136_4_n139, _add_0_root_add_136_4_n138, _add_0_root_add_136_4_n137, _add_0_root_add_136_4_n136, _add_0_root_add_136_4_n135, _add_0_root_add_136_4_n134, _add_0_root_add_136_4_n133, _add_0_root_add_136_4_n132, _add_0_root_add_136_4_n131, _add_0_root_add_136_4_n130, _add_0_root_add_136_4_n129, _add_0_root_add_136_4_n128, _add_0_root_add_136_4_n127, _add_0_root_add_136_4_n126, _add_0_root_add_136_4_n125, _add_0_root_add_136_4_n124, _add_0_root_add_136_4_n123, _add_0_root_add_136_4_n122, _add_0_root_add_136_4_n121, _add_0_root_add_136_4_n120, _add_0_root_add_136_4_n119, _add_0_root_add_136_4_n118, _add_0_root_add_136_4_n117, _add_0_root_add_136_4_n116, _add_0_root_add_136_4_n115, _add_0_root_add_136_4_n114, _add_0_root_add_136_4_n113, 
  _add_0_root_add_136_4_n112, _add_0_root_add_136_4_n111, _add_0_root_add_136_4_n110, _add_0_root_add_136_4_n109, _add_0_root_add_136_4_n108, _add_0_root_add_136_4_n107, _add_0_root_add_136_4_n106, _add_0_root_add_136_4_n105, _add_0_root_add_136_4_n104, _add_0_root_add_136_4_n103, _add_0_root_add_136_4_n102, _add_0_root_add_136_4_n101, _add_0_root_add_136_4_n100, _add_0_root_add_136_4_n99, _add_0_root_add_136_4_n98, _add_0_root_add_136_4_n97, _add_0_root_add_136_4_n96, _add_0_root_add_136_4_n95, _add_0_root_add_136_4_n94, _add_0_root_add_136_4_n93, _add_0_root_add_136_4_n92, _add_0_root_add_136_4_n91, _add_0_root_add_136_4_n90, _add_0_root_add_136_4_n89, _add_0_root_add_136_4_n88, _add_0_root_add_136_4_n87, _add_0_root_add_136_4_n86, _add_0_root_add_136_4_n85, _add_0_root_add_136_4_n84, _add_0_root_add_136_4_n83, _add_0_root_add_136_4_n82, _add_0_root_add_136_4_n81, _add_0_root_add_136_4_n77, _add_0_root_add_136_4_n75, _add_0_root_add_136_4_n73, _add_0_root_add_136_4_n72, _add_0_root_add_136_4_n71, _add_0_root_add_136_4_n70, _add_0_root_add_136_4_n66, _add_0_root_add_136_4_n65, _add_0_root_add_136_4_n64, _add_0_root_add_136_4_n63, _add_0_root_add_136_4_n62, _add_0_root_add_136_4_n61, _add_0_root_add_136_4_n60, _add_0_root_add_136_4_n59, _add_0_root_add_136_4_n58, _add_0_root_add_136_4_n57, _add_0_root_add_136_4_n56, _add_0_root_add_136_4_n55, 
  _add_0_root_add_136_4_n54, _add_0_root_add_136_4_n53, _add_0_root_add_136_4_n52, _add_0_root_add_136_4_n51, _add_0_root_add_136_4_n50, _add_0_root_add_136_4_n49, _add_0_root_add_136_4_n48, _add_0_root_add_136_4_n47, _add_0_root_add_136_4_n46, _add_0_root_add_136_4_n45, _add_0_root_add_136_4_n44, _add_0_root_add_136_4_n43, _add_0_root_add_136_4_n42, _add_0_root_add_136_4_n41, _add_0_root_add_136_4_n40, _add_0_root_add_136_4_n39, _add_0_root_add_136_4_n38, _add_0_root_add_136_4_n37, _add_0_root_add_136_4_n36, _add_0_root_add_136_4_n34, _add_0_root_add_136_4_n33, _add_0_root_add_136_4_n32, _add_0_root_add_136_4_n30, _add_0_root_add_136_4_n29, _add_0_root_add_136_4_n28, _add_0_root_add_136_4_n27, _add_0_root_add_136_4_n26, _add_0_root_add_136_4_n25, _add_0_root_add_136_4_n24, _add_0_root_add_136_4_n23, _add_0_root_add_136_4_n22, _add_0_root_add_136_4_n21, _add_0_root_add_136_4_n20, _add_0_root_add_136_4_n19, _add_0_root_add_136_4_n18, _add_0_root_add_136_4_n17, _add_0_root_add_136_4_n16, _add_0_root_add_136_4_n15, _add_0_root_add_136_4_n14, _add_0_root_add_136_4_n13, _add_0_root_add_136_4_n12, _add_0_root_add_136_4_n11, _add_0_root_add_136_4_n10, _add_0_root_add_136_4_n9, _add_0_root_add_136_4_n8, _add_0_root_add_136_4_n7, _add_0_root_add_136_4_n6, _add_0_root_add_136_4_n5, _add_0_root_add_136_4_n4, _add_0_root_add_136_4_n3, 
  _add_0_root_add_136_4_n2, _add_0_root_add_136_4_n1 ;
CLKBUFX1 gbuf_d_1(.A(n13067), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(cmd_o[1]));
CLKBUFX1 gbuf_qn_1(.A(qn_in_1), .Y(n345));
CLKBUFX1 gbuf_d_2(.A(n13128), .Y(d_out_2));
CLKBUFX1 gbuf_q_2(.A(q_in_2), .Y(round[0]));
CLKBUFX1 gbuf_qn_2(.A(qn_in_2), .Y(n13112));
CLKBUFX1 gbuf_d_3(.A(N1720), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(n13069));
CLKBUFX1 gbuf_qn_3(.A(qn_in_3), .Y(n13114));
CLKBUFX1 gbuf_d_4(.A(n13065), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(cmd_o[0]));
CLKBUFX1 gbuf_qn_4(.A(qn_in_4), .Y(n347));
CLKBUFX1 gbuf_d_5(.A(n4528), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(n14963));
CLKBUFX1 gbuf_d_6(.A(n4272), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(n14964));
CLKBUFX1 gbuf_d_7(.A(n4240), .Y(d_out_7));
CLKBUFX1 gbuf_q_7(.A(q_in_7), .Y(n14965));
CLKBUFX1 gbuf_d_8(.A(n4208), .Y(d_out_8));
CLKBUFX1 gbuf_q_8(.A(q_in_8), .Y(n14966));
CLKBUFX1 gbuf_d_9(.A(n4176), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(n14967));
CLKBUFX1 gbuf_d_10(.A(n4144), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(n14968));
CLKBUFX1 gbuf_d_11(.A(n4112), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(n14969));
CLKBUFX1 gbuf_qn_11(.A(qn_in_11), .Y(n12976));
CLKBUFX1 gbuf_d_12(.A(n4080), .Y(d_out_12));
CLKBUFX1 gbuf_q_12(.A(q_in_12), .Y(n14970));
CLKBUFX1 gbuf_d_13(.A(n4048), .Y(d_out_13));
CLKBUFX1 gbuf_q_13(.A(q_in_13), .Y(n14971));
CLKBUFX1 gbuf_d_14(.A(n4526), .Y(d_out_14));
CLKBUFX1 gbuf_q_14(.A(q_in_14), .Y(Wt[1]));
CLKBUFX1 gbuf_d_15(.A(n4494), .Y(d_out_15));
CLKBUFX1 gbuf_q_15(.A(q_in_15), .Y(n14934));
CLKBUFX1 gbuf_d_16(.A(n4462), .Y(d_out_16));
CLKBUFX1 gbuf_q_16(.A(q_in_16), .Y(n14972));
CLKBUFX1 gbuf_qn_16(.A(qn_in_16), .Y(n8320));
CLKBUFX1 gbuf_d_17(.A(n4430), .Y(d_out_17));
CLKBUFX1 gbuf_q_17(.A(q_in_17), .Y(n14973));
CLKBUFX1 gbuf_d_18(.A(n4398), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(n14974));
CLKBUFX1 gbuf_d_19(.A(n4366), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(n14975));
CLKBUFX1 gbuf_d_20(.A(n4334), .Y(d_out_20));
CLKBUFX1 gbuf_q_20(.A(q_in_20), .Y(n14976));
CLKBUFX1 gbuf_d_21(.A(n4303), .Y(d_out_21));
CLKBUFX1 gbuf_q_21(.A(q_in_21), .Y(n14977));
CLKBUFX1 gbuf_d_22(.A(n4271), .Y(d_out_22));
CLKBUFX1 gbuf_q_22(.A(q_in_22), .Y(n14978));
CLKBUFX1 gbuf_d_23(.A(n4239), .Y(d_out_23));
CLKBUFX1 gbuf_q_23(.A(q_in_23), .Y(n14979));
CLKBUFX1 gbuf_d_24(.A(n4207), .Y(d_out_24));
CLKBUFX1 gbuf_q_24(.A(q_in_24), .Y(n14980));
CLKBUFX1 gbuf_d_25(.A(n4175), .Y(d_out_25));
CLKBUFX1 gbuf_q_25(.A(q_in_25), .Y(n14981));
CLKBUFX1 gbuf_d_26(.A(n4143), .Y(d_out_26));
CLKBUFX1 gbuf_q_26(.A(q_in_26), .Y(n14982));
CLKBUFX1 gbuf_d_27(.A(n4111), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(n14983));
CLKBUFX1 gbuf_qn_27(.A(qn_in_27), .Y(n12974));
CLKBUFX1 gbuf_d_28(.A(n4079), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(n14984));
CLKBUFX1 gbuf_d_29(.A(n4047), .Y(d_out_29));
CLKBUFX1 gbuf_q_29(.A(q_in_29), .Y(n14985));
CLKBUFX1 gbuf_d_30(.A(n4525), .Y(d_out_30));
CLKBUFX1 gbuf_q_30(.A(q_in_30), .Y(Wt[2]));
CLKBUFX1 gbuf_d_31(.A(n4493), .Y(d_out_31));
CLKBUFX1 gbuf_q_31(.A(q_in_31), .Y(n14935));
CLKBUFX1 gbuf_d_32(.A(n4461), .Y(d_out_32));
CLKBUFX1 gbuf_q_32(.A(q_in_32), .Y(n14986));
CLKBUFX1 gbuf_qn_32(.A(qn_in_32), .Y(n8318));
CLKBUFX1 gbuf_d_33(.A(n4429), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(n14987));
CLKBUFX1 gbuf_d_34(.A(n4397), .Y(d_out_34));
CLKBUFX1 gbuf_q_34(.A(q_in_34), .Y(n14988));
CLKBUFX1 gbuf_d_35(.A(n4365), .Y(d_out_35));
CLKBUFX1 gbuf_q_35(.A(q_in_35), .Y(n14989));
CLKBUFX1 gbuf_d_36(.A(n4333), .Y(d_out_36));
CLKBUFX1 gbuf_q_36(.A(q_in_36), .Y(n14990));
CLKBUFX1 gbuf_d_37(.A(n4302), .Y(d_out_37));
CLKBUFX1 gbuf_q_37(.A(q_in_37), .Y(n14991));
CLKBUFX1 gbuf_d_38(.A(n4270), .Y(d_out_38));
CLKBUFX1 gbuf_q_38(.A(q_in_38), .Y(n14992));
CLKBUFX1 gbuf_d_39(.A(n4238), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(n14993));
CLKBUFX1 gbuf_d_40(.A(n4206), .Y(d_out_40));
CLKBUFX1 gbuf_q_40(.A(q_in_40), .Y(n14994));
CLKBUFX1 gbuf_d_41(.A(n4174), .Y(d_out_41));
CLKBUFX1 gbuf_q_41(.A(q_in_41), .Y(n14995));
CLKBUFX1 gbuf_d_42(.A(n4142), .Y(d_out_42));
CLKBUFX1 gbuf_q_42(.A(q_in_42), .Y(n14996));
CLKBUFX1 gbuf_d_43(.A(n4110), .Y(d_out_43));
CLKBUFX1 gbuf_q_43(.A(q_in_43), .Y(n14997));
CLKBUFX1 gbuf_qn_43(.A(qn_in_43), .Y(n12972));
CLKBUFX1 gbuf_d_44(.A(n4078), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(n14998));
CLKBUFX1 gbuf_d_45(.A(n4046), .Y(d_out_45));
CLKBUFX1 gbuf_q_45(.A(q_in_45), .Y(n14999));
CLKBUFX1 gbuf_d_46(.A(n4524), .Y(d_out_46));
CLKBUFX1 gbuf_q_46(.A(q_in_46), .Y(Wt[3]));
CLKBUFX1 gbuf_d_47(.A(n4492), .Y(d_out_47));
CLKBUFX1 gbuf_q_47(.A(q_in_47), .Y(n14936));
CLKBUFX1 gbuf_d_48(.A(n4460), .Y(d_out_48));
CLKBUFX1 gbuf_q_48(.A(q_in_48), .Y(n15000));
CLKBUFX1 gbuf_qn_48(.A(qn_in_48), .Y(n8316));
CLKBUFX1 gbuf_d_49(.A(n4428), .Y(d_out_49));
CLKBUFX1 gbuf_q_49(.A(q_in_49), .Y(n15001));
CLKBUFX1 gbuf_d_50(.A(n4396), .Y(d_out_50));
CLKBUFX1 gbuf_q_50(.A(q_in_50), .Y(n15002));
CLKBUFX1 gbuf_d_51(.A(n4364), .Y(d_out_51));
CLKBUFX1 gbuf_q_51(.A(q_in_51), .Y(n15003));
CLKBUFX1 gbuf_d_52(.A(n4332), .Y(d_out_52));
CLKBUFX1 gbuf_q_52(.A(q_in_52), .Y(n15004));
CLKBUFX1 gbuf_d_53(.A(n4301), .Y(d_out_53));
CLKBUFX1 gbuf_q_53(.A(q_in_53), .Y(n15005));
CLKBUFX1 gbuf_d_54(.A(n4269), .Y(d_out_54));
CLKBUFX1 gbuf_q_54(.A(q_in_54), .Y(n15006));
CLKBUFX1 gbuf_d_55(.A(n4237), .Y(d_out_55));
CLKBUFX1 gbuf_q_55(.A(q_in_55), .Y(n15007));
CLKBUFX1 gbuf_d_56(.A(n4205), .Y(d_out_56));
CLKBUFX1 gbuf_q_56(.A(q_in_56), .Y(n15008));
CLKBUFX1 gbuf_d_57(.A(n4173), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(n15009));
CLKBUFX1 gbuf_d_58(.A(n4141), .Y(d_out_58));
CLKBUFX1 gbuf_q_58(.A(q_in_58), .Y(n15010));
CLKBUFX1 gbuf_d_59(.A(n4109), .Y(d_out_59));
CLKBUFX1 gbuf_q_59(.A(q_in_59), .Y(n15011));
CLKBUFX1 gbuf_qn_59(.A(qn_in_59), .Y(n12970));
CLKBUFX1 gbuf_d_60(.A(n4077), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(n15012));
CLKBUFX1 gbuf_d_61(.A(n4045), .Y(d_out_61));
CLKBUFX1 gbuf_q_61(.A(q_in_61), .Y(n15013));
CLKBUFX1 gbuf_d_62(.A(n4523), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(Wt[4]));
CLKBUFX1 gbuf_d_63(.A(n4491), .Y(d_out_63));
CLKBUFX1 gbuf_q_63(.A(q_in_63), .Y(n14937));
CLKBUFX1 gbuf_d_64(.A(n4459), .Y(d_out_64));
CLKBUFX1 gbuf_q_64(.A(q_in_64), .Y(n15014));
CLKBUFX1 gbuf_qn_64(.A(qn_in_64), .Y(n8314));
CLKBUFX1 gbuf_d_65(.A(n4427), .Y(d_out_65));
CLKBUFX1 gbuf_q_65(.A(q_in_65), .Y(n15015));
CLKBUFX1 gbuf_d_66(.A(n4395), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(n15016));
CLKBUFX1 gbuf_d_67(.A(n4363), .Y(d_out_67));
CLKBUFX1 gbuf_q_67(.A(q_in_67), .Y(n15017));
CLKBUFX1 gbuf_d_68(.A(n4331), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(n15018));
CLKBUFX1 gbuf_d_69(.A(n4300), .Y(d_out_69));
CLKBUFX1 gbuf_q_69(.A(q_in_69), .Y(n15019));
CLKBUFX1 gbuf_d_70(.A(n4268), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(n15020));
CLKBUFX1 gbuf_d_71(.A(n4236), .Y(d_out_71));
CLKBUFX1 gbuf_q_71(.A(q_in_71), .Y(n15021));
CLKBUFX1 gbuf_d_72(.A(n4204), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(n15022));
CLKBUFX1 gbuf_d_73(.A(n4172), .Y(d_out_73));
CLKBUFX1 gbuf_q_73(.A(q_in_73), .Y(n15023));
CLKBUFX1 gbuf_d_74(.A(n4140), .Y(d_out_74));
CLKBUFX1 gbuf_q_74(.A(q_in_74), .Y(n15024));
CLKBUFX1 gbuf_d_75(.A(n4108), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(n15025));
CLKBUFX1 gbuf_qn_75(.A(qn_in_75), .Y(n12968));
CLKBUFX1 gbuf_d_76(.A(n4076), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(n15026));
CLKBUFX1 gbuf_d_77(.A(n4044), .Y(d_out_77));
CLKBUFX1 gbuf_q_77(.A(q_in_77), .Y(n15027));
CLKBUFX1 gbuf_d_78(.A(n4522), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(Wt[5]));
CLKBUFX1 gbuf_d_79(.A(n4490), .Y(d_out_79));
CLKBUFX1 gbuf_q_79(.A(q_in_79), .Y(n14938));
CLKBUFX1 gbuf_d_80(.A(n4458), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(n15028));
CLKBUFX1 gbuf_qn_80(.A(qn_in_80), .Y(n8312));
CLKBUFX1 gbuf_d_81(.A(n4426), .Y(d_out_81));
CLKBUFX1 gbuf_q_81(.A(q_in_81), .Y(n15029));
CLKBUFX1 gbuf_d_82(.A(n4394), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(n15030));
CLKBUFX1 gbuf_d_83(.A(n4362), .Y(d_out_83));
CLKBUFX1 gbuf_q_83(.A(q_in_83), .Y(n15031));
CLKBUFX1 gbuf_d_84(.A(n4330), .Y(d_out_84));
CLKBUFX1 gbuf_q_84(.A(q_in_84), .Y(n15032));
CLKBUFX1 gbuf_d_85(.A(n4299), .Y(d_out_85));
CLKBUFX1 gbuf_q_85(.A(q_in_85), .Y(n15033));
CLKBUFX1 gbuf_d_86(.A(n4267), .Y(d_out_86));
CLKBUFX1 gbuf_q_86(.A(q_in_86), .Y(n15034));
CLKBUFX1 gbuf_d_87(.A(n4235), .Y(d_out_87));
CLKBUFX1 gbuf_q_87(.A(q_in_87), .Y(n15035));
CLKBUFX1 gbuf_d_88(.A(n4203), .Y(d_out_88));
CLKBUFX1 gbuf_q_88(.A(q_in_88), .Y(n15036));
CLKBUFX1 gbuf_d_89(.A(n4171), .Y(d_out_89));
CLKBUFX1 gbuf_q_89(.A(q_in_89), .Y(n15037));
CLKBUFX1 gbuf_d_90(.A(n4139), .Y(d_out_90));
CLKBUFX1 gbuf_q_90(.A(q_in_90), .Y(n15038));
CLKBUFX1 gbuf_d_91(.A(n4107), .Y(d_out_91));
CLKBUFX1 gbuf_q_91(.A(q_in_91), .Y(n15039));
CLKBUFX1 gbuf_qn_91(.A(qn_in_91), .Y(n12966));
CLKBUFX1 gbuf_d_92(.A(n4075), .Y(d_out_92));
CLKBUFX1 gbuf_q_92(.A(q_in_92), .Y(n15040));
CLKBUFX1 gbuf_d_93(.A(n4043), .Y(d_out_93));
CLKBUFX1 gbuf_q_93(.A(q_in_93), .Y(n15041));
CLKBUFX1 gbuf_d_94(.A(n4521), .Y(d_out_94));
CLKBUFX1 gbuf_q_94(.A(q_in_94), .Y(Wt[6]));
CLKBUFX1 gbuf_d_95(.A(n4489), .Y(d_out_95));
CLKBUFX1 gbuf_q_95(.A(q_in_95), .Y(n14939));
CLKBUFX1 gbuf_d_96(.A(n4457), .Y(d_out_96));
CLKBUFX1 gbuf_q_96(.A(q_in_96), .Y(n15042));
CLKBUFX1 gbuf_qn_96(.A(qn_in_96), .Y(n8310));
CLKBUFX1 gbuf_d_97(.A(n4425), .Y(d_out_97));
CLKBUFX1 gbuf_q_97(.A(q_in_97), .Y(n15043));
CLKBUFX1 gbuf_d_98(.A(n4393), .Y(d_out_98));
CLKBUFX1 gbuf_q_98(.A(q_in_98), .Y(n15044));
CLKBUFX1 gbuf_d_99(.A(n4361), .Y(d_out_99));
CLKBUFX1 gbuf_q_99(.A(q_in_99), .Y(n15045));
CLKBUFX1 gbuf_d_100(.A(n4329), .Y(d_out_100));
CLKBUFX1 gbuf_q_100(.A(q_in_100), .Y(n15046));
CLKBUFX1 gbuf_d_101(.A(n4298), .Y(d_out_101));
CLKBUFX1 gbuf_q_101(.A(q_in_101), .Y(n15047));
CLKBUFX1 gbuf_d_102(.A(n4266), .Y(d_out_102));
CLKBUFX1 gbuf_q_102(.A(q_in_102), .Y(n15048));
CLKBUFX1 gbuf_d_103(.A(n4234), .Y(d_out_103));
CLKBUFX1 gbuf_q_103(.A(q_in_103), .Y(n15049));
CLKBUFX1 gbuf_d_104(.A(n4202), .Y(d_out_104));
CLKBUFX1 gbuf_q_104(.A(q_in_104), .Y(n15050));
CLKBUFX1 gbuf_d_105(.A(n4170), .Y(d_out_105));
CLKBUFX1 gbuf_q_105(.A(q_in_105), .Y(n15051));
CLKBUFX1 gbuf_d_106(.A(n4138), .Y(d_out_106));
CLKBUFX1 gbuf_q_106(.A(q_in_106), .Y(n15052));
CLKBUFX1 gbuf_d_107(.A(n4106), .Y(d_out_107));
CLKBUFX1 gbuf_q_107(.A(q_in_107), .Y(n15053));
CLKBUFX1 gbuf_qn_107(.A(qn_in_107), .Y(n12964));
CLKBUFX1 gbuf_d_108(.A(n4074), .Y(d_out_108));
CLKBUFX1 gbuf_q_108(.A(q_in_108), .Y(n15054));
CLKBUFX1 gbuf_d_109(.A(n4042), .Y(d_out_109));
CLKBUFX1 gbuf_q_109(.A(q_in_109), .Y(n15055));
CLKBUFX1 gbuf_d_110(.A(n4520), .Y(d_out_110));
CLKBUFX1 gbuf_q_110(.A(q_in_110), .Y(Wt[7]));
CLKBUFX1 gbuf_d_111(.A(n4488), .Y(d_out_111));
CLKBUFX1 gbuf_q_111(.A(q_in_111), .Y(n14940));
CLKBUFX1 gbuf_d_112(.A(n4456), .Y(d_out_112));
CLKBUFX1 gbuf_q_112(.A(q_in_112), .Y(n15056));
CLKBUFX1 gbuf_qn_112(.A(qn_in_112), .Y(n8308));
CLKBUFX1 gbuf_d_113(.A(n4424), .Y(d_out_113));
CLKBUFX1 gbuf_q_113(.A(q_in_113), .Y(n15057));
CLKBUFX1 gbuf_d_114(.A(n4392), .Y(d_out_114));
CLKBUFX1 gbuf_q_114(.A(q_in_114), .Y(n15058));
CLKBUFX1 gbuf_d_115(.A(n4360), .Y(d_out_115));
CLKBUFX1 gbuf_q_115(.A(q_in_115), .Y(n15059));
CLKBUFX1 gbuf_d_116(.A(n4328), .Y(d_out_116));
CLKBUFX1 gbuf_q_116(.A(q_in_116), .Y(n15060));
CLKBUFX1 gbuf_d_117(.A(n4297), .Y(d_out_117));
CLKBUFX1 gbuf_q_117(.A(q_in_117), .Y(n15061));
CLKBUFX1 gbuf_d_118(.A(n4265), .Y(d_out_118));
CLKBUFX1 gbuf_q_118(.A(q_in_118), .Y(n15062));
CLKBUFX1 gbuf_d_119(.A(n4233), .Y(d_out_119));
CLKBUFX1 gbuf_q_119(.A(q_in_119), .Y(n15063));
CLKBUFX1 gbuf_d_120(.A(n4201), .Y(d_out_120));
CLKBUFX1 gbuf_q_120(.A(q_in_120), .Y(n15064));
CLKBUFX1 gbuf_d_121(.A(n4169), .Y(d_out_121));
CLKBUFX1 gbuf_q_121(.A(q_in_121), .Y(n15065));
CLKBUFX1 gbuf_d_122(.A(n4137), .Y(d_out_122));
CLKBUFX1 gbuf_q_122(.A(q_in_122), .Y(n15066));
CLKBUFX1 gbuf_d_123(.A(n4105), .Y(d_out_123));
CLKBUFX1 gbuf_q_123(.A(q_in_123), .Y(n15067));
CLKBUFX1 gbuf_qn_123(.A(qn_in_123), .Y(n12962));
CLKBUFX1 gbuf_d_124(.A(n4073), .Y(d_out_124));
CLKBUFX1 gbuf_q_124(.A(q_in_124), .Y(n15068));
CLKBUFX1 gbuf_d_125(.A(n4041), .Y(d_out_125));
CLKBUFX1 gbuf_q_125(.A(q_in_125), .Y(n15069));
CLKBUFX1 gbuf_d_126(.A(n4519), .Y(d_out_126));
CLKBUFX1 gbuf_q_126(.A(q_in_126), .Y(Wt[8]));
CLKBUFX1 gbuf_d_127(.A(n4487), .Y(d_out_127));
CLKBUFX1 gbuf_q_127(.A(q_in_127), .Y(n14941));
CLKBUFX1 gbuf_d_128(.A(n4455), .Y(d_out_128));
CLKBUFX1 gbuf_q_128(.A(q_in_128), .Y(n15070));
CLKBUFX1 gbuf_qn_128(.A(qn_in_128), .Y(n8306));
CLKBUFX1 gbuf_d_129(.A(n4423), .Y(d_out_129));
CLKBUFX1 gbuf_q_129(.A(q_in_129), .Y(n15071));
CLKBUFX1 gbuf_d_130(.A(n4391), .Y(d_out_130));
CLKBUFX1 gbuf_q_130(.A(q_in_130), .Y(n15072));
CLKBUFX1 gbuf_d_131(.A(n4359), .Y(d_out_131));
CLKBUFX1 gbuf_q_131(.A(q_in_131), .Y(n15073));
CLKBUFX1 gbuf_d_132(.A(n4327), .Y(d_out_132));
CLKBUFX1 gbuf_q_132(.A(q_in_132), .Y(n15074));
CLKBUFX1 gbuf_d_133(.A(n4296), .Y(d_out_133));
CLKBUFX1 gbuf_q_133(.A(q_in_133), .Y(n15075));
CLKBUFX1 gbuf_d_134(.A(n4264), .Y(d_out_134));
CLKBUFX1 gbuf_q_134(.A(q_in_134), .Y(n15076));
CLKBUFX1 gbuf_d_135(.A(n4232), .Y(d_out_135));
CLKBUFX1 gbuf_q_135(.A(q_in_135), .Y(n15077));
CLKBUFX1 gbuf_d_136(.A(n4200), .Y(d_out_136));
CLKBUFX1 gbuf_q_136(.A(q_in_136), .Y(n15078));
CLKBUFX1 gbuf_d_137(.A(n4168), .Y(d_out_137));
CLKBUFX1 gbuf_q_137(.A(q_in_137), .Y(n15079));
CLKBUFX1 gbuf_d_138(.A(n4136), .Y(d_out_138));
CLKBUFX1 gbuf_q_138(.A(q_in_138), .Y(n15080));
CLKBUFX1 gbuf_d_139(.A(n4104), .Y(d_out_139));
CLKBUFX1 gbuf_q_139(.A(q_in_139), .Y(n15081));
CLKBUFX1 gbuf_qn_139(.A(qn_in_139), .Y(n12960));
CLKBUFX1 gbuf_d_140(.A(n4072), .Y(d_out_140));
CLKBUFX1 gbuf_q_140(.A(q_in_140), .Y(n15082));
CLKBUFX1 gbuf_d_141(.A(n4040), .Y(d_out_141));
CLKBUFX1 gbuf_q_141(.A(q_in_141), .Y(n15083));
CLKBUFX1 gbuf_d_142(.A(n4518), .Y(d_out_142));
CLKBUFX1 gbuf_q_142(.A(q_in_142), .Y(Wt[9]));
CLKBUFX1 gbuf_d_143(.A(n4486), .Y(d_out_143));
CLKBUFX1 gbuf_q_143(.A(q_in_143), .Y(n14942));
CLKBUFX1 gbuf_d_144(.A(n4454), .Y(d_out_144));
CLKBUFX1 gbuf_q_144(.A(q_in_144), .Y(n15084));
CLKBUFX1 gbuf_qn_144(.A(qn_in_144), .Y(n8304));
CLKBUFX1 gbuf_d_145(.A(n4422), .Y(d_out_145));
CLKBUFX1 gbuf_q_145(.A(q_in_145), .Y(n15085));
CLKBUFX1 gbuf_d_146(.A(n4390), .Y(d_out_146));
CLKBUFX1 gbuf_q_146(.A(q_in_146), .Y(n15086));
CLKBUFX1 gbuf_d_147(.A(n4358), .Y(d_out_147));
CLKBUFX1 gbuf_q_147(.A(q_in_147), .Y(n15087));
CLKBUFX1 gbuf_d_148(.A(n4326), .Y(d_out_148));
CLKBUFX1 gbuf_q_148(.A(q_in_148), .Y(n15088));
CLKBUFX1 gbuf_d_149(.A(n4295), .Y(d_out_149));
CLKBUFX1 gbuf_q_149(.A(q_in_149), .Y(n15089));
CLKBUFX1 gbuf_d_150(.A(n4263), .Y(d_out_150));
CLKBUFX1 gbuf_q_150(.A(q_in_150), .Y(n15090));
CLKBUFX1 gbuf_d_151(.A(n4231), .Y(d_out_151));
CLKBUFX1 gbuf_q_151(.A(q_in_151), .Y(n15091));
CLKBUFX1 gbuf_d_152(.A(n4199), .Y(d_out_152));
CLKBUFX1 gbuf_q_152(.A(q_in_152), .Y(n15092));
CLKBUFX1 gbuf_d_153(.A(n4167), .Y(d_out_153));
CLKBUFX1 gbuf_q_153(.A(q_in_153), .Y(n15093));
CLKBUFX1 gbuf_d_154(.A(n4135), .Y(d_out_154));
CLKBUFX1 gbuf_q_154(.A(q_in_154), .Y(n15094));
CLKBUFX1 gbuf_d_155(.A(n4103), .Y(d_out_155));
CLKBUFX1 gbuf_q_155(.A(q_in_155), .Y(n15095));
CLKBUFX1 gbuf_qn_155(.A(qn_in_155), .Y(n12958));
CLKBUFX1 gbuf_d_156(.A(n4071), .Y(d_out_156));
CLKBUFX1 gbuf_q_156(.A(q_in_156), .Y(n15096));
CLKBUFX1 gbuf_d_157(.A(n4039), .Y(d_out_157));
CLKBUFX1 gbuf_q_157(.A(q_in_157), .Y(n15097));
CLKBUFX1 gbuf_d_158(.A(n4517), .Y(d_out_158));
CLKBUFX1 gbuf_q_158(.A(q_in_158), .Y(Wt[10]));
CLKBUFX1 gbuf_d_159(.A(n4485), .Y(d_out_159));
CLKBUFX1 gbuf_q_159(.A(q_in_159), .Y(n14943));
CLKBUFX1 gbuf_d_160(.A(n4453), .Y(d_out_160));
CLKBUFX1 gbuf_q_160(.A(q_in_160), .Y(n15098));
CLKBUFX1 gbuf_qn_160(.A(qn_in_160), .Y(n8302));
CLKBUFX1 gbuf_d_161(.A(n4421), .Y(d_out_161));
CLKBUFX1 gbuf_q_161(.A(q_in_161), .Y(n15099));
CLKBUFX1 gbuf_d_162(.A(n4389), .Y(d_out_162));
CLKBUFX1 gbuf_q_162(.A(q_in_162), .Y(n15100));
CLKBUFX1 gbuf_d_163(.A(n4357), .Y(d_out_163));
CLKBUFX1 gbuf_q_163(.A(q_in_163), .Y(n15101));
CLKBUFX1 gbuf_d_164(.A(n4325), .Y(d_out_164));
CLKBUFX1 gbuf_q_164(.A(q_in_164), .Y(n15102));
CLKBUFX1 gbuf_d_165(.A(n4294), .Y(d_out_165));
CLKBUFX1 gbuf_q_165(.A(q_in_165), .Y(n15103));
CLKBUFX1 gbuf_d_166(.A(n4262), .Y(d_out_166));
CLKBUFX1 gbuf_q_166(.A(q_in_166), .Y(n15104));
CLKBUFX1 gbuf_d_167(.A(n4230), .Y(d_out_167));
CLKBUFX1 gbuf_q_167(.A(q_in_167), .Y(n15105));
CLKBUFX1 gbuf_d_168(.A(n4198), .Y(d_out_168));
CLKBUFX1 gbuf_q_168(.A(q_in_168), .Y(n15106));
CLKBUFX1 gbuf_d_169(.A(n4166), .Y(d_out_169));
CLKBUFX1 gbuf_q_169(.A(q_in_169), .Y(n15107));
CLKBUFX1 gbuf_d_170(.A(n4134), .Y(d_out_170));
CLKBUFX1 gbuf_q_170(.A(q_in_170), .Y(n15108));
CLKBUFX1 gbuf_d_171(.A(n4102), .Y(d_out_171));
CLKBUFX1 gbuf_q_171(.A(q_in_171), .Y(n15109));
CLKBUFX1 gbuf_qn_171(.A(qn_in_171), .Y(n12956));
CLKBUFX1 gbuf_d_172(.A(n4070), .Y(d_out_172));
CLKBUFX1 gbuf_q_172(.A(q_in_172), .Y(n15110));
CLKBUFX1 gbuf_d_173(.A(n4038), .Y(d_out_173));
CLKBUFX1 gbuf_q_173(.A(q_in_173), .Y(n15111));
CLKBUFX1 gbuf_d_174(.A(n4516), .Y(d_out_174));
CLKBUFX1 gbuf_q_174(.A(q_in_174), .Y(Wt[11]));
CLKBUFX1 gbuf_d_175(.A(n4484), .Y(d_out_175));
CLKBUFX1 gbuf_q_175(.A(q_in_175), .Y(n14944));
CLKBUFX1 gbuf_d_176(.A(n4452), .Y(d_out_176));
CLKBUFX1 gbuf_q_176(.A(q_in_176), .Y(n15112));
CLKBUFX1 gbuf_qn_176(.A(qn_in_176), .Y(n8300));
CLKBUFX1 gbuf_d_177(.A(n4420), .Y(d_out_177));
CLKBUFX1 gbuf_q_177(.A(q_in_177), .Y(n15113));
CLKBUFX1 gbuf_d_178(.A(n4388), .Y(d_out_178));
CLKBUFX1 gbuf_q_178(.A(q_in_178), .Y(n15114));
CLKBUFX1 gbuf_d_179(.A(n4356), .Y(d_out_179));
CLKBUFX1 gbuf_q_179(.A(q_in_179), .Y(n15115));
CLKBUFX1 gbuf_d_180(.A(n4324), .Y(d_out_180));
CLKBUFX1 gbuf_q_180(.A(q_in_180), .Y(n15116));
CLKBUFX1 gbuf_d_181(.A(n4293), .Y(d_out_181));
CLKBUFX1 gbuf_q_181(.A(q_in_181), .Y(n15117));
CLKBUFX1 gbuf_d_182(.A(n4261), .Y(d_out_182));
CLKBUFX1 gbuf_q_182(.A(q_in_182), .Y(n15118));
CLKBUFX1 gbuf_d_183(.A(n4229), .Y(d_out_183));
CLKBUFX1 gbuf_q_183(.A(q_in_183), .Y(n15119));
CLKBUFX1 gbuf_d_184(.A(n4197), .Y(d_out_184));
CLKBUFX1 gbuf_q_184(.A(q_in_184), .Y(n15120));
CLKBUFX1 gbuf_d_185(.A(n4165), .Y(d_out_185));
CLKBUFX1 gbuf_q_185(.A(q_in_185), .Y(n15121));
CLKBUFX1 gbuf_d_186(.A(n4133), .Y(d_out_186));
CLKBUFX1 gbuf_q_186(.A(q_in_186), .Y(n15122));
CLKBUFX1 gbuf_d_187(.A(n4101), .Y(d_out_187));
CLKBUFX1 gbuf_q_187(.A(q_in_187), .Y(n15123));
CLKBUFX1 gbuf_qn_187(.A(qn_in_187), .Y(n12954));
CLKBUFX1 gbuf_d_188(.A(n4069), .Y(d_out_188));
CLKBUFX1 gbuf_q_188(.A(q_in_188), .Y(n15124));
CLKBUFX1 gbuf_d_189(.A(n4037), .Y(d_out_189));
CLKBUFX1 gbuf_q_189(.A(q_in_189), .Y(n15125));
CLKBUFX1 gbuf_d_190(.A(n4515), .Y(d_out_190));
CLKBUFX1 gbuf_q_190(.A(q_in_190), .Y(Wt[12]));
CLKBUFX1 gbuf_d_191(.A(n4483), .Y(d_out_191));
CLKBUFX1 gbuf_q_191(.A(q_in_191), .Y(n14945));
CLKBUFX1 gbuf_d_192(.A(n4451), .Y(d_out_192));
CLKBUFX1 gbuf_q_192(.A(q_in_192), .Y(n15126));
CLKBUFX1 gbuf_qn_192(.A(qn_in_192), .Y(n8298));
CLKBUFX1 gbuf_d_193(.A(n4419), .Y(d_out_193));
CLKBUFX1 gbuf_q_193(.A(q_in_193), .Y(n15127));
CLKBUFX1 gbuf_d_194(.A(n4387), .Y(d_out_194));
CLKBUFX1 gbuf_q_194(.A(q_in_194), .Y(n15128));
CLKBUFX1 gbuf_d_195(.A(n4355), .Y(d_out_195));
CLKBUFX1 gbuf_q_195(.A(q_in_195), .Y(n15129));
CLKBUFX1 gbuf_d_196(.A(n4323), .Y(d_out_196));
CLKBUFX1 gbuf_q_196(.A(q_in_196), .Y(n15130));
CLKBUFX1 gbuf_d_197(.A(n4292), .Y(d_out_197));
CLKBUFX1 gbuf_q_197(.A(q_in_197), .Y(n15131));
CLKBUFX1 gbuf_d_198(.A(n4260), .Y(d_out_198));
CLKBUFX1 gbuf_q_198(.A(q_in_198), .Y(n15132));
CLKBUFX1 gbuf_d_199(.A(n4228), .Y(d_out_199));
CLKBUFX1 gbuf_q_199(.A(q_in_199), .Y(n15133));
CLKBUFX1 gbuf_d_200(.A(n4196), .Y(d_out_200));
CLKBUFX1 gbuf_q_200(.A(q_in_200), .Y(n15134));
CLKBUFX1 gbuf_d_201(.A(n4164), .Y(d_out_201));
CLKBUFX1 gbuf_q_201(.A(q_in_201), .Y(n15135));
CLKBUFX1 gbuf_d_202(.A(n4132), .Y(d_out_202));
CLKBUFX1 gbuf_q_202(.A(q_in_202), .Y(n15136));
CLKBUFX1 gbuf_d_203(.A(n4100), .Y(d_out_203));
CLKBUFX1 gbuf_q_203(.A(q_in_203), .Y(n15137));
CLKBUFX1 gbuf_qn_203(.A(qn_in_203), .Y(n12952));
CLKBUFX1 gbuf_d_204(.A(n4068), .Y(d_out_204));
CLKBUFX1 gbuf_q_204(.A(q_in_204), .Y(n15138));
CLKBUFX1 gbuf_d_205(.A(n4036), .Y(d_out_205));
CLKBUFX1 gbuf_q_205(.A(q_in_205), .Y(n15139));
CLKBUFX1 gbuf_d_206(.A(n4514), .Y(d_out_206));
CLKBUFX1 gbuf_q_206(.A(q_in_206), .Y(Wt[13]));
CLKBUFX1 gbuf_d_207(.A(n4482), .Y(d_out_207));
CLKBUFX1 gbuf_q_207(.A(q_in_207), .Y(n14946));
CLKBUFX1 gbuf_d_208(.A(n4450), .Y(d_out_208));
CLKBUFX1 gbuf_q_208(.A(q_in_208), .Y(n15140));
CLKBUFX1 gbuf_qn_208(.A(qn_in_208), .Y(n8296));
CLKBUFX1 gbuf_d_209(.A(n4418), .Y(d_out_209));
CLKBUFX1 gbuf_q_209(.A(q_in_209), .Y(n15141));
CLKBUFX1 gbuf_d_210(.A(n4386), .Y(d_out_210));
CLKBUFX1 gbuf_q_210(.A(q_in_210), .Y(n15142));
CLKBUFX1 gbuf_d_211(.A(n4354), .Y(d_out_211));
CLKBUFX1 gbuf_q_211(.A(q_in_211), .Y(n15143));
CLKBUFX1 gbuf_d_212(.A(n4322), .Y(d_out_212));
CLKBUFX1 gbuf_q_212(.A(q_in_212), .Y(n15144));
CLKBUFX1 gbuf_d_213(.A(n4291), .Y(d_out_213));
CLKBUFX1 gbuf_q_213(.A(q_in_213), .Y(n15145));
CLKBUFX1 gbuf_d_214(.A(n4259), .Y(d_out_214));
CLKBUFX1 gbuf_q_214(.A(q_in_214), .Y(n15146));
CLKBUFX1 gbuf_d_215(.A(n4227), .Y(d_out_215));
CLKBUFX1 gbuf_q_215(.A(q_in_215), .Y(n15147));
CLKBUFX1 gbuf_d_216(.A(n4195), .Y(d_out_216));
CLKBUFX1 gbuf_q_216(.A(q_in_216), .Y(n15148));
CLKBUFX1 gbuf_d_217(.A(n4163), .Y(d_out_217));
CLKBUFX1 gbuf_q_217(.A(q_in_217), .Y(n15149));
CLKBUFX1 gbuf_d_218(.A(n4131), .Y(d_out_218));
CLKBUFX1 gbuf_q_218(.A(q_in_218), .Y(n15150));
CLKBUFX1 gbuf_d_219(.A(n4099), .Y(d_out_219));
CLKBUFX1 gbuf_q_219(.A(q_in_219), .Y(n15151));
CLKBUFX1 gbuf_qn_219(.A(qn_in_219), .Y(n12950));
CLKBUFX1 gbuf_d_220(.A(n4067), .Y(d_out_220));
CLKBUFX1 gbuf_q_220(.A(q_in_220), .Y(n15152));
CLKBUFX1 gbuf_d_221(.A(n4035), .Y(d_out_221));
CLKBUFX1 gbuf_q_221(.A(q_in_221), .Y(n15153));
CLKBUFX1 gbuf_d_222(.A(n4513), .Y(d_out_222));
CLKBUFX1 gbuf_q_222(.A(q_in_222), .Y(Wt[14]));
CLKBUFX1 gbuf_d_223(.A(n4481), .Y(d_out_223));
CLKBUFX1 gbuf_q_223(.A(q_in_223), .Y(n14947));
CLKBUFX1 gbuf_d_224(.A(n4449), .Y(d_out_224));
CLKBUFX1 gbuf_q_224(.A(q_in_224), .Y(n15154));
CLKBUFX1 gbuf_qn_224(.A(qn_in_224), .Y(n8294));
CLKBUFX1 gbuf_d_225(.A(n4417), .Y(d_out_225));
CLKBUFX1 gbuf_q_225(.A(q_in_225), .Y(n15155));
CLKBUFX1 gbuf_d_226(.A(n4385), .Y(d_out_226));
CLKBUFX1 gbuf_q_226(.A(q_in_226), .Y(n15156));
CLKBUFX1 gbuf_d_227(.A(n4353), .Y(d_out_227));
CLKBUFX1 gbuf_q_227(.A(q_in_227), .Y(n15157));
CLKBUFX1 gbuf_d_228(.A(n4321), .Y(d_out_228));
CLKBUFX1 gbuf_q_228(.A(q_in_228), .Y(n15158));
CLKBUFX1 gbuf_d_229(.A(n4290), .Y(d_out_229));
CLKBUFX1 gbuf_q_229(.A(q_in_229), .Y(n15159));
CLKBUFX1 gbuf_d_230(.A(n4258), .Y(d_out_230));
CLKBUFX1 gbuf_q_230(.A(q_in_230), .Y(n15160));
CLKBUFX1 gbuf_d_231(.A(n4226), .Y(d_out_231));
CLKBUFX1 gbuf_q_231(.A(q_in_231), .Y(n15161));
CLKBUFX1 gbuf_d_232(.A(n4194), .Y(d_out_232));
CLKBUFX1 gbuf_q_232(.A(q_in_232), .Y(n15162));
CLKBUFX1 gbuf_d_233(.A(n4162), .Y(d_out_233));
CLKBUFX1 gbuf_q_233(.A(q_in_233), .Y(n15163));
CLKBUFX1 gbuf_d_234(.A(n4130), .Y(d_out_234));
CLKBUFX1 gbuf_q_234(.A(q_in_234), .Y(n15164));
CLKBUFX1 gbuf_d_235(.A(n4098), .Y(d_out_235));
CLKBUFX1 gbuf_q_235(.A(q_in_235), .Y(n15165));
CLKBUFX1 gbuf_qn_235(.A(qn_in_235), .Y(n12948));
CLKBUFX1 gbuf_d_236(.A(n4066), .Y(d_out_236));
CLKBUFX1 gbuf_q_236(.A(q_in_236), .Y(n15166));
CLKBUFX1 gbuf_d_237(.A(n4034), .Y(d_out_237));
CLKBUFX1 gbuf_q_237(.A(q_in_237), .Y(n15167));
CLKBUFX1 gbuf_d_238(.A(n4512), .Y(d_out_238));
CLKBUFX1 gbuf_q_238(.A(q_in_238), .Y(Wt[15]));
CLKBUFX1 gbuf_d_239(.A(n4480), .Y(d_out_239));
CLKBUFX1 gbuf_q_239(.A(q_in_239), .Y(n14948));
CLKBUFX1 gbuf_d_240(.A(n4448), .Y(d_out_240));
CLKBUFX1 gbuf_q_240(.A(q_in_240), .Y(n15168));
CLKBUFX1 gbuf_qn_240(.A(qn_in_240), .Y(n8292));
CLKBUFX1 gbuf_d_241(.A(n4416), .Y(d_out_241));
CLKBUFX1 gbuf_q_241(.A(q_in_241), .Y(n15169));
CLKBUFX1 gbuf_d_242(.A(n4384), .Y(d_out_242));
CLKBUFX1 gbuf_q_242(.A(q_in_242), .Y(n15170));
CLKBUFX1 gbuf_d_243(.A(n4352), .Y(d_out_243));
CLKBUFX1 gbuf_q_243(.A(q_in_243), .Y(n15171));
CLKBUFX1 gbuf_d_244(.A(n4320), .Y(d_out_244));
CLKBUFX1 gbuf_q_244(.A(q_in_244), .Y(n15172));
CLKBUFX1 gbuf_d_245(.A(n4289), .Y(d_out_245));
CLKBUFX1 gbuf_q_245(.A(q_in_245), .Y(n15173));
CLKBUFX1 gbuf_d_246(.A(n4257), .Y(d_out_246));
CLKBUFX1 gbuf_q_246(.A(q_in_246), .Y(n15174));
CLKBUFX1 gbuf_d_247(.A(n4225), .Y(d_out_247));
CLKBUFX1 gbuf_q_247(.A(q_in_247), .Y(n15175));
CLKBUFX1 gbuf_d_248(.A(n4193), .Y(d_out_248));
CLKBUFX1 gbuf_q_248(.A(q_in_248), .Y(n15176));
CLKBUFX1 gbuf_d_249(.A(n4161), .Y(d_out_249));
CLKBUFX1 gbuf_q_249(.A(q_in_249), .Y(n15177));
CLKBUFX1 gbuf_d_250(.A(n4129), .Y(d_out_250));
CLKBUFX1 gbuf_q_250(.A(q_in_250), .Y(n15178));
CLKBUFX1 gbuf_d_251(.A(n4097), .Y(d_out_251));
CLKBUFX1 gbuf_q_251(.A(q_in_251), .Y(n15179));
CLKBUFX1 gbuf_qn_251(.A(qn_in_251), .Y(n12946));
CLKBUFX1 gbuf_d_252(.A(n4065), .Y(d_out_252));
CLKBUFX1 gbuf_q_252(.A(q_in_252), .Y(n15180));
CLKBUFX1 gbuf_d_253(.A(n4033), .Y(d_out_253));
CLKBUFX1 gbuf_q_253(.A(q_in_253), .Y(n15181));
CLKBUFX1 gbuf_d_254(.A(n4511), .Y(d_out_254));
CLKBUFX1 gbuf_q_254(.A(q_in_254), .Y(Wt[16]));
CLKBUFX1 gbuf_d_255(.A(n4479), .Y(d_out_255));
CLKBUFX1 gbuf_q_255(.A(q_in_255), .Y(n14949));
CLKBUFX1 gbuf_d_256(.A(n4447), .Y(d_out_256));
CLKBUFX1 gbuf_q_256(.A(q_in_256), .Y(n15182));
CLKBUFX1 gbuf_qn_256(.A(qn_in_256), .Y(n8290));
CLKBUFX1 gbuf_d_257(.A(n4415), .Y(d_out_257));
CLKBUFX1 gbuf_q_257(.A(q_in_257), .Y(n15183));
CLKBUFX1 gbuf_d_258(.A(n4383), .Y(d_out_258));
CLKBUFX1 gbuf_q_258(.A(q_in_258), .Y(n15184));
CLKBUFX1 gbuf_d_259(.A(n4351), .Y(d_out_259));
CLKBUFX1 gbuf_q_259(.A(q_in_259), .Y(n15185));
CLKBUFX1 gbuf_d_260(.A(n4319), .Y(d_out_260));
CLKBUFX1 gbuf_q_260(.A(q_in_260), .Y(n15186));
CLKBUFX1 gbuf_d_261(.A(n4288), .Y(d_out_261));
CLKBUFX1 gbuf_q_261(.A(q_in_261), .Y(n15187));
CLKBUFX1 gbuf_d_262(.A(n4256), .Y(d_out_262));
CLKBUFX1 gbuf_q_262(.A(q_in_262), .Y(n15188));
CLKBUFX1 gbuf_d_263(.A(n4224), .Y(d_out_263));
CLKBUFX1 gbuf_q_263(.A(q_in_263), .Y(n15189));
CLKBUFX1 gbuf_d_264(.A(n4192), .Y(d_out_264));
CLKBUFX1 gbuf_q_264(.A(q_in_264), .Y(n15190));
CLKBUFX1 gbuf_d_265(.A(n4160), .Y(d_out_265));
CLKBUFX1 gbuf_q_265(.A(q_in_265), .Y(n15191));
CLKBUFX1 gbuf_d_266(.A(n4128), .Y(d_out_266));
CLKBUFX1 gbuf_q_266(.A(q_in_266), .Y(n15192));
CLKBUFX1 gbuf_d_267(.A(n4096), .Y(d_out_267));
CLKBUFX1 gbuf_q_267(.A(q_in_267), .Y(n15193));
CLKBUFX1 gbuf_qn_267(.A(qn_in_267), .Y(n12944));
CLKBUFX1 gbuf_d_268(.A(n4064), .Y(d_out_268));
CLKBUFX1 gbuf_q_268(.A(q_in_268), .Y(n15194));
CLKBUFX1 gbuf_d_269(.A(n4032), .Y(d_out_269));
CLKBUFX1 gbuf_q_269(.A(q_in_269), .Y(n15195));
CLKBUFX1 gbuf_d_270(.A(n4510), .Y(d_out_270));
CLKBUFX1 gbuf_q_270(.A(q_in_270), .Y(Wt[17]));
CLKBUFX1 gbuf_d_271(.A(n4478), .Y(d_out_271));
CLKBUFX1 gbuf_q_271(.A(q_in_271), .Y(n14950));
CLKBUFX1 gbuf_d_272(.A(n4446), .Y(d_out_272));
CLKBUFX1 gbuf_q_272(.A(q_in_272), .Y(n15196));
CLKBUFX1 gbuf_qn_272(.A(qn_in_272), .Y(n8288));
CLKBUFX1 gbuf_d_273(.A(n4414), .Y(d_out_273));
CLKBUFX1 gbuf_q_273(.A(q_in_273), .Y(n15197));
CLKBUFX1 gbuf_d_274(.A(n4382), .Y(d_out_274));
CLKBUFX1 gbuf_q_274(.A(q_in_274), .Y(n15198));
CLKBUFX1 gbuf_d_275(.A(n4350), .Y(d_out_275));
CLKBUFX1 gbuf_q_275(.A(q_in_275), .Y(n15199));
CLKBUFX1 gbuf_d_276(.A(n4318), .Y(d_out_276));
CLKBUFX1 gbuf_q_276(.A(q_in_276), .Y(n15200));
CLKBUFX1 gbuf_d_277(.A(n4287), .Y(d_out_277));
CLKBUFX1 gbuf_q_277(.A(q_in_277), .Y(n15201));
CLKBUFX1 gbuf_d_278(.A(n4255), .Y(d_out_278));
CLKBUFX1 gbuf_q_278(.A(q_in_278), .Y(n15202));
CLKBUFX1 gbuf_d_279(.A(n4223), .Y(d_out_279));
CLKBUFX1 gbuf_q_279(.A(q_in_279), .Y(n15203));
CLKBUFX1 gbuf_d_280(.A(n4191), .Y(d_out_280));
CLKBUFX1 gbuf_q_280(.A(q_in_280), .Y(n15204));
CLKBUFX1 gbuf_d_281(.A(n4159), .Y(d_out_281));
CLKBUFX1 gbuf_q_281(.A(q_in_281), .Y(n15205));
CLKBUFX1 gbuf_d_282(.A(n4127), .Y(d_out_282));
CLKBUFX1 gbuf_q_282(.A(q_in_282), .Y(n15206));
CLKBUFX1 gbuf_d_283(.A(n4095), .Y(d_out_283));
CLKBUFX1 gbuf_q_283(.A(q_in_283), .Y(n15207));
CLKBUFX1 gbuf_qn_283(.A(qn_in_283), .Y(n12942));
CLKBUFX1 gbuf_d_284(.A(n4063), .Y(d_out_284));
CLKBUFX1 gbuf_q_284(.A(q_in_284), .Y(n15208));
CLKBUFX1 gbuf_d_285(.A(n4031), .Y(d_out_285));
CLKBUFX1 gbuf_q_285(.A(q_in_285), .Y(n15209));
CLKBUFX1 gbuf_d_286(.A(n4509), .Y(d_out_286));
CLKBUFX1 gbuf_q_286(.A(q_in_286), .Y(Wt[18]));
CLKBUFX1 gbuf_d_287(.A(n4477), .Y(d_out_287));
CLKBUFX1 gbuf_q_287(.A(q_in_287), .Y(n15210));
CLKBUFX1 gbuf_d_288(.A(n4445), .Y(d_out_288));
CLKBUFX1 gbuf_q_288(.A(q_in_288), .Y(n15211));
CLKBUFX1 gbuf_qn_288(.A(qn_in_288), .Y(n8286));
CLKBUFX1 gbuf_d_289(.A(n4413), .Y(d_out_289));
CLKBUFX1 gbuf_q_289(.A(q_in_289), .Y(n15212));
CLKBUFX1 gbuf_d_290(.A(n4381), .Y(d_out_290));
CLKBUFX1 gbuf_q_290(.A(q_in_290), .Y(n15213));
CLKBUFX1 gbuf_d_291(.A(n4349), .Y(d_out_291));
CLKBUFX1 gbuf_q_291(.A(q_in_291), .Y(n15214));
CLKBUFX1 gbuf_d_292(.A(n4317), .Y(d_out_292));
CLKBUFX1 gbuf_q_292(.A(q_in_292), .Y(n15215));
CLKBUFX1 gbuf_d_293(.A(n4286), .Y(d_out_293));
CLKBUFX1 gbuf_q_293(.A(q_in_293), .Y(n15216));
CLKBUFX1 gbuf_d_294(.A(n4254), .Y(d_out_294));
CLKBUFX1 gbuf_q_294(.A(q_in_294), .Y(n15217));
CLKBUFX1 gbuf_d_295(.A(n4222), .Y(d_out_295));
CLKBUFX1 gbuf_q_295(.A(q_in_295), .Y(n15218));
CLKBUFX1 gbuf_d_296(.A(n4190), .Y(d_out_296));
CLKBUFX1 gbuf_q_296(.A(q_in_296), .Y(n15219));
CLKBUFX1 gbuf_d_297(.A(n4158), .Y(d_out_297));
CLKBUFX1 gbuf_q_297(.A(q_in_297), .Y(n15220));
CLKBUFX1 gbuf_d_298(.A(n4126), .Y(d_out_298));
CLKBUFX1 gbuf_q_298(.A(q_in_298), .Y(n15221));
CLKBUFX1 gbuf_d_299(.A(n4094), .Y(d_out_299));
CLKBUFX1 gbuf_q_299(.A(q_in_299), .Y(n15222));
CLKBUFX1 gbuf_qn_299(.A(qn_in_299), .Y(n12940));
CLKBUFX1 gbuf_d_300(.A(n4062), .Y(d_out_300));
CLKBUFX1 gbuf_q_300(.A(q_in_300), .Y(n15223));
CLKBUFX1 gbuf_d_301(.A(n4030), .Y(d_out_301));
CLKBUFX1 gbuf_q_301(.A(q_in_301), .Y(n15224));
CLKBUFX1 gbuf_d_302(.A(n4508), .Y(d_out_302));
CLKBUFX1 gbuf_q_302(.A(q_in_302), .Y(Wt[19]));
CLKBUFX1 gbuf_d_303(.A(n4476), .Y(d_out_303));
CLKBUFX1 gbuf_q_303(.A(q_in_303), .Y(n15225));
CLKBUFX1 gbuf_d_304(.A(n4444), .Y(d_out_304));
CLKBUFX1 gbuf_q_304(.A(q_in_304), .Y(n15226));
CLKBUFX1 gbuf_qn_304(.A(qn_in_304), .Y(n8284));
CLKBUFX1 gbuf_d_305(.A(n4412), .Y(d_out_305));
CLKBUFX1 gbuf_q_305(.A(q_in_305), .Y(n15227));
CLKBUFX1 gbuf_d_306(.A(n4380), .Y(d_out_306));
CLKBUFX1 gbuf_q_306(.A(q_in_306), .Y(n15228));
CLKBUFX1 gbuf_d_307(.A(n4348), .Y(d_out_307));
CLKBUFX1 gbuf_q_307(.A(q_in_307), .Y(n15229));
CLKBUFX1 gbuf_d_308(.A(n4316), .Y(d_out_308));
CLKBUFX1 gbuf_q_308(.A(q_in_308), .Y(n15230));
CLKBUFX1 gbuf_d_309(.A(n4285), .Y(d_out_309));
CLKBUFX1 gbuf_q_309(.A(q_in_309), .Y(n15231));
CLKBUFX1 gbuf_d_310(.A(n4253), .Y(d_out_310));
CLKBUFX1 gbuf_q_310(.A(q_in_310), .Y(n15232));
CLKBUFX1 gbuf_d_311(.A(n4221), .Y(d_out_311));
CLKBUFX1 gbuf_q_311(.A(q_in_311), .Y(n15233));
CLKBUFX1 gbuf_d_312(.A(n4189), .Y(d_out_312));
CLKBUFX1 gbuf_q_312(.A(q_in_312), .Y(n15234));
CLKBUFX1 gbuf_d_313(.A(n4157), .Y(d_out_313));
CLKBUFX1 gbuf_q_313(.A(q_in_313), .Y(n15235));
CLKBUFX1 gbuf_d_314(.A(n4125), .Y(d_out_314));
CLKBUFX1 gbuf_q_314(.A(q_in_314), .Y(n15236));
CLKBUFX1 gbuf_d_315(.A(n4093), .Y(d_out_315));
CLKBUFX1 gbuf_q_315(.A(q_in_315), .Y(n15237));
CLKBUFX1 gbuf_qn_315(.A(qn_in_315), .Y(n12938));
CLKBUFX1 gbuf_d_316(.A(n4061), .Y(d_out_316));
CLKBUFX1 gbuf_q_316(.A(q_in_316), .Y(n15238));
CLKBUFX1 gbuf_d_317(.A(n4029), .Y(d_out_317));
CLKBUFX1 gbuf_q_317(.A(q_in_317), .Y(n15239));
CLKBUFX1 gbuf_d_318(.A(n4507), .Y(d_out_318));
CLKBUFX1 gbuf_q_318(.A(q_in_318), .Y(Wt[20]));
CLKBUFX1 gbuf_d_319(.A(n4475), .Y(d_out_319));
CLKBUFX1 gbuf_q_319(.A(q_in_319), .Y(n15240));
CLKBUFX1 gbuf_d_320(.A(n4443), .Y(d_out_320));
CLKBUFX1 gbuf_q_320(.A(q_in_320), .Y(n15241));
CLKBUFX1 gbuf_qn_320(.A(qn_in_320), .Y(n8282));
CLKBUFX1 gbuf_d_321(.A(n4411), .Y(d_out_321));
CLKBUFX1 gbuf_q_321(.A(q_in_321), .Y(n15242));
CLKBUFX1 gbuf_d_322(.A(n4379), .Y(d_out_322));
CLKBUFX1 gbuf_q_322(.A(q_in_322), .Y(n15243));
CLKBUFX1 gbuf_d_323(.A(n4347), .Y(d_out_323));
CLKBUFX1 gbuf_q_323(.A(q_in_323), .Y(n15244));
CLKBUFX1 gbuf_d_324(.A(n4315), .Y(d_out_324));
CLKBUFX1 gbuf_q_324(.A(q_in_324), .Y(n15245));
CLKBUFX1 gbuf_d_325(.A(n4284), .Y(d_out_325));
CLKBUFX1 gbuf_q_325(.A(q_in_325), .Y(n15246));
CLKBUFX1 gbuf_d_326(.A(n4252), .Y(d_out_326));
CLKBUFX1 gbuf_q_326(.A(q_in_326), .Y(n15247));
CLKBUFX1 gbuf_d_327(.A(n4220), .Y(d_out_327));
CLKBUFX1 gbuf_q_327(.A(q_in_327), .Y(n15248));
CLKBUFX1 gbuf_d_328(.A(n4188), .Y(d_out_328));
CLKBUFX1 gbuf_q_328(.A(q_in_328), .Y(n15249));
CLKBUFX1 gbuf_d_329(.A(n4156), .Y(d_out_329));
CLKBUFX1 gbuf_q_329(.A(q_in_329), .Y(n15250));
CLKBUFX1 gbuf_d_330(.A(n4124), .Y(d_out_330));
CLKBUFX1 gbuf_q_330(.A(q_in_330), .Y(n15251));
CLKBUFX1 gbuf_d_331(.A(n4092), .Y(d_out_331));
CLKBUFX1 gbuf_q_331(.A(q_in_331), .Y(n15252));
CLKBUFX1 gbuf_qn_331(.A(qn_in_331), .Y(n12936));
CLKBUFX1 gbuf_d_332(.A(n4060), .Y(d_out_332));
CLKBUFX1 gbuf_q_332(.A(q_in_332), .Y(n15253));
CLKBUFX1 gbuf_d_333(.A(n4028), .Y(d_out_333));
CLKBUFX1 gbuf_q_333(.A(q_in_333), .Y(n15254));
CLKBUFX1 gbuf_d_334(.A(n4506), .Y(d_out_334));
CLKBUFX1 gbuf_q_334(.A(q_in_334), .Y(Wt[21]));
CLKBUFX1 gbuf_d_335(.A(n4474), .Y(d_out_335));
CLKBUFX1 gbuf_q_335(.A(q_in_335), .Y(n15255));
CLKBUFX1 gbuf_d_336(.A(n4442), .Y(d_out_336));
CLKBUFX1 gbuf_q_336(.A(q_in_336), .Y(n15256));
CLKBUFX1 gbuf_qn_336(.A(qn_in_336), .Y(n8280));
CLKBUFX1 gbuf_d_337(.A(n4410), .Y(d_out_337));
CLKBUFX1 gbuf_q_337(.A(q_in_337), .Y(n15257));
CLKBUFX1 gbuf_d_338(.A(n4378), .Y(d_out_338));
CLKBUFX1 gbuf_q_338(.A(q_in_338), .Y(n15258));
CLKBUFX1 gbuf_d_339(.A(n4346), .Y(d_out_339));
CLKBUFX1 gbuf_q_339(.A(q_in_339), .Y(n15259));
CLKBUFX1 gbuf_d_340(.A(n4314), .Y(d_out_340));
CLKBUFX1 gbuf_q_340(.A(q_in_340), .Y(n15260));
CLKBUFX1 gbuf_d_341(.A(n4283), .Y(d_out_341));
CLKBUFX1 gbuf_q_341(.A(q_in_341), .Y(n15261));
CLKBUFX1 gbuf_d_342(.A(n4251), .Y(d_out_342));
CLKBUFX1 gbuf_q_342(.A(q_in_342), .Y(n15262));
CLKBUFX1 gbuf_d_343(.A(n4219), .Y(d_out_343));
CLKBUFX1 gbuf_q_343(.A(q_in_343), .Y(n15263));
CLKBUFX1 gbuf_d_344(.A(n4187), .Y(d_out_344));
CLKBUFX1 gbuf_q_344(.A(q_in_344), .Y(n15264));
CLKBUFX1 gbuf_d_345(.A(n4155), .Y(d_out_345));
CLKBUFX1 gbuf_q_345(.A(q_in_345), .Y(n15265));
CLKBUFX1 gbuf_d_346(.A(n4123), .Y(d_out_346));
CLKBUFX1 gbuf_q_346(.A(q_in_346), .Y(n15266));
CLKBUFX1 gbuf_d_347(.A(n4091), .Y(d_out_347));
CLKBUFX1 gbuf_q_347(.A(q_in_347), .Y(n15267));
CLKBUFX1 gbuf_qn_347(.A(qn_in_347), .Y(n12934));
CLKBUFX1 gbuf_d_348(.A(n4059), .Y(d_out_348));
CLKBUFX1 gbuf_q_348(.A(q_in_348), .Y(n15268));
CLKBUFX1 gbuf_d_349(.A(n4027), .Y(d_out_349));
CLKBUFX1 gbuf_q_349(.A(q_in_349), .Y(n15269));
CLKBUFX1 gbuf_d_350(.A(n4505), .Y(d_out_350));
CLKBUFX1 gbuf_q_350(.A(q_in_350), .Y(Wt[22]));
CLKBUFX1 gbuf_d_351(.A(n4473), .Y(d_out_351));
CLKBUFX1 gbuf_q_351(.A(q_in_351), .Y(n15270));
CLKBUFX1 gbuf_d_352(.A(n4441), .Y(d_out_352));
CLKBUFX1 gbuf_q_352(.A(q_in_352), .Y(n15271));
CLKBUFX1 gbuf_qn_352(.A(qn_in_352), .Y(n8278));
CLKBUFX1 gbuf_d_353(.A(n4409), .Y(d_out_353));
CLKBUFX1 gbuf_q_353(.A(q_in_353), .Y(n15272));
CLKBUFX1 gbuf_d_354(.A(n4377), .Y(d_out_354));
CLKBUFX1 gbuf_q_354(.A(q_in_354), .Y(n15273));
CLKBUFX1 gbuf_d_355(.A(n4345), .Y(d_out_355));
CLKBUFX1 gbuf_q_355(.A(q_in_355), .Y(n15274));
CLKBUFX1 gbuf_d_356(.A(n4313), .Y(d_out_356));
CLKBUFX1 gbuf_q_356(.A(q_in_356), .Y(n15275));
CLKBUFX1 gbuf_d_357(.A(n4282), .Y(d_out_357));
CLKBUFX1 gbuf_q_357(.A(q_in_357), .Y(n15276));
CLKBUFX1 gbuf_d_358(.A(n4250), .Y(d_out_358));
CLKBUFX1 gbuf_q_358(.A(q_in_358), .Y(n15277));
CLKBUFX1 gbuf_d_359(.A(n4218), .Y(d_out_359));
CLKBUFX1 gbuf_q_359(.A(q_in_359), .Y(n15278));
CLKBUFX1 gbuf_d_360(.A(n4186), .Y(d_out_360));
CLKBUFX1 gbuf_q_360(.A(q_in_360), .Y(n15279));
CLKBUFX1 gbuf_d_361(.A(n4154), .Y(d_out_361));
CLKBUFX1 gbuf_q_361(.A(q_in_361), .Y(n15280));
CLKBUFX1 gbuf_d_362(.A(n4122), .Y(d_out_362));
CLKBUFX1 gbuf_q_362(.A(q_in_362), .Y(n15281));
CLKBUFX1 gbuf_d_363(.A(n4090), .Y(d_out_363));
CLKBUFX1 gbuf_q_363(.A(q_in_363), .Y(n15282));
CLKBUFX1 gbuf_qn_363(.A(qn_in_363), .Y(n12932));
CLKBUFX1 gbuf_d_364(.A(n4058), .Y(d_out_364));
CLKBUFX1 gbuf_q_364(.A(q_in_364), .Y(n15283));
CLKBUFX1 gbuf_d_365(.A(n4026), .Y(d_out_365));
CLKBUFX1 gbuf_q_365(.A(q_in_365), .Y(n15284));
CLKBUFX1 gbuf_d_366(.A(n4504), .Y(d_out_366));
CLKBUFX1 gbuf_q_366(.A(q_in_366), .Y(Wt[23]));
CLKBUFX1 gbuf_d_367(.A(n4472), .Y(d_out_367));
CLKBUFX1 gbuf_q_367(.A(q_in_367), .Y(n15285));
CLKBUFX1 gbuf_d_368(.A(n4440), .Y(d_out_368));
CLKBUFX1 gbuf_q_368(.A(q_in_368), .Y(n15286));
CLKBUFX1 gbuf_qn_368(.A(qn_in_368), .Y(n8276));
CLKBUFX1 gbuf_d_369(.A(n4408), .Y(d_out_369));
CLKBUFX1 gbuf_q_369(.A(q_in_369), .Y(n15287));
CLKBUFX1 gbuf_d_370(.A(n4376), .Y(d_out_370));
CLKBUFX1 gbuf_q_370(.A(q_in_370), .Y(n15288));
CLKBUFX1 gbuf_d_371(.A(n4344), .Y(d_out_371));
CLKBUFX1 gbuf_q_371(.A(q_in_371), .Y(n15289));
CLKBUFX1 gbuf_d_372(.A(n4312), .Y(d_out_372));
CLKBUFX1 gbuf_q_372(.A(q_in_372), .Y(n15290));
CLKBUFX1 gbuf_d_373(.A(n4281), .Y(d_out_373));
CLKBUFX1 gbuf_q_373(.A(q_in_373), .Y(n15291));
CLKBUFX1 gbuf_d_374(.A(n4249), .Y(d_out_374));
CLKBUFX1 gbuf_q_374(.A(q_in_374), .Y(n15292));
CLKBUFX1 gbuf_d_375(.A(n4217), .Y(d_out_375));
CLKBUFX1 gbuf_q_375(.A(q_in_375), .Y(n15293));
CLKBUFX1 gbuf_d_376(.A(n4185), .Y(d_out_376));
CLKBUFX1 gbuf_q_376(.A(q_in_376), .Y(n15294));
CLKBUFX1 gbuf_d_377(.A(n4153), .Y(d_out_377));
CLKBUFX1 gbuf_q_377(.A(q_in_377), .Y(n15295));
CLKBUFX1 gbuf_d_378(.A(n4121), .Y(d_out_378));
CLKBUFX1 gbuf_q_378(.A(q_in_378), .Y(n15296));
CLKBUFX1 gbuf_d_379(.A(n4089), .Y(d_out_379));
CLKBUFX1 gbuf_q_379(.A(q_in_379), .Y(n15297));
CLKBUFX1 gbuf_qn_379(.A(qn_in_379), .Y(n12930));
CLKBUFX1 gbuf_d_380(.A(n4057), .Y(d_out_380));
CLKBUFX1 gbuf_q_380(.A(q_in_380), .Y(n15298));
CLKBUFX1 gbuf_d_381(.A(n4025), .Y(d_out_381));
CLKBUFX1 gbuf_q_381(.A(q_in_381), .Y(n15299));
CLKBUFX1 gbuf_d_382(.A(n4503), .Y(d_out_382));
CLKBUFX1 gbuf_q_382(.A(q_in_382), .Y(Wt[24]));
CLKBUFX1 gbuf_d_383(.A(n4471), .Y(d_out_383));
CLKBUFX1 gbuf_q_383(.A(q_in_383), .Y(n15300));
CLKBUFX1 gbuf_d_384(.A(n4439), .Y(d_out_384));
CLKBUFX1 gbuf_q_384(.A(q_in_384), .Y(n15301));
CLKBUFX1 gbuf_qn_384(.A(qn_in_384), .Y(n8274));
CLKBUFX1 gbuf_d_385(.A(n4407), .Y(d_out_385));
CLKBUFX1 gbuf_q_385(.A(q_in_385), .Y(n15302));
CLKBUFX1 gbuf_d_386(.A(n4375), .Y(d_out_386));
CLKBUFX1 gbuf_q_386(.A(q_in_386), .Y(n15303));
CLKBUFX1 gbuf_d_387(.A(n4343), .Y(d_out_387));
CLKBUFX1 gbuf_q_387(.A(q_in_387), .Y(n15304));
CLKBUFX1 gbuf_d_388(.A(n4311), .Y(d_out_388));
CLKBUFX1 gbuf_q_388(.A(q_in_388), .Y(n15305));
CLKBUFX1 gbuf_d_389(.A(n4280), .Y(d_out_389));
CLKBUFX1 gbuf_q_389(.A(q_in_389), .Y(n15306));
CLKBUFX1 gbuf_d_390(.A(n4248), .Y(d_out_390));
CLKBUFX1 gbuf_q_390(.A(q_in_390), .Y(n15307));
CLKBUFX1 gbuf_d_391(.A(n4216), .Y(d_out_391));
CLKBUFX1 gbuf_q_391(.A(q_in_391), .Y(n15308));
CLKBUFX1 gbuf_d_392(.A(n4184), .Y(d_out_392));
CLKBUFX1 gbuf_q_392(.A(q_in_392), .Y(n15309));
CLKBUFX1 gbuf_d_393(.A(n4152), .Y(d_out_393));
CLKBUFX1 gbuf_q_393(.A(q_in_393), .Y(n15310));
CLKBUFX1 gbuf_d_394(.A(n4120), .Y(d_out_394));
CLKBUFX1 gbuf_q_394(.A(q_in_394), .Y(n15311));
CLKBUFX1 gbuf_d_395(.A(n4088), .Y(d_out_395));
CLKBUFX1 gbuf_q_395(.A(q_in_395), .Y(n15312));
CLKBUFX1 gbuf_qn_395(.A(qn_in_395), .Y(n12928));
CLKBUFX1 gbuf_d_396(.A(n4056), .Y(d_out_396));
CLKBUFX1 gbuf_q_396(.A(q_in_396), .Y(n15313));
CLKBUFX1 gbuf_d_397(.A(n4024), .Y(d_out_397));
CLKBUFX1 gbuf_q_397(.A(q_in_397), .Y(n15314));
CLKBUFX1 gbuf_d_398(.A(n4502), .Y(d_out_398));
CLKBUFX1 gbuf_q_398(.A(q_in_398), .Y(Wt[25]));
CLKBUFX1 gbuf_d_399(.A(n4470), .Y(d_out_399));
CLKBUFX1 gbuf_q_399(.A(q_in_399), .Y(n15315));
CLKBUFX1 gbuf_d_400(.A(n4438), .Y(d_out_400));
CLKBUFX1 gbuf_q_400(.A(q_in_400), .Y(n15316));
CLKBUFX1 gbuf_qn_400(.A(qn_in_400), .Y(n8272));
CLKBUFX1 gbuf_d_401(.A(n4406), .Y(d_out_401));
CLKBUFX1 gbuf_q_401(.A(q_in_401), .Y(n15317));
CLKBUFX1 gbuf_d_402(.A(n4374), .Y(d_out_402));
CLKBUFX1 gbuf_q_402(.A(q_in_402), .Y(n15318));
CLKBUFX1 gbuf_d_403(.A(n4342), .Y(d_out_403));
CLKBUFX1 gbuf_q_403(.A(q_in_403), .Y(n15319));
CLKBUFX1 gbuf_d_404(.A(n4310), .Y(d_out_404));
CLKBUFX1 gbuf_q_404(.A(q_in_404), .Y(n15320));
CLKBUFX1 gbuf_d_405(.A(n4279), .Y(d_out_405));
CLKBUFX1 gbuf_q_405(.A(q_in_405), .Y(n15321));
CLKBUFX1 gbuf_d_406(.A(n4247), .Y(d_out_406));
CLKBUFX1 gbuf_q_406(.A(q_in_406), .Y(n15322));
CLKBUFX1 gbuf_d_407(.A(n4215), .Y(d_out_407));
CLKBUFX1 gbuf_q_407(.A(q_in_407), .Y(n15323));
CLKBUFX1 gbuf_d_408(.A(n4183), .Y(d_out_408));
CLKBUFX1 gbuf_q_408(.A(q_in_408), .Y(n15324));
CLKBUFX1 gbuf_d_409(.A(n4151), .Y(d_out_409));
CLKBUFX1 gbuf_q_409(.A(q_in_409), .Y(n15325));
CLKBUFX1 gbuf_d_410(.A(n4119), .Y(d_out_410));
CLKBUFX1 gbuf_q_410(.A(q_in_410), .Y(n15326));
CLKBUFX1 gbuf_d_411(.A(n4087), .Y(d_out_411));
CLKBUFX1 gbuf_q_411(.A(q_in_411), .Y(n15327));
CLKBUFX1 gbuf_qn_411(.A(qn_in_411), .Y(n12926));
CLKBUFX1 gbuf_d_412(.A(n4055), .Y(d_out_412));
CLKBUFX1 gbuf_q_412(.A(q_in_412), .Y(n15328));
CLKBUFX1 gbuf_d_413(.A(n4023), .Y(d_out_413));
CLKBUFX1 gbuf_q_413(.A(q_in_413), .Y(n15329));
CLKBUFX1 gbuf_d_414(.A(n4501), .Y(d_out_414));
CLKBUFX1 gbuf_q_414(.A(q_in_414), .Y(Wt[26]));
CLKBUFX1 gbuf_d_415(.A(n4469), .Y(d_out_415));
CLKBUFX1 gbuf_q_415(.A(q_in_415), .Y(n15330));
CLKBUFX1 gbuf_d_416(.A(n4437), .Y(d_out_416));
CLKBUFX1 gbuf_q_416(.A(q_in_416), .Y(n15331));
CLKBUFX1 gbuf_qn_416(.A(qn_in_416), .Y(n8270));
CLKBUFX1 gbuf_d_417(.A(n4405), .Y(d_out_417));
CLKBUFX1 gbuf_q_417(.A(q_in_417), .Y(n15332));
CLKBUFX1 gbuf_d_418(.A(n4373), .Y(d_out_418));
CLKBUFX1 gbuf_q_418(.A(q_in_418), .Y(n15333));
CLKBUFX1 gbuf_d_419(.A(n4341), .Y(d_out_419));
CLKBUFX1 gbuf_q_419(.A(q_in_419), .Y(n15334));
CLKBUFX1 gbuf_d_420(.A(n4309), .Y(d_out_420));
CLKBUFX1 gbuf_q_420(.A(q_in_420), .Y(n15335));
CLKBUFX1 gbuf_d_421(.A(n4278), .Y(d_out_421));
CLKBUFX1 gbuf_q_421(.A(q_in_421), .Y(n15336));
CLKBUFX1 gbuf_d_422(.A(n4246), .Y(d_out_422));
CLKBUFX1 gbuf_q_422(.A(q_in_422), .Y(n15337));
CLKBUFX1 gbuf_d_423(.A(n4214), .Y(d_out_423));
CLKBUFX1 gbuf_q_423(.A(q_in_423), .Y(n15338));
CLKBUFX1 gbuf_d_424(.A(n4182), .Y(d_out_424));
CLKBUFX1 gbuf_q_424(.A(q_in_424), .Y(n15339));
CLKBUFX1 gbuf_d_425(.A(n4150), .Y(d_out_425));
CLKBUFX1 gbuf_q_425(.A(q_in_425), .Y(n15340));
CLKBUFX1 gbuf_d_426(.A(n4118), .Y(d_out_426));
CLKBUFX1 gbuf_q_426(.A(q_in_426), .Y(n15341));
CLKBUFX1 gbuf_d_427(.A(n4086), .Y(d_out_427));
CLKBUFX1 gbuf_q_427(.A(q_in_427), .Y(n15342));
CLKBUFX1 gbuf_qn_427(.A(qn_in_427), .Y(n12924));
CLKBUFX1 gbuf_d_428(.A(n4054), .Y(d_out_428));
CLKBUFX1 gbuf_q_428(.A(q_in_428), .Y(n15343));
CLKBUFX1 gbuf_d_429(.A(n4022), .Y(d_out_429));
CLKBUFX1 gbuf_q_429(.A(q_in_429), .Y(n15344));
CLKBUFX1 gbuf_d_430(.A(n4500), .Y(d_out_430));
CLKBUFX1 gbuf_q_430(.A(q_in_430), .Y(Wt[27]));
CLKBUFX1 gbuf_d_431(.A(n4468), .Y(d_out_431));
CLKBUFX1 gbuf_q_431(.A(q_in_431), .Y(n15345));
CLKBUFX1 gbuf_d_432(.A(n4436), .Y(d_out_432));
CLKBUFX1 gbuf_q_432(.A(q_in_432), .Y(n15346));
CLKBUFX1 gbuf_qn_432(.A(qn_in_432), .Y(n8268));
CLKBUFX1 gbuf_d_433(.A(n4404), .Y(d_out_433));
CLKBUFX1 gbuf_q_433(.A(q_in_433), .Y(n15347));
CLKBUFX1 gbuf_d_434(.A(n4372), .Y(d_out_434));
CLKBUFX1 gbuf_q_434(.A(q_in_434), .Y(n15348));
CLKBUFX1 gbuf_d_435(.A(n4340), .Y(d_out_435));
CLKBUFX1 gbuf_q_435(.A(q_in_435), .Y(n15349));
CLKBUFX1 gbuf_d_436(.A(n4308), .Y(d_out_436));
CLKBUFX1 gbuf_q_436(.A(q_in_436), .Y(n15350));
CLKBUFX1 gbuf_d_437(.A(n4277), .Y(d_out_437));
CLKBUFX1 gbuf_q_437(.A(q_in_437), .Y(n15351));
CLKBUFX1 gbuf_d_438(.A(n4245), .Y(d_out_438));
CLKBUFX1 gbuf_q_438(.A(q_in_438), .Y(n15352));
CLKBUFX1 gbuf_d_439(.A(n4213), .Y(d_out_439));
CLKBUFX1 gbuf_q_439(.A(q_in_439), .Y(n15353));
CLKBUFX1 gbuf_d_440(.A(n4181), .Y(d_out_440));
CLKBUFX1 gbuf_q_440(.A(q_in_440), .Y(n15354));
CLKBUFX1 gbuf_d_441(.A(n4149), .Y(d_out_441));
CLKBUFX1 gbuf_q_441(.A(q_in_441), .Y(n15355));
CLKBUFX1 gbuf_d_442(.A(n4117), .Y(d_out_442));
CLKBUFX1 gbuf_q_442(.A(q_in_442), .Y(n15356));
CLKBUFX1 gbuf_d_443(.A(n4085), .Y(d_out_443));
CLKBUFX1 gbuf_q_443(.A(q_in_443), .Y(n15357));
CLKBUFX1 gbuf_qn_443(.A(qn_in_443), .Y(n12922));
CLKBUFX1 gbuf_d_444(.A(n4053), .Y(d_out_444));
CLKBUFX1 gbuf_q_444(.A(q_in_444), .Y(n15358));
CLKBUFX1 gbuf_d_445(.A(n4021), .Y(d_out_445));
CLKBUFX1 gbuf_q_445(.A(q_in_445), .Y(n15359));
CLKBUFX1 gbuf_d_446(.A(n4499), .Y(d_out_446));
CLKBUFX1 gbuf_q_446(.A(q_in_446), .Y(Wt[28]));
CLKBUFX1 gbuf_d_447(.A(n4467), .Y(d_out_447));
CLKBUFX1 gbuf_q_447(.A(q_in_447), .Y(n15360));
CLKBUFX1 gbuf_d_448(.A(n4435), .Y(d_out_448));
CLKBUFX1 gbuf_q_448(.A(q_in_448), .Y(n15361));
CLKBUFX1 gbuf_qn_448(.A(qn_in_448), .Y(n8266));
CLKBUFX1 gbuf_d_449(.A(n4403), .Y(d_out_449));
CLKBUFX1 gbuf_q_449(.A(q_in_449), .Y(n15362));
CLKBUFX1 gbuf_d_450(.A(n4371), .Y(d_out_450));
CLKBUFX1 gbuf_q_450(.A(q_in_450), .Y(n15363));
CLKBUFX1 gbuf_d_451(.A(n4339), .Y(d_out_451));
CLKBUFX1 gbuf_q_451(.A(q_in_451), .Y(n15364));
CLKBUFX1 gbuf_d_452(.A(n4307), .Y(d_out_452));
CLKBUFX1 gbuf_q_452(.A(q_in_452), .Y(n15365));
CLKBUFX1 gbuf_d_453(.A(n4276), .Y(d_out_453));
CLKBUFX1 gbuf_q_453(.A(q_in_453), .Y(n15366));
CLKBUFX1 gbuf_d_454(.A(n4244), .Y(d_out_454));
CLKBUFX1 gbuf_q_454(.A(q_in_454), .Y(n15367));
CLKBUFX1 gbuf_d_455(.A(n4212), .Y(d_out_455));
CLKBUFX1 gbuf_q_455(.A(q_in_455), .Y(n15368));
CLKBUFX1 gbuf_d_456(.A(n4180), .Y(d_out_456));
CLKBUFX1 gbuf_q_456(.A(q_in_456), .Y(n15369));
CLKBUFX1 gbuf_d_457(.A(n4148), .Y(d_out_457));
CLKBUFX1 gbuf_q_457(.A(q_in_457), .Y(n15370));
CLKBUFX1 gbuf_d_458(.A(n4116), .Y(d_out_458));
CLKBUFX1 gbuf_q_458(.A(q_in_458), .Y(n15371));
CLKBUFX1 gbuf_d_459(.A(n4084), .Y(d_out_459));
CLKBUFX1 gbuf_q_459(.A(q_in_459), .Y(n15372));
CLKBUFX1 gbuf_qn_459(.A(qn_in_459), .Y(n12920));
CLKBUFX1 gbuf_d_460(.A(n4052), .Y(d_out_460));
CLKBUFX1 gbuf_q_460(.A(q_in_460), .Y(n15373));
CLKBUFX1 gbuf_d_461(.A(n4020), .Y(d_out_461));
CLKBUFX1 gbuf_q_461(.A(q_in_461), .Y(n15374));
CLKBUFX1 gbuf_d_462(.A(n4498), .Y(d_out_462));
CLKBUFX1 gbuf_q_462(.A(q_in_462), .Y(Wt[29]));
CLKBUFX1 gbuf_d_463(.A(n4466), .Y(d_out_463));
CLKBUFX1 gbuf_q_463(.A(q_in_463), .Y(n15375));
CLKBUFX1 gbuf_d_464(.A(n4434), .Y(d_out_464));
CLKBUFX1 gbuf_q_464(.A(q_in_464), .Y(n15376));
CLKBUFX1 gbuf_qn_464(.A(qn_in_464), .Y(n8264));
CLKBUFX1 gbuf_d_465(.A(n4402), .Y(d_out_465));
CLKBUFX1 gbuf_q_465(.A(q_in_465), .Y(n15377));
CLKBUFX1 gbuf_d_466(.A(n4370), .Y(d_out_466));
CLKBUFX1 gbuf_q_466(.A(q_in_466), .Y(n15378));
CLKBUFX1 gbuf_d_467(.A(n4338), .Y(d_out_467));
CLKBUFX1 gbuf_q_467(.A(q_in_467), .Y(n15379));
CLKBUFX1 gbuf_d_468(.A(n4306), .Y(d_out_468));
CLKBUFX1 gbuf_q_468(.A(q_in_468), .Y(n15380));
CLKBUFX1 gbuf_d_469(.A(n4275), .Y(d_out_469));
CLKBUFX1 gbuf_q_469(.A(q_in_469), .Y(n15381));
CLKBUFX1 gbuf_d_470(.A(n4243), .Y(d_out_470));
CLKBUFX1 gbuf_q_470(.A(q_in_470), .Y(n15382));
CLKBUFX1 gbuf_d_471(.A(n4211), .Y(d_out_471));
CLKBUFX1 gbuf_q_471(.A(q_in_471), .Y(n15383));
CLKBUFX1 gbuf_d_472(.A(n4179), .Y(d_out_472));
CLKBUFX1 gbuf_q_472(.A(q_in_472), .Y(n15384));
CLKBUFX1 gbuf_d_473(.A(n4147), .Y(d_out_473));
CLKBUFX1 gbuf_q_473(.A(q_in_473), .Y(n15385));
CLKBUFX1 gbuf_d_474(.A(n4115), .Y(d_out_474));
CLKBUFX1 gbuf_q_474(.A(q_in_474), .Y(n15386));
CLKBUFX1 gbuf_d_475(.A(n4083), .Y(d_out_475));
CLKBUFX1 gbuf_q_475(.A(q_in_475), .Y(n15387));
CLKBUFX1 gbuf_qn_475(.A(qn_in_475), .Y(n12918));
CLKBUFX1 gbuf_d_476(.A(n4051), .Y(d_out_476));
CLKBUFX1 gbuf_q_476(.A(q_in_476), .Y(n15388));
CLKBUFX1 gbuf_d_477(.A(n4019), .Y(d_out_477));
CLKBUFX1 gbuf_q_477(.A(q_in_477), .Y(n15389));
CLKBUFX1 gbuf_d_478(.A(n4497), .Y(d_out_478));
CLKBUFX1 gbuf_q_478(.A(q_in_478), .Y(Wt[30]));
CLKBUFX1 gbuf_d_479(.A(n4465), .Y(d_out_479));
CLKBUFX1 gbuf_q_479(.A(q_in_479), .Y(n15390));
CLKBUFX1 gbuf_d_480(.A(n4433), .Y(d_out_480));
CLKBUFX1 gbuf_q_480(.A(q_in_480), .Y(n15391));
CLKBUFX1 gbuf_qn_480(.A(qn_in_480), .Y(n8262));
CLKBUFX1 gbuf_d_481(.A(n4401), .Y(d_out_481));
CLKBUFX1 gbuf_q_481(.A(q_in_481), .Y(n15392));
CLKBUFX1 gbuf_d_482(.A(n4369), .Y(d_out_482));
CLKBUFX1 gbuf_q_482(.A(q_in_482), .Y(n15393));
CLKBUFX1 gbuf_d_483(.A(n4337), .Y(d_out_483));
CLKBUFX1 gbuf_q_483(.A(q_in_483), .Y(n15394));
CLKBUFX1 gbuf_d_484(.A(n4305), .Y(d_out_484));
CLKBUFX1 gbuf_q_484(.A(q_in_484), .Y(n15395));
CLKBUFX1 gbuf_d_485(.A(n4274), .Y(d_out_485));
CLKBUFX1 gbuf_q_485(.A(q_in_485), .Y(n15396));
CLKBUFX1 gbuf_d_486(.A(n4242), .Y(d_out_486));
CLKBUFX1 gbuf_q_486(.A(q_in_486), .Y(n15397));
CLKBUFX1 gbuf_d_487(.A(n4210), .Y(d_out_487));
CLKBUFX1 gbuf_q_487(.A(q_in_487), .Y(n15398));
CLKBUFX1 gbuf_d_488(.A(n4178), .Y(d_out_488));
CLKBUFX1 gbuf_q_488(.A(q_in_488), .Y(n15399));
CLKBUFX1 gbuf_d_489(.A(n4146), .Y(d_out_489));
CLKBUFX1 gbuf_q_489(.A(q_in_489), .Y(n15400));
CLKBUFX1 gbuf_d_490(.A(n4114), .Y(d_out_490));
CLKBUFX1 gbuf_q_490(.A(q_in_490), .Y(n15401));
CLKBUFX1 gbuf_d_491(.A(n4082), .Y(d_out_491));
CLKBUFX1 gbuf_q_491(.A(q_in_491), .Y(n15402));
CLKBUFX1 gbuf_qn_491(.A(qn_in_491), .Y(n12916));
CLKBUFX1 gbuf_d_492(.A(n4050), .Y(d_out_492));
CLKBUFX1 gbuf_q_492(.A(q_in_492), .Y(n15403));
CLKBUFX1 gbuf_d_493(.A(n4018), .Y(d_out_493));
CLKBUFX1 gbuf_q_493(.A(q_in_493), .Y(n15404));
CLKBUFX1 gbuf_d_494(.A(n4496), .Y(d_out_494));
CLKBUFX1 gbuf_q_494(.A(q_in_494), .Y(Wt[31]));
CLKBUFX1 gbuf_d_495(.A(n4464), .Y(d_out_495));
CLKBUFX1 gbuf_q_495(.A(q_in_495), .Y(n15405));
CLKBUFX1 gbuf_d_496(.A(n4432), .Y(d_out_496));
CLKBUFX1 gbuf_q_496(.A(q_in_496), .Y(n15406));
CLKBUFX1 gbuf_qn_496(.A(qn_in_496), .Y(n8323));
CLKBUFX1 gbuf_d_497(.A(n4400), .Y(d_out_497));
CLKBUFX1 gbuf_q_497(.A(q_in_497), .Y(n15407));
CLKBUFX1 gbuf_d_498(.A(n4368), .Y(d_out_498));
CLKBUFX1 gbuf_q_498(.A(q_in_498), .Y(n15408));
CLKBUFX1 gbuf_d_499(.A(n4336), .Y(d_out_499));
CLKBUFX1 gbuf_q_499(.A(q_in_499), .Y(n15409));
CLKBUFX1 gbuf_d_500(.A(n4304), .Y(d_out_500));
CLKBUFX1 gbuf_q_500(.A(q_in_500), .Y(n15410));
CLKBUFX1 gbuf_d_501(.A(n4273), .Y(d_out_501));
CLKBUFX1 gbuf_q_501(.A(q_in_501), .Y(n15411));
CLKBUFX1 gbuf_d_502(.A(n4241), .Y(d_out_502));
CLKBUFX1 gbuf_q_502(.A(q_in_502), .Y(n15412));
CLKBUFX1 gbuf_d_503(.A(n4209), .Y(d_out_503));
CLKBUFX1 gbuf_q_503(.A(q_in_503), .Y(n15413));
CLKBUFX1 gbuf_d_504(.A(n4177), .Y(d_out_504));
CLKBUFX1 gbuf_q_504(.A(q_in_504), .Y(n15414));
CLKBUFX1 gbuf_d_505(.A(n4145), .Y(d_out_505));
CLKBUFX1 gbuf_q_505(.A(q_in_505), .Y(n15415));
CLKBUFX1 gbuf_d_506(.A(n4113), .Y(d_out_506));
CLKBUFX1 gbuf_q_506(.A(q_in_506), .Y(n15416));
CLKBUFX1 gbuf_d_507(.A(n4081), .Y(d_out_507));
CLKBUFX1 gbuf_q_507(.A(q_in_507), .Y(n15417));
CLKBUFX1 gbuf_qn_507(.A(qn_in_507), .Y(n12978));
CLKBUFX1 gbuf_d_508(.A(n4049), .Y(d_out_508));
CLKBUFX1 gbuf_q_508(.A(q_in_508), .Y(n15418));
CLKBUFX1 gbuf_d_509(.A(n4017), .Y(d_out_509));
CLKBUFX1 gbuf_q_509(.A(q_in_509), .Y(n15419));
CLKBUFX1 gbuf_d_510(.A(n4527), .Y(d_out_510));
CLKBUFX1 gbuf_q_510(.A(q_in_510), .Y(Wt[0]));
CLKBUFX1 gbuf_d_511(.A(n4495), .Y(d_out_511));
CLKBUFX1 gbuf_q_511(.A(q_in_511), .Y(n14951));
CLKBUFX1 gbuf_d_512(.A(n4463), .Y(d_out_512));
CLKBUFX1 gbuf_q_512(.A(q_in_512), .Y(n15420));
CLKBUFX1 gbuf_qn_512(.A(qn_in_512), .Y(n8322));
CLKBUFX1 gbuf_d_513(.A(n4431), .Y(d_out_513));
CLKBUFX1 gbuf_q_513(.A(q_in_513), .Y(n15421));
CLKBUFX1 gbuf_d_514(.A(n4399), .Y(d_out_514));
CLKBUFX1 gbuf_q_514(.A(q_in_514), .Y(n15422));
CLKBUFX1 gbuf_d_515(.A(n4367), .Y(d_out_515));
CLKBUFX1 gbuf_q_515(.A(q_in_515), .Y(n15423));
CLKBUFX1 gbuf_d_516(.A(n4335), .Y(d_out_516));
CLKBUFX1 gbuf_q_516(.A(q_in_516), .Y(n15424));
CLKBUFX1 gbuf_d_517(.A(n3953), .Y(d_out_517));
CLKBUFX1 gbuf_q_517(.A(q_in_517), .Y(H0[31]));
CLKBUFX1 gbuf_d_518(.A(n4016), .Y(d_out_518));
CLKBUFX1 gbuf_q_518(.A(q_in_518), .Y(SHA1_result_128));
CLKBUFX1 gbuf_qn_518(.A(qn_in_518), .Y(n12851));
CLKBUFX1 gbuf_d_519(.A(n4015), .Y(d_out_519));
CLKBUFX1 gbuf_q_519(.A(q_in_519), .Y(SHA1_result_129));
CLKBUFX1 gbuf_qn_519(.A(qn_in_519), .Y(n12853));
CLKBUFX1 gbuf_d_520(.A(n3983), .Y(d_out_520));
CLKBUFX1 gbuf_q_520(.A(q_in_520), .Y(H0[1]));
CLKBUFX1 gbuf_d_521(.A(n4014), .Y(d_out_521));
CLKBUFX1 gbuf_q_521(.A(q_in_521), .Y(SHA1_result_130));
CLKBUFX1 gbuf_qn_521(.A(qn_in_521), .Y(n12855));
CLKBUFX1 gbuf_d_522(.A(n3982), .Y(d_out_522));
CLKBUFX1 gbuf_q_522(.A(q_in_522), .Y(H0[2]));
CLKBUFX1 gbuf_d_523(.A(n4013), .Y(d_out_523));
CLKBUFX1 gbuf_q_523(.A(q_in_523), .Y(SHA1_result_131));
CLKBUFX1 gbuf_qn_523(.A(qn_in_523), .Y(n12857));
CLKBUFX1 gbuf_d_524(.A(n3981), .Y(d_out_524));
CLKBUFX1 gbuf_q_524(.A(q_in_524), .Y(H0[3]));
CLKBUFX1 gbuf_d_525(.A(n4012), .Y(d_out_525));
CLKBUFX1 gbuf_q_525(.A(q_in_525), .Y(SHA1_result_132));
CLKBUFX1 gbuf_qn_525(.A(qn_in_525), .Y(n12859));
CLKBUFX1 gbuf_d_526(.A(n3980), .Y(d_out_526));
CLKBUFX1 gbuf_q_526(.A(q_in_526), .Y(H0[4]));
CLKBUFX1 gbuf_d_527(.A(n4011), .Y(d_out_527));
CLKBUFX1 gbuf_q_527(.A(q_in_527), .Y(SHA1_result_133));
CLKBUFX1 gbuf_qn_527(.A(qn_in_527), .Y(n12861));
CLKBUFX1 gbuf_d_528(.A(n3979), .Y(d_out_528));
CLKBUFX1 gbuf_q_528(.A(q_in_528), .Y(H0[5]));
CLKBUFX1 gbuf_d_529(.A(n4010), .Y(d_out_529));
CLKBUFX1 gbuf_q_529(.A(q_in_529), .Y(SHA1_result_134));
CLKBUFX1 gbuf_qn_529(.A(qn_in_529), .Y(n12863));
CLKBUFX1 gbuf_d_530(.A(n3978), .Y(d_out_530));
CLKBUFX1 gbuf_q_530(.A(q_in_530), .Y(H0[6]));
CLKBUFX1 gbuf_d_531(.A(n4009), .Y(d_out_531));
CLKBUFX1 gbuf_q_531(.A(q_in_531), .Y(SHA1_result_135));
CLKBUFX1 gbuf_qn_531(.A(qn_in_531), .Y(n12865));
CLKBUFX1 gbuf_d_532(.A(n3977), .Y(d_out_532));
CLKBUFX1 gbuf_q_532(.A(q_in_532), .Y(H0[7]));
CLKBUFX1 gbuf_d_533(.A(n4008), .Y(d_out_533));
CLKBUFX1 gbuf_q_533(.A(q_in_533), .Y(SHA1_result_136));
CLKBUFX1 gbuf_qn_533(.A(qn_in_533), .Y(n12867));
CLKBUFX1 gbuf_d_534(.A(n3976), .Y(d_out_534));
CLKBUFX1 gbuf_q_534(.A(q_in_534), .Y(H0[8]));
CLKBUFX1 gbuf_d_535(.A(n3975), .Y(d_out_535));
CLKBUFX1 gbuf_q_535(.A(q_in_535), .Y(H0[9]));
CLKBUFX1 gbuf_d_536(.A(n4006), .Y(d_out_536));
CLKBUFX1 gbuf_q_536(.A(q_in_536), .Y(n14440));
CLKBUFX1 gbuf_qn_536(.A(qn_in_536), .Y(n12871));
CLKBUFX1 gbuf_d_537(.A(n3974), .Y(d_out_537));
CLKBUFX1 gbuf_q_537(.A(q_in_537), .Y(H0[10]));
CLKBUFX1 gbuf_d_538(.A(n3973), .Y(d_out_538));
CLKBUFX1 gbuf_q_538(.A(q_in_538), .Y(H0[11]));
CLKBUFX1 gbuf_d_539(.A(n3972), .Y(d_out_539));
CLKBUFX1 gbuf_q_539(.A(q_in_539), .Y(H0[12]));
CLKBUFX1 gbuf_d_540(.A(n3971), .Y(d_out_540));
CLKBUFX1 gbuf_q_540(.A(q_in_540), .Y(H0[13]));
CLKBUFX1 gbuf_d_541(.A(n3970), .Y(d_out_541));
CLKBUFX1 gbuf_q_541(.A(q_in_541), .Y(H0[14]));
CLKBUFX1 gbuf_d_542(.A(n3969), .Y(d_out_542));
CLKBUFX1 gbuf_q_542(.A(q_in_542), .Y(H0[15]));
CLKBUFX1 gbuf_d_543(.A(n3968), .Y(d_out_543));
CLKBUFX1 gbuf_q_543(.A(q_in_543), .Y(H0[16]));
CLKBUFX1 gbuf_d_544(.A(n3967), .Y(d_out_544));
CLKBUFX1 gbuf_q_544(.A(q_in_544), .Y(H0[17]));
CLKBUFX1 gbuf_d_545(.A(n3966), .Y(d_out_545));
CLKBUFX1 gbuf_q_545(.A(q_in_545), .Y(H0[18]));
CLKBUFX1 gbuf_d_546(.A(n3965), .Y(d_out_546));
CLKBUFX1 gbuf_q_546(.A(q_in_546), .Y(H0[19]));
CLKBUFX1 gbuf_d_547(.A(n3996), .Y(d_out_547));
CLKBUFX1 gbuf_q_547(.A(q_in_547), .Y(SHA1_result_148));
CLKBUFX1 gbuf_qn_547(.A(qn_in_547), .Y(n12891));
CLKBUFX1 gbuf_d_548(.A(n3964), .Y(d_out_548));
CLKBUFX1 gbuf_q_548(.A(q_in_548), .Y(H0[20]));
CLKBUFX1 gbuf_d_549(.A(n3963), .Y(d_out_549));
CLKBUFX1 gbuf_q_549(.A(q_in_549), .Y(H0[21]));
CLKBUFX1 gbuf_d_550(.A(n3962), .Y(d_out_550));
CLKBUFX1 gbuf_q_550(.A(q_in_550), .Y(H0[22]));
CLKBUFX1 gbuf_d_551(.A(n3961), .Y(d_out_551));
CLKBUFX1 gbuf_q_551(.A(q_in_551), .Y(H0[23]));
CLKBUFX1 gbuf_d_552(.A(n3960), .Y(d_out_552));
CLKBUFX1 gbuf_q_552(.A(q_in_552), .Y(H0[24]));
CLKBUFX1 gbuf_d_553(.A(n3959), .Y(d_out_553));
CLKBUFX1 gbuf_q_553(.A(q_in_553), .Y(H0[25]));
CLKBUFX1 gbuf_d_554(.A(n3958), .Y(d_out_554));
CLKBUFX1 gbuf_q_554(.A(q_in_554), .Y(H0[26]));
CLKBUFX1 gbuf_d_555(.A(n3957), .Y(d_out_555));
CLKBUFX1 gbuf_q_555(.A(q_in_555), .Y(H0[27]));
CLKBUFX1 gbuf_d_556(.A(n3956), .Y(d_out_556));
CLKBUFX1 gbuf_q_556(.A(q_in_556), .Y(H0[28]));
CLKBUFX1 gbuf_d_557(.A(n3955), .Y(d_out_557));
CLKBUFX1 gbuf_q_557(.A(q_in_557), .Y(H0[29]));
CLKBUFX1 gbuf_d_558(.A(n3922), .Y(d_out_558));
CLKBUFX1 gbuf_q_558(.A(q_in_558), .Y(next_C[28]));
CLKBUFX1 gbuf_qn_558(.A(qn_in_558), .Y(n13007));
CLKBUFX1 gbuf_d_559(.A(n3698), .Y(d_out_559));
CLKBUFX1 gbuf_q_559(.A(q_in_559), .Y(H1[30]));
CLKBUFX1 gbuf_d_560(.A(n3952), .Y(d_out_560));
CLKBUFX1 gbuf_q_560(.A(q_in_560), .Y(next_C[30]));
CLKBUFX1 gbuf_qn_560(.A(qn_in_560), .Y(n13084));
CLKBUFX1 gbuf_d_561(.A(n3728), .Y(d_out_561));
CLKBUFX1 gbuf_q_561(.A(q_in_561), .Y(H1[0]));
CLKBUFX1 gbuf_d_562(.A(n3727), .Y(d_out_562));
CLKBUFX1 gbuf_q_562(.A(q_in_562), .Y(H1[1]));
CLKBUFX1 gbuf_d_563(.A(n3950), .Y(d_out_563));
CLKBUFX1 gbuf_q_563(.A(q_in_563), .Y(next_C[0]));
CLKBUFX1 gbuf_qn_563(.A(qn_in_563), .Y(n13083));
CLKBUFX1 gbuf_d_564(.A(n3726), .Y(d_out_564));
CLKBUFX1 gbuf_q_564(.A(q_in_564), .Y(H1[2]));
CLKBUFX1 gbuf_d_565(.A(n3725), .Y(d_out_565));
CLKBUFX1 gbuf_q_565(.A(q_in_565), .Y(H1[3]));
CLKBUFX1 gbuf_d_566(.A(n3948), .Y(d_out_566));
CLKBUFX1 gbuf_q_566(.A(q_in_566), .Y(next_C[2]));
CLKBUFX1 gbuf_qn_566(.A(qn_in_566), .Y(n13015));
CLKBUFX1 gbuf_d_567(.A(n3724), .Y(d_out_567));
CLKBUFX1 gbuf_q_567(.A(q_in_567), .Y(H1[4]));
CLKBUFX1 gbuf_d_568(.A(n3723), .Y(d_out_568));
CLKBUFX1 gbuf_q_568(.A(q_in_568), .Y(H1[5]));
CLKBUFX1 gbuf_d_569(.A(n3946), .Y(d_out_569));
CLKBUFX1 gbuf_q_569(.A(q_in_569), .Y(next_C[4]));
CLKBUFX1 gbuf_qn_569(.A(qn_in_569), .Y(n13000));
CLKBUFX1 gbuf_d_570(.A(n3722), .Y(d_out_570));
CLKBUFX1 gbuf_q_570(.A(q_in_570), .Y(H1[6]));
CLKBUFX1 gbuf_d_571(.A(n3945), .Y(d_out_571));
CLKBUFX1 gbuf_q_571(.A(q_in_571), .Y(next_C[5]));
CLKBUFX1 gbuf_qn_571(.A(qn_in_571), .Y(n13019));
CLKBUFX1 gbuf_d_572(.A(n3721), .Y(d_out_572));
CLKBUFX1 gbuf_q_572(.A(q_in_572), .Y(H1[7]));
CLKBUFX1 gbuf_d_573(.A(n3944), .Y(d_out_573));
CLKBUFX1 gbuf_q_573(.A(q_in_573), .Y(next_C[6]));
CLKBUFX1 gbuf_qn_573(.A(qn_in_573), .Y(n13020));
CLKBUFX1 gbuf_d_574(.A(n3720), .Y(d_out_574));
CLKBUFX1 gbuf_q_574(.A(q_in_574), .Y(H1[8]));
CLKBUFX1 gbuf_d_575(.A(n3943), .Y(d_out_575));
CLKBUFX1 gbuf_q_575(.A(q_in_575), .Y(next_C[7]));
CLKBUFX1 gbuf_qn_575(.A(qn_in_575), .Y(n13079));
CLKBUFX1 gbuf_d_576(.A(n3719), .Y(d_out_576));
CLKBUFX1 gbuf_q_576(.A(q_in_576), .Y(H1[9]));
CLKBUFX1 gbuf_d_577(.A(n3942), .Y(d_out_577));
CLKBUFX1 gbuf_q_577(.A(q_in_577), .Y(next_C[8]));
CLKBUFX1 gbuf_qn_577(.A(qn_in_577), .Y(n13098));
CLKBUFX1 gbuf_d_578(.A(n3718), .Y(d_out_578));
CLKBUFX1 gbuf_q_578(.A(q_in_578), .Y(H1[10]));
CLKBUFX1 gbuf_d_579(.A(n3941), .Y(d_out_579));
CLKBUFX1 gbuf_q_579(.A(q_in_579), .Y(next_C[9]));
CLKBUFX1 gbuf_qn_579(.A(qn_in_579), .Y(n13001));
CLKBUFX1 gbuf_d_580(.A(n3717), .Y(d_out_580));
CLKBUFX1 gbuf_q_580(.A(q_in_580), .Y(H1[11]));
CLKBUFX1 gbuf_d_581(.A(n3940), .Y(d_out_581));
CLKBUFX1 gbuf_q_581(.A(q_in_581), .Y(next_C[10]));
CLKBUFX1 gbuf_qn_581(.A(qn_in_581), .Y(n13016));
CLKBUFX1 gbuf_d_582(.A(n3716), .Y(d_out_582));
CLKBUFX1 gbuf_q_582(.A(q_in_582), .Y(H1[12]));
CLKBUFX1 gbuf_d_583(.A(n3939), .Y(d_out_583));
CLKBUFX1 gbuf_q_583(.A(q_in_583), .Y(next_C[11]));
CLKBUFX1 gbuf_qn_583(.A(qn_in_583), .Y(n13022));
CLKBUFX1 gbuf_d_584(.A(n3715), .Y(d_out_584));
CLKBUFX1 gbuf_q_584(.A(q_in_584), .Y(H1[13]));
CLKBUFX1 gbuf_d_585(.A(n3938), .Y(d_out_585));
CLKBUFX1 gbuf_q_585(.A(q_in_585), .Y(next_C[12]));
CLKBUFX1 gbuf_qn_585(.A(qn_in_585), .Y(n13005));
CLKBUFX1 gbuf_d_586(.A(n3714), .Y(d_out_586));
CLKBUFX1 gbuf_q_586(.A(q_in_586), .Y(H1[14]));
CLKBUFX1 gbuf_d_587(.A(n3937), .Y(d_out_587));
CLKBUFX1 gbuf_q_587(.A(q_in_587), .Y(next_C[13]));
CLKBUFX1 gbuf_qn_587(.A(qn_in_587), .Y(n13021));
CLKBUFX1 gbuf_d_588(.A(n3713), .Y(d_out_588));
CLKBUFX1 gbuf_q_588(.A(q_in_588), .Y(H1[15]));
CLKBUFX1 gbuf_d_589(.A(n3936), .Y(d_out_589));
CLKBUFX1 gbuf_q_589(.A(q_in_589), .Y(next_C[14]));
CLKBUFX1 gbuf_qn_589(.A(qn_in_589), .Y(n13018));
CLKBUFX1 gbuf_d_590(.A(n3712), .Y(d_out_590));
CLKBUFX1 gbuf_q_590(.A(q_in_590), .Y(H1[16]));
CLKBUFX1 gbuf_d_591(.A(n3935), .Y(d_out_591));
CLKBUFX1 gbuf_q_591(.A(q_in_591), .Y(next_C[15]));
CLKBUFX1 gbuf_qn_591(.A(qn_in_591), .Y(n13023));
CLKBUFX1 gbuf_d_592(.A(n3711), .Y(d_out_592));
CLKBUFX1 gbuf_q_592(.A(q_in_592), .Y(H1[17]));
CLKBUFX1 gbuf_d_593(.A(n3934), .Y(d_out_593));
CLKBUFX1 gbuf_q_593(.A(q_in_593), .Y(next_C[16]));
CLKBUFX1 gbuf_qn_593(.A(qn_in_593), .Y(n13004));
CLKBUFX1 gbuf_d_594(.A(n3710), .Y(d_out_594));
CLKBUFX1 gbuf_q_594(.A(q_in_594), .Y(H1[18]));
CLKBUFX1 gbuf_d_595(.A(n3709), .Y(d_out_595));
CLKBUFX1 gbuf_q_595(.A(q_in_595), .Y(H1[19]));
CLKBUFX1 gbuf_d_596(.A(n3932), .Y(d_out_596));
CLKBUFX1 gbuf_q_596(.A(q_in_596), .Y(next_C[18]));
CLKBUFX1 gbuf_qn_596(.A(qn_in_596), .Y(n13012));
CLKBUFX1 gbuf_d_597(.A(n3708), .Y(d_out_597));
CLKBUFX1 gbuf_q_597(.A(q_in_597), .Y(H1[20]));
CLKBUFX1 gbuf_d_598(.A(n3931), .Y(d_out_598));
CLKBUFX1 gbuf_q_598(.A(q_in_598), .Y(next_C[19]));
CLKBUFX1 gbuf_qn_598(.A(qn_in_598), .Y(n13011));
CLKBUFX1 gbuf_d_599(.A(n3707), .Y(d_out_599));
CLKBUFX1 gbuf_q_599(.A(q_in_599), .Y(H1[21]));
CLKBUFX1 gbuf_d_600(.A(n3930), .Y(d_out_600));
CLKBUFX1 gbuf_q_600(.A(q_in_600), .Y(next_C[20]));
CLKBUFX1 gbuf_qn_600(.A(qn_in_600), .Y(n13006));
CLKBUFX1 gbuf_d_601(.A(n3706), .Y(d_out_601));
CLKBUFX1 gbuf_q_601(.A(q_in_601), .Y(H1[22]));
CLKBUFX1 gbuf_d_602(.A(n3705), .Y(d_out_602));
CLKBUFX1 gbuf_q_602(.A(q_in_602), .Y(H1[23]));
CLKBUFX1 gbuf_d_603(.A(n3928), .Y(d_out_603));
CLKBUFX1 gbuf_q_603(.A(q_in_603), .Y(next_C[22]));
CLKBUFX1 gbuf_qn_603(.A(qn_in_603), .Y(n13010));
CLKBUFX1 gbuf_d_604(.A(n3704), .Y(d_out_604));
CLKBUFX1 gbuf_q_604(.A(q_in_604), .Y(H1[24]));
CLKBUFX1 gbuf_d_605(.A(n3927), .Y(d_out_605));
CLKBUFX1 gbuf_q_605(.A(q_in_605), .Y(next_C[23]));
CLKBUFX1 gbuf_qn_605(.A(qn_in_605), .Y(n13009));
CLKBUFX1 gbuf_d_606(.A(n3703), .Y(d_out_606));
CLKBUFX1 gbuf_q_606(.A(q_in_606), .Y(H1[25]));
CLKBUFX1 gbuf_d_607(.A(n3926), .Y(d_out_607));
CLKBUFX1 gbuf_q_607(.A(q_in_607), .Y(next_C[24]));
CLKBUFX1 gbuf_qn_607(.A(qn_in_607), .Y(n13003));
CLKBUFX1 gbuf_d_608(.A(n3702), .Y(d_out_608));
CLKBUFX1 gbuf_q_608(.A(q_in_608), .Y(H1[26]));
CLKBUFX1 gbuf_d_609(.A(n3925), .Y(d_out_609));
CLKBUFX1 gbuf_q_609(.A(q_in_609), .Y(next_C[25]));
CLKBUFX1 gbuf_qn_609(.A(qn_in_609), .Y(n13008));
CLKBUFX1 gbuf_d_610(.A(n3701), .Y(d_out_610));
CLKBUFX1 gbuf_q_610(.A(q_in_610), .Y(H1[27]));
CLKBUFX1 gbuf_d_611(.A(n3924), .Y(d_out_611));
CLKBUFX1 gbuf_q_611(.A(q_in_611), .Y(next_C[26]));
CLKBUFX1 gbuf_qn_611(.A(qn_in_611), .Y(n13014));
CLKBUFX1 gbuf_d_612(.A(n3700), .Y(d_out_612));
CLKBUFX1 gbuf_q_612(.A(q_in_612), .Y(H1[28]));
CLKBUFX1 gbuf_d_613(.A(n3923), .Y(d_out_613));
CLKBUFX1 gbuf_q_613(.A(q_in_613), .Y(next_C[27]));
CLKBUFX1 gbuf_qn_613(.A(qn_in_613), .Y(n13013));
CLKBUFX1 gbuf_d_614(.A(n3699), .Y(d_out_614));
CLKBUFX1 gbuf_q_614(.A(q_in_614), .Y(H1[29]));
CLKBUFX1 gbuf_d_615(.A(n3921), .Y(d_out_615));
CLKBUFX1 gbuf_q_615(.A(q_in_615), .Y(next_C[29]));
CLKBUFX1 gbuf_qn_615(.A(qn_in_615), .Y(n13002));
CLKBUFX1 gbuf_d_616(.A(n3697), .Y(d_out_616));
CLKBUFX1 gbuf_q_616(.A(q_in_616), .Y(H1[31]));
CLKBUFX1 gbuf_d_617(.A(n3892), .Y(d_out_617));
CLKBUFX1 gbuf_q_617(.A(q_in_617), .Y(SHA1_result[92]));
CLKBUFX1 gbuf_qn_617(.A(qn_in_617), .Y(n447));
CLKBUFX1 gbuf_d_618(.A(n3732), .Y(d_out_618));
CLKBUFX1 gbuf_q_618(.A(q_in_618), .Y(H2[28]));
CLKBUFX1 gbuf_d_619(.A(n3920), .Y(d_out_619));
CLKBUFX1 gbuf_q_619(.A(q_in_619), .Y(SHA1_result[64]));
CLKBUFX1 gbuf_qn_619(.A(qn_in_619), .Y(n475));
CLKBUFX1 gbuf_d_620(.A(n3760), .Y(d_out_620));
CLKBUFX1 gbuf_q_620(.A(q_in_620), .Y(H2[0]));
CLKBUFX1 gbuf_d_621(.A(n3918), .Y(d_out_621));
CLKBUFX1 gbuf_q_621(.A(q_in_621), .Y(SHA1_result[66]));
CLKBUFX1 gbuf_qn_621(.A(qn_in_621), .Y(n473));
CLKBUFX1 gbuf_d_622(.A(n3917), .Y(d_out_622));
CLKBUFX1 gbuf_q_622(.A(q_in_622), .Y(SHA1_result[67]));
CLKBUFX1 gbuf_qn_622(.A(qn_in_622), .Y(n472));
CLKBUFX1 gbuf_d_623(.A(n3916), .Y(d_out_623));
CLKBUFX1 gbuf_q_623(.A(q_in_623), .Y(SHA1_result[68]));
CLKBUFX1 gbuf_qn_623(.A(qn_in_623), .Y(n471));
CLKBUFX1 gbuf_d_624(.A(n3915), .Y(d_out_624));
CLKBUFX1 gbuf_q_624(.A(q_in_624), .Y(SHA1_result[69]));
CLKBUFX1 gbuf_qn_624(.A(qn_in_624), .Y(n470));
CLKBUFX1 gbuf_d_625(.A(n3914), .Y(d_out_625));
CLKBUFX1 gbuf_q_625(.A(q_in_625), .Y(SHA1_result[70]));
CLKBUFX1 gbuf_d_626(.A(n3913), .Y(d_out_626));
CLKBUFX1 gbuf_q_626(.A(q_in_626), .Y(SHA1_result[71]));
CLKBUFX1 gbuf_qn_626(.A(qn_in_626), .Y(n468));
CLKBUFX1 gbuf_d_627(.A(n3912), .Y(d_out_627));
CLKBUFX1 gbuf_q_627(.A(q_in_627), .Y(SHA1_result[72]));
CLKBUFX1 gbuf_qn_627(.A(qn_in_627), .Y(n467));
CLKBUFX1 gbuf_d_628(.A(n3752), .Y(d_out_628));
CLKBUFX1 gbuf_q_628(.A(q_in_628), .Y(H2[8]));
CLKBUFX1 gbuf_d_629(.A(n3911), .Y(d_out_629));
CLKBUFX1 gbuf_q_629(.A(q_in_629), .Y(SHA1_result[73]));
CLKBUFX1 gbuf_qn_629(.A(qn_in_629), .Y(n466));
CLKBUFX1 gbuf_d_630(.A(n3751), .Y(d_out_630));
CLKBUFX1 gbuf_q_630(.A(q_in_630), .Y(H2[9]));
CLKBUFX1 gbuf_d_631(.A(n3910), .Y(d_out_631));
CLKBUFX1 gbuf_q_631(.A(q_in_631), .Y(SHA1_result[74]));
CLKBUFX1 gbuf_qn_631(.A(qn_in_631), .Y(n465));
CLKBUFX1 gbuf_d_632(.A(n3909), .Y(d_out_632));
CLKBUFX1 gbuf_q_632(.A(q_in_632), .Y(SHA1_result[75]));
CLKBUFX1 gbuf_qn_632(.A(qn_in_632), .Y(n464));
CLKBUFX1 gbuf_d_633(.A(n3908), .Y(d_out_633));
CLKBUFX1 gbuf_q_633(.A(q_in_633), .Y(SHA1_result[76]));
CLKBUFX1 gbuf_qn_633(.A(qn_in_633), .Y(n463));
CLKBUFX1 gbuf_d_634(.A(n3748), .Y(d_out_634));
CLKBUFX1 gbuf_q_634(.A(q_in_634), .Y(H2[12]));
CLKBUFX1 gbuf_d_635(.A(n3907), .Y(d_out_635));
CLKBUFX1 gbuf_q_635(.A(q_in_635), .Y(SHA1_result[77]));
CLKBUFX1 gbuf_qn_635(.A(qn_in_635), .Y(n462));
CLKBUFX1 gbuf_d_636(.A(n3747), .Y(d_out_636));
CLKBUFX1 gbuf_q_636(.A(q_in_636), .Y(H2[13]));
CLKBUFX1 gbuf_d_637(.A(n3906), .Y(d_out_637));
CLKBUFX1 gbuf_q_637(.A(q_in_637), .Y(SHA1_result[78]));
CLKBUFX1 gbuf_qn_637(.A(qn_in_637), .Y(n461));
CLKBUFX1 gbuf_d_638(.A(n3746), .Y(d_out_638));
CLKBUFX1 gbuf_q_638(.A(q_in_638), .Y(H2[14]));
CLKBUFX1 gbuf_d_639(.A(n3905), .Y(d_out_639));
CLKBUFX1 gbuf_q_639(.A(q_in_639), .Y(SHA1_result[79]));
CLKBUFX1 gbuf_qn_639(.A(qn_in_639), .Y(n460));
CLKBUFX1 gbuf_d_640(.A(n3745), .Y(d_out_640));
CLKBUFX1 gbuf_q_640(.A(q_in_640), .Y(H2[15]));
CLKBUFX1 gbuf_d_641(.A(n3904), .Y(d_out_641));
CLKBUFX1 gbuf_q_641(.A(q_in_641), .Y(SHA1_result[80]));
CLKBUFX1 gbuf_qn_641(.A(qn_in_641), .Y(n459));
CLKBUFX1 gbuf_d_642(.A(n3744), .Y(d_out_642));
CLKBUFX1 gbuf_q_642(.A(q_in_642), .Y(H2[16]));
CLKBUFX1 gbuf_d_643(.A(n3903), .Y(d_out_643));
CLKBUFX1 gbuf_q_643(.A(q_in_643), .Y(SHA1_result[81]));
CLKBUFX1 gbuf_qn_643(.A(qn_in_643), .Y(n458));
CLKBUFX1 gbuf_d_644(.A(n3743), .Y(d_out_644));
CLKBUFX1 gbuf_q_644(.A(q_in_644), .Y(H2[17]));
CLKBUFX1 gbuf_d_645(.A(n3902), .Y(d_out_645));
CLKBUFX1 gbuf_q_645(.A(q_in_645), .Y(SHA1_result[82]));
CLKBUFX1 gbuf_qn_645(.A(qn_in_645), .Y(n457));
CLKBUFX1 gbuf_d_646(.A(n3742), .Y(d_out_646));
CLKBUFX1 gbuf_q_646(.A(q_in_646), .Y(H2[18]));
CLKBUFX1 gbuf_d_647(.A(n3901), .Y(d_out_647));
CLKBUFX1 gbuf_q_647(.A(q_in_647), .Y(SHA1_result[83]));
CLKBUFX1 gbuf_qn_647(.A(qn_in_647), .Y(n456));
CLKBUFX1 gbuf_d_648(.A(n3741), .Y(d_out_648));
CLKBUFX1 gbuf_q_648(.A(q_in_648), .Y(H2[19]));
CLKBUFX1 gbuf_d_649(.A(n3900), .Y(d_out_649));
CLKBUFX1 gbuf_q_649(.A(q_in_649), .Y(SHA1_result[84]));
CLKBUFX1 gbuf_qn_649(.A(qn_in_649), .Y(n455));
CLKBUFX1 gbuf_d_650(.A(n3740), .Y(d_out_650));
CLKBUFX1 gbuf_q_650(.A(q_in_650), .Y(H2[20]));
CLKBUFX1 gbuf_d_651(.A(n3899), .Y(d_out_651));
CLKBUFX1 gbuf_q_651(.A(q_in_651), .Y(SHA1_result[85]));
CLKBUFX1 gbuf_qn_651(.A(qn_in_651), .Y(n454));
CLKBUFX1 gbuf_d_652(.A(n3739), .Y(d_out_652));
CLKBUFX1 gbuf_q_652(.A(q_in_652), .Y(H2[21]));
CLKBUFX1 gbuf_d_653(.A(n3898), .Y(d_out_653));
CLKBUFX1 gbuf_q_653(.A(q_in_653), .Y(SHA1_result[86]));
CLKBUFX1 gbuf_qn_653(.A(qn_in_653), .Y(n453));
CLKBUFX1 gbuf_d_654(.A(n3738), .Y(d_out_654));
CLKBUFX1 gbuf_q_654(.A(q_in_654), .Y(H2[22]));
CLKBUFX1 gbuf_d_655(.A(n3897), .Y(d_out_655));
CLKBUFX1 gbuf_q_655(.A(q_in_655), .Y(SHA1_result[87]));
CLKBUFX1 gbuf_qn_655(.A(qn_in_655), .Y(n452));
CLKBUFX1 gbuf_d_656(.A(n3737), .Y(d_out_656));
CLKBUFX1 gbuf_q_656(.A(q_in_656), .Y(H2[23]));
CLKBUFX1 gbuf_d_657(.A(n3896), .Y(d_out_657));
CLKBUFX1 gbuf_q_657(.A(q_in_657), .Y(SHA1_result[88]));
CLKBUFX1 gbuf_qn_657(.A(qn_in_657), .Y(n451));
CLKBUFX1 gbuf_d_658(.A(n3736), .Y(d_out_658));
CLKBUFX1 gbuf_q_658(.A(q_in_658), .Y(H2[24]));
CLKBUFX1 gbuf_d_659(.A(n3895), .Y(d_out_659));
CLKBUFX1 gbuf_q_659(.A(q_in_659), .Y(SHA1_result[89]));
CLKBUFX1 gbuf_qn_659(.A(qn_in_659), .Y(n450));
CLKBUFX1 gbuf_d_660(.A(n3735), .Y(d_out_660));
CLKBUFX1 gbuf_q_660(.A(q_in_660), .Y(H2[25]));
CLKBUFX1 gbuf_d_661(.A(n3894), .Y(d_out_661));
CLKBUFX1 gbuf_q_661(.A(q_in_661), .Y(SHA1_result[90]));
CLKBUFX1 gbuf_qn_661(.A(qn_in_661), .Y(n449));
CLKBUFX1 gbuf_d_662(.A(n3734), .Y(d_out_662));
CLKBUFX1 gbuf_q_662(.A(q_in_662), .Y(H2[26]));
CLKBUFX1 gbuf_d_663(.A(n3893), .Y(d_out_663));
CLKBUFX1 gbuf_q_663(.A(q_in_663), .Y(SHA1_result[91]));
CLKBUFX1 gbuf_qn_663(.A(qn_in_663), .Y(n448));
CLKBUFX1 gbuf_d_664(.A(n3733), .Y(d_out_664));
CLKBUFX1 gbuf_q_664(.A(q_in_664), .Y(H2[27]));
CLKBUFX1 gbuf_d_665(.A(n3891), .Y(d_out_665));
CLKBUFX1 gbuf_q_665(.A(q_in_665), .Y(SHA1_result[93]));
CLKBUFX1 gbuf_qn_665(.A(qn_in_665), .Y(n446));
CLKBUFX1 gbuf_d_666(.A(n3731), .Y(d_out_666));
CLKBUFX1 gbuf_q_666(.A(q_in_666), .Y(H2[29]));
CLKBUFX1 gbuf_d_667(.A(n3890), .Y(d_out_667));
CLKBUFX1 gbuf_q_667(.A(q_in_667), .Y(SHA1_result[94]));
CLKBUFX1 gbuf_qn_667(.A(qn_in_667), .Y(n445));
CLKBUFX1 gbuf_d_668(.A(n3730), .Y(d_out_668));
CLKBUFX1 gbuf_q_668(.A(q_in_668), .Y(H2[30]));
CLKBUFX1 gbuf_d_669(.A(n3889), .Y(d_out_669));
CLKBUFX1 gbuf_q_669(.A(q_in_669), .Y(SHA1_result[95]));
CLKBUFX1 gbuf_qn_669(.A(qn_in_669), .Y(n444));
CLKBUFX1 gbuf_d_670(.A(n3729), .Y(d_out_670));
CLKBUFX1 gbuf_q_670(.A(q_in_670), .Y(H2[31]));
CLKBUFX1 gbuf_d_671(.A(n3860), .Y(d_out_671));
CLKBUFX1 gbuf_q_671(.A(q_in_671), .Y(SHA1_result[60]));
CLKBUFX1 gbuf_d_672(.A(n3888), .Y(d_out_672));
CLKBUFX1 gbuf_q_672(.A(q_in_672), .Y(SHA1_result[32]));
CLKBUFX1 gbuf_qn_672(.A(qn_in_672), .Y(n443));
CLKBUFX1 gbuf_d_673(.A(n3887), .Y(d_out_673));
CLKBUFX1 gbuf_q_673(.A(q_in_673), .Y(SHA1_result[33]));
CLKBUFX1 gbuf_qn_673(.A(qn_in_673), .Y(n442));
CLKBUFX1 gbuf_d_674(.A(n3855), .Y(d_out_674));
CLKBUFX1 gbuf_q_674(.A(q_in_674), .Y(H3[1]));
CLKBUFX1 gbuf_d_675(.A(n3886), .Y(d_out_675));
CLKBUFX1 gbuf_q_675(.A(q_in_675), .Y(SHA1_result[34]));
CLKBUFX1 gbuf_d_676(.A(n3885), .Y(d_out_676));
CLKBUFX1 gbuf_q_676(.A(q_in_676), .Y(SHA1_result[35]));
CLKBUFX1 gbuf_qn_676(.A(qn_in_676), .Y(n440));
CLKBUFX1 gbuf_d_677(.A(n3884), .Y(d_out_677));
CLKBUFX1 gbuf_q_677(.A(q_in_677), .Y(SHA1_result[36]));
CLKBUFX1 gbuf_d_678(.A(n3883), .Y(d_out_678));
CLKBUFX1 gbuf_q_678(.A(q_in_678), .Y(SHA1_result[37]));
CLKBUFX1 gbuf_qn_678(.A(qn_in_678), .Y(n438));
CLKBUFX1 gbuf_d_679(.A(n3882), .Y(d_out_679));
CLKBUFX1 gbuf_q_679(.A(q_in_679), .Y(SHA1_result[38]));
CLKBUFX1 gbuf_qn_679(.A(qn_in_679), .Y(n437));
CLKBUFX1 gbuf_d_680(.A(n3881), .Y(d_out_680));
CLKBUFX1 gbuf_q_680(.A(q_in_680), .Y(SHA1_result[39]));
CLKBUFX1 gbuf_d_681(.A(n3880), .Y(d_out_681));
CLKBUFX1 gbuf_q_681(.A(q_in_681), .Y(SHA1_result[40]));
CLKBUFX1 gbuf_d_682(.A(n3848), .Y(d_out_682));
CLKBUFX1 gbuf_q_682(.A(q_in_682), .Y(H3[8]));
CLKBUFX1 gbuf_d_683(.A(n3847), .Y(d_out_683));
CLKBUFX1 gbuf_q_683(.A(q_in_683), .Y(H3[9]));
CLKBUFX1 gbuf_d_684(.A(n3878), .Y(d_out_684));
CLKBUFX1 gbuf_q_684(.A(q_in_684), .Y(SHA1_result[42]));
CLKBUFX1 gbuf_qn_684(.A(qn_in_684), .Y(n433));
CLKBUFX1 gbuf_d_685(.A(n3877), .Y(d_out_685));
CLKBUFX1 gbuf_q_685(.A(q_in_685), .Y(n14810));
CLKBUFX1 gbuf_d_686(.A(n3845), .Y(d_out_686));
CLKBUFX1 gbuf_q_686(.A(q_in_686), .Y(H3[11]));
CLKBUFX1 gbuf_d_687(.A(n3876), .Y(d_out_687));
CLKBUFX1 gbuf_q_687(.A(q_in_687), .Y(n14817));
CLKBUFX1 gbuf_d_688(.A(n3875), .Y(d_out_688));
CLKBUFX1 gbuf_q_688(.A(q_in_688), .Y(SHA1_result[45]));
CLKBUFX1 gbuf_d_689(.A(n3843), .Y(d_out_689));
CLKBUFX1 gbuf_q_689(.A(q_in_689), .Y(H3[13]));
CLKBUFX1 gbuf_d_690(.A(n3874), .Y(d_out_690));
CLKBUFX1 gbuf_q_690(.A(q_in_690), .Y(n14830));
CLKBUFX1 gbuf_d_691(.A(n3873), .Y(d_out_691));
CLKBUFX1 gbuf_q_691(.A(q_in_691), .Y(SHA1_result[47]));
CLKBUFX1 gbuf_d_692(.A(n3841), .Y(d_out_692));
CLKBUFX1 gbuf_q_692(.A(q_in_692), .Y(H3[15]));
CLKBUFX1 gbuf_d_693(.A(n3872), .Y(d_out_693));
CLKBUFX1 gbuf_q_693(.A(q_in_693), .Y(SHA1_result[48]));
CLKBUFX1 gbuf_d_694(.A(n3840), .Y(d_out_694));
CLKBUFX1 gbuf_q_694(.A(q_in_694), .Y(H3[16]));
CLKBUFX1 gbuf_d_695(.A(n3871), .Y(d_out_695));
CLKBUFX1 gbuf_q_695(.A(q_in_695), .Y(SHA1_result[49]));
CLKBUFX1 gbuf_d_696(.A(n3870), .Y(d_out_696));
CLKBUFX1 gbuf_q_696(.A(q_in_696), .Y(SHA1_result[50]));
CLKBUFX1 gbuf_d_697(.A(n3838), .Y(d_out_697));
CLKBUFX1 gbuf_q_697(.A(q_in_697), .Y(H3[18]));
CLKBUFX1 gbuf_d_698(.A(n3869), .Y(d_out_698));
CLKBUFX1 gbuf_q_698(.A(q_in_698), .Y(SHA1_result[51]));
CLKBUFX1 gbuf_d_699(.A(n3837), .Y(d_out_699));
CLKBUFX1 gbuf_q_699(.A(q_in_699), .Y(H3[19]));
CLKBUFX1 gbuf_d_700(.A(n3868), .Y(d_out_700));
CLKBUFX1 gbuf_q_700(.A(q_in_700), .Y(SHA1_result[52]));
CLKBUFX1 gbuf_qn_700(.A(qn_in_700), .Y(n423));
CLKBUFX1 gbuf_d_701(.A(n3867), .Y(d_out_701));
CLKBUFX1 gbuf_q_701(.A(q_in_701), .Y(SHA1_result[53]));
CLKBUFX1 gbuf_qn_701(.A(qn_in_701), .Y(n422));
CLKBUFX1 gbuf_d_702(.A(n3866), .Y(d_out_702));
CLKBUFX1 gbuf_q_702(.A(q_in_702), .Y(n14681));
CLKBUFX1 gbuf_d_703(.A(n3834), .Y(d_out_703));
CLKBUFX1 gbuf_q_703(.A(q_in_703), .Y(H3[22]));
CLKBUFX1 gbuf_d_704(.A(n3865), .Y(d_out_704));
CLKBUFX1 gbuf_q_704(.A(q_in_704), .Y(SHA1_result[55]));
CLKBUFX1 gbuf_d_705(.A(n3833), .Y(d_out_705));
CLKBUFX1 gbuf_q_705(.A(q_in_705), .Y(H3[23]));
CLKBUFX1 gbuf_d_706(.A(n3864), .Y(d_out_706));
CLKBUFX1 gbuf_q_706(.A(q_in_706), .Y(SHA1_result[56]));
CLKBUFX1 gbuf_d_707(.A(n3832), .Y(d_out_707));
CLKBUFX1 gbuf_q_707(.A(q_in_707), .Y(H3[24]));
CLKBUFX1 gbuf_d_708(.A(n3863), .Y(d_out_708));
CLKBUFX1 gbuf_q_708(.A(q_in_708), .Y(SHA1_result[57]));
CLKBUFX1 gbuf_d_709(.A(n3831), .Y(d_out_709));
CLKBUFX1 gbuf_q_709(.A(q_in_709), .Y(H3[25]));
CLKBUFX1 gbuf_d_710(.A(n3862), .Y(d_out_710));
CLKBUFX1 gbuf_q_710(.A(q_in_710), .Y(SHA1_result[58]));
CLKBUFX1 gbuf_d_711(.A(n3830), .Y(d_out_711));
CLKBUFX1 gbuf_q_711(.A(q_in_711), .Y(H3[26]));
CLKBUFX1 gbuf_d_712(.A(n3861), .Y(d_out_712));
CLKBUFX1 gbuf_q_712(.A(q_in_712), .Y(SHA1_result[59]));
CLKBUFX1 gbuf_d_713(.A(n3829), .Y(d_out_713));
CLKBUFX1 gbuf_q_713(.A(q_in_713), .Y(H3[27]));
CLKBUFX1 gbuf_d_714(.A(n3859), .Y(d_out_714));
CLKBUFX1 gbuf_q_714(.A(q_in_714), .Y(SHA1_result[61]));
CLKBUFX1 gbuf_d_715(.A(n3827), .Y(d_out_715));
CLKBUFX1 gbuf_q_715(.A(q_in_715), .Y(H3[29]));
CLKBUFX1 gbuf_d_716(.A(n3858), .Y(d_out_716));
CLKBUFX1 gbuf_q_716(.A(q_in_716), .Y(SHA1_result[62]));
CLKBUFX1 gbuf_d_717(.A(n3826), .Y(d_out_717));
CLKBUFX1 gbuf_q_717(.A(q_in_717), .Y(H3[30]));
CLKBUFX1 gbuf_d_718(.A(n3857), .Y(d_out_718));
CLKBUFX1 gbuf_q_718(.A(q_in_718), .Y(SHA1_result[63]));
CLKBUFX1 gbuf_qn_718(.A(qn_in_718), .Y(n412));
CLKBUFX1 gbuf_d_719(.A(n3793), .Y(d_out_719));
CLKBUFX1 gbuf_q_719(.A(q_in_719), .Y(SHA1_result[31]));
CLKBUFX1 gbuf_d_720(.A(n3824), .Y(d_out_720));
CLKBUFX1 gbuf_q_720(.A(q_in_720), .Y(SHA1_result[0]));
CLKBUFX1 gbuf_d_721(.A(n3792), .Y(d_out_721));
CLKBUFX1 gbuf_q_721(.A(q_in_721), .Y(H4[0]));
CLKBUFX1 gbuf_d_722(.A(n3823), .Y(d_out_722));
CLKBUFX1 gbuf_q_722(.A(q_in_722), .Y(SHA1_result[1]));
CLKBUFX1 gbuf_d_723(.A(n3791), .Y(d_out_723));
CLKBUFX1 gbuf_q_723(.A(q_in_723), .Y(H4[1]));
CLKBUFX1 gbuf_d_724(.A(n3822), .Y(d_out_724));
CLKBUFX1 gbuf_q_724(.A(q_in_724), .Y(SHA1_result[2]));
CLKBUFX1 gbuf_d_725(.A(n3790), .Y(d_out_725));
CLKBUFX1 gbuf_q_725(.A(q_in_725), .Y(H4[2]));
CLKBUFX1 gbuf_d_726(.A(n3821), .Y(d_out_726));
CLKBUFX1 gbuf_q_726(.A(q_in_726), .Y(SHA1_result[3]));
CLKBUFX1 gbuf_d_727(.A(n3789), .Y(d_out_727));
CLKBUFX1 gbuf_q_727(.A(q_in_727), .Y(H4[3]));
CLKBUFX1 gbuf_d_728(.A(n3820), .Y(d_out_728));
CLKBUFX1 gbuf_q_728(.A(q_in_728), .Y(SHA1_result[4]));
CLKBUFX1 gbuf_d_729(.A(n3788), .Y(d_out_729));
CLKBUFX1 gbuf_q_729(.A(q_in_729), .Y(H4[4]));
CLKBUFX1 gbuf_d_730(.A(n3819), .Y(d_out_730));
CLKBUFX1 gbuf_q_730(.A(q_in_730), .Y(SHA1_result[5]));
CLKBUFX1 gbuf_d_731(.A(n3787), .Y(d_out_731));
CLKBUFX1 gbuf_q_731(.A(q_in_731), .Y(H4[5]));
CLKBUFX1 gbuf_d_732(.A(n3818), .Y(d_out_732));
CLKBUFX1 gbuf_q_732(.A(q_in_732), .Y(SHA1_result[6]));
CLKBUFX1 gbuf_d_733(.A(n3786), .Y(d_out_733));
CLKBUFX1 gbuf_q_733(.A(q_in_733), .Y(H4[6]));
CLKBUFX1 gbuf_d_734(.A(n3817), .Y(d_out_734));
CLKBUFX1 gbuf_q_734(.A(q_in_734), .Y(SHA1_result[7]));
CLKBUFX1 gbuf_d_735(.A(n3785), .Y(d_out_735));
CLKBUFX1 gbuf_q_735(.A(q_in_735), .Y(H4[7]));
CLKBUFX1 gbuf_d_736(.A(n3816), .Y(d_out_736));
CLKBUFX1 gbuf_q_736(.A(q_in_736), .Y(SHA1_result[8]));
CLKBUFX1 gbuf_d_737(.A(n3784), .Y(d_out_737));
CLKBUFX1 gbuf_q_737(.A(q_in_737), .Y(H4[8]));
CLKBUFX1 gbuf_d_738(.A(n3815), .Y(d_out_738));
CLKBUFX1 gbuf_q_738(.A(q_in_738), .Y(SHA1_result[9]));
CLKBUFX1 gbuf_d_739(.A(n3783), .Y(d_out_739));
CLKBUFX1 gbuf_q_739(.A(q_in_739), .Y(H4[9]));
CLKBUFX1 gbuf_d_740(.A(n3814), .Y(d_out_740));
CLKBUFX1 gbuf_q_740(.A(q_in_740), .Y(SHA1_result[10]));
CLKBUFX1 gbuf_d_741(.A(n3782), .Y(d_out_741));
CLKBUFX1 gbuf_q_741(.A(q_in_741), .Y(H4[10]));
CLKBUFX1 gbuf_d_742(.A(n3813), .Y(d_out_742));
CLKBUFX1 gbuf_q_742(.A(q_in_742), .Y(SHA1_result[11]));
CLKBUFX1 gbuf_d_743(.A(n3781), .Y(d_out_743));
CLKBUFX1 gbuf_q_743(.A(q_in_743), .Y(H4[11]));
CLKBUFX1 gbuf_d_744(.A(n3812), .Y(d_out_744));
CLKBUFX1 gbuf_q_744(.A(q_in_744), .Y(SHA1_result[12]));
CLKBUFX1 gbuf_d_745(.A(n3780), .Y(d_out_745));
CLKBUFX1 gbuf_q_745(.A(q_in_745), .Y(H4[12]));
CLKBUFX1 gbuf_d_746(.A(n3811), .Y(d_out_746));
CLKBUFX1 gbuf_q_746(.A(q_in_746), .Y(SHA1_result[13]));
CLKBUFX1 gbuf_d_747(.A(n3779), .Y(d_out_747));
CLKBUFX1 gbuf_q_747(.A(q_in_747), .Y(H4[13]));
CLKBUFX1 gbuf_d_748(.A(n3810), .Y(d_out_748));
CLKBUFX1 gbuf_q_748(.A(q_in_748), .Y(SHA1_result[14]));
CLKBUFX1 gbuf_d_749(.A(n3778), .Y(d_out_749));
CLKBUFX1 gbuf_q_749(.A(q_in_749), .Y(H4[14]));
CLKBUFX1 gbuf_d_750(.A(n3809), .Y(d_out_750));
CLKBUFX1 gbuf_q_750(.A(q_in_750), .Y(SHA1_result[15]));
CLKBUFX1 gbuf_d_751(.A(n3777), .Y(d_out_751));
CLKBUFX1 gbuf_q_751(.A(q_in_751), .Y(H4[15]));
CLKBUFX1 gbuf_d_752(.A(n3808), .Y(d_out_752));
CLKBUFX1 gbuf_q_752(.A(q_in_752), .Y(SHA1_result[16]));
CLKBUFX1 gbuf_d_753(.A(n3776), .Y(d_out_753));
CLKBUFX1 gbuf_q_753(.A(q_in_753), .Y(H4[16]));
CLKBUFX1 gbuf_d_754(.A(n3807), .Y(d_out_754));
CLKBUFX1 gbuf_q_754(.A(q_in_754), .Y(SHA1_result[17]));
CLKBUFX1 gbuf_d_755(.A(n3775), .Y(d_out_755));
CLKBUFX1 gbuf_q_755(.A(q_in_755), .Y(H4[17]));
CLKBUFX1 gbuf_d_756(.A(n3806), .Y(d_out_756));
CLKBUFX1 gbuf_q_756(.A(q_in_756), .Y(SHA1_result[18]));
CLKBUFX1 gbuf_d_757(.A(n3774), .Y(d_out_757));
CLKBUFX1 gbuf_q_757(.A(q_in_757), .Y(H4[18]));
CLKBUFX1 gbuf_d_758(.A(n3805), .Y(d_out_758));
CLKBUFX1 gbuf_q_758(.A(q_in_758), .Y(SHA1_result[19]));
CLKBUFX1 gbuf_d_759(.A(n3773), .Y(d_out_759));
CLKBUFX1 gbuf_q_759(.A(q_in_759), .Y(H4[19]));
CLKBUFX1 gbuf_d_760(.A(n3804), .Y(d_out_760));
CLKBUFX1 gbuf_q_760(.A(q_in_760), .Y(SHA1_result[20]));
CLKBUFX1 gbuf_d_761(.A(n3772), .Y(d_out_761));
CLKBUFX1 gbuf_q_761(.A(q_in_761), .Y(H4[20]));
CLKBUFX1 gbuf_d_762(.A(n3803), .Y(d_out_762));
CLKBUFX1 gbuf_q_762(.A(q_in_762), .Y(SHA1_result[21]));
CLKBUFX1 gbuf_d_763(.A(n3771), .Y(d_out_763));
CLKBUFX1 gbuf_q_763(.A(q_in_763), .Y(H4[21]));
CLKBUFX1 gbuf_d_764(.A(n3802), .Y(d_out_764));
CLKBUFX1 gbuf_q_764(.A(q_in_764), .Y(SHA1_result[22]));
CLKBUFX1 gbuf_d_765(.A(n3770), .Y(d_out_765));
CLKBUFX1 gbuf_q_765(.A(q_in_765), .Y(H4[22]));
CLKBUFX1 gbuf_d_766(.A(n3801), .Y(d_out_766));
CLKBUFX1 gbuf_q_766(.A(q_in_766), .Y(SHA1_result[23]));
CLKBUFX1 gbuf_d_767(.A(n3800), .Y(d_out_767));
CLKBUFX1 gbuf_q_767(.A(q_in_767), .Y(SHA1_result[24]));
CLKBUFX1 gbuf_d_768(.A(n3799), .Y(d_out_768));
CLKBUFX1 gbuf_q_768(.A(q_in_768), .Y(SHA1_result[25]));
CLKBUFX1 gbuf_d_769(.A(n3798), .Y(d_out_769));
CLKBUFX1 gbuf_q_769(.A(q_in_769), .Y(SHA1_result[26]));
CLKBUFX1 gbuf_d_770(.A(n3766), .Y(d_out_770));
CLKBUFX1 gbuf_q_770(.A(q_in_770), .Y(H4[26]));
CLKBUFX1 gbuf_d_771(.A(n3797), .Y(d_out_771));
CLKBUFX1 gbuf_q_771(.A(q_in_771), .Y(SHA1_result[27]));
CLKBUFX1 gbuf_d_772(.A(n3765), .Y(d_out_772));
CLKBUFX1 gbuf_q_772(.A(q_in_772), .Y(H4[27]));
CLKBUFX1 gbuf_d_773(.A(n3796), .Y(d_out_773));
CLKBUFX1 gbuf_q_773(.A(q_in_773), .Y(SHA1_result[28]));
CLKBUFX1 gbuf_d_774(.A(n3764), .Y(d_out_774));
CLKBUFX1 gbuf_q_774(.A(q_in_774), .Y(H4[28]));
CLKBUFX1 gbuf_d_775(.A(n3795), .Y(d_out_775));
CLKBUFX1 gbuf_q_775(.A(q_in_775), .Y(SHA1_result[29]));
CLKBUFX1 gbuf_d_776(.A(n3763), .Y(d_out_776));
CLKBUFX1 gbuf_q_776(.A(q_in_776), .Y(H4[29]));
CLKBUFX1 gbuf_d_777(.A(n3794), .Y(d_out_777));
CLKBUFX1 gbuf_q_777(.A(q_in_777), .Y(SHA1_result[30]));
CLKBUFX1 gbuf_d_778(.A(n3825), .Y(d_out_778));
CLKBUFX1 gbuf_q_778(.A(q_in_778), .Y(H3[31]));
CLKBUFX1 gbuf_d_779(.A(n3954), .Y(d_out_779));
CLKBUFX1 gbuf_q_779(.A(q_in_779), .Y(H0[30]));
CLKBUFX1 gbuf_d_780(.A(n3662), .Y(d_out_780));
CLKBUFX1 gbuf_q_780(.A(q_in_780), .Y(text_o[31]));
CLKBUFX1 gbuf_qn_780(.A(qn_in_780), .Y(n12914));
CLKBUFX1 gbuf_d_781(.A(n3663), .Y(d_out_781));
CLKBUFX1 gbuf_q_781(.A(q_in_781), .Y(text_o[30]));
CLKBUFX1 gbuf_qn_781(.A(qn_in_781), .Y(n12912));
CLKBUFX1 gbuf_d_782(.A(n3664), .Y(d_out_782));
CLKBUFX1 gbuf_q_782(.A(q_in_782), .Y(text_o[29]));
CLKBUFX1 gbuf_qn_782(.A(qn_in_782), .Y(n12910));
CLKBUFX1 gbuf_d_783(.A(n3665), .Y(d_out_783));
CLKBUFX1 gbuf_q_783(.A(q_in_783), .Y(text_o[28]));
CLKBUFX1 gbuf_qn_783(.A(qn_in_783), .Y(n12908));
CLKBUFX1 gbuf_d_784(.A(n3666), .Y(d_out_784));
CLKBUFX1 gbuf_q_784(.A(q_in_784), .Y(text_o[27]));
CLKBUFX1 gbuf_qn_784(.A(qn_in_784), .Y(n12906));
CLKBUFX1 gbuf_d_785(.A(n3667), .Y(d_out_785));
CLKBUFX1 gbuf_q_785(.A(q_in_785), .Y(text_o[26]));
CLKBUFX1 gbuf_qn_785(.A(qn_in_785), .Y(n12904));
CLKBUFX1 gbuf_d_786(.A(n3668), .Y(d_out_786));
CLKBUFX1 gbuf_q_786(.A(q_in_786), .Y(text_o[25]));
CLKBUFX1 gbuf_qn_786(.A(qn_in_786), .Y(n12902));
CLKBUFX1 gbuf_d_787(.A(n3669), .Y(d_out_787));
CLKBUFX1 gbuf_q_787(.A(q_in_787), .Y(text_o[24]));
CLKBUFX1 gbuf_qn_787(.A(qn_in_787), .Y(n12900));
CLKBUFX1 gbuf_d_788(.A(n3670), .Y(d_out_788));
CLKBUFX1 gbuf_q_788(.A(q_in_788), .Y(text_o[23]));
CLKBUFX1 gbuf_qn_788(.A(qn_in_788), .Y(n12898));
CLKBUFX1 gbuf_d_789(.A(n3671), .Y(d_out_789));
CLKBUFX1 gbuf_q_789(.A(q_in_789), .Y(text_o[22]));
CLKBUFX1 gbuf_qn_789(.A(qn_in_789), .Y(n12896));
CLKBUFX1 gbuf_d_790(.A(n3672), .Y(d_out_790));
CLKBUFX1 gbuf_q_790(.A(q_in_790), .Y(text_o[21]));
CLKBUFX1 gbuf_qn_790(.A(qn_in_790), .Y(n12894));
CLKBUFX1 gbuf_d_791(.A(n3673), .Y(d_out_791));
CLKBUFX1 gbuf_q_791(.A(q_in_791), .Y(text_o[20]));
CLKBUFX1 gbuf_qn_791(.A(qn_in_791), .Y(n12892));
CLKBUFX1 gbuf_d_792(.A(n3674), .Y(d_out_792));
CLKBUFX1 gbuf_q_792(.A(q_in_792), .Y(text_o[19]));
CLKBUFX1 gbuf_qn_792(.A(qn_in_792), .Y(n12890));
CLKBUFX1 gbuf_d_793(.A(n3675), .Y(d_out_793));
CLKBUFX1 gbuf_q_793(.A(q_in_793), .Y(text_o[18]));
CLKBUFX1 gbuf_qn_793(.A(qn_in_793), .Y(n12888));
CLKBUFX1 gbuf_d_794(.A(n3676), .Y(d_out_794));
CLKBUFX1 gbuf_q_794(.A(q_in_794), .Y(text_o[17]));
CLKBUFX1 gbuf_qn_794(.A(qn_in_794), .Y(n12886));
CLKBUFX1 gbuf_d_795(.A(n3677), .Y(d_out_795));
CLKBUFX1 gbuf_q_795(.A(q_in_795), .Y(text_o[16]));
CLKBUFX1 gbuf_qn_795(.A(qn_in_795), .Y(n12884));
CLKBUFX1 gbuf_d_796(.A(n3678), .Y(d_out_796));
CLKBUFX1 gbuf_q_796(.A(q_in_796), .Y(text_o[15]));
CLKBUFX1 gbuf_qn_796(.A(qn_in_796), .Y(n12882));
CLKBUFX1 gbuf_d_797(.A(n3679), .Y(d_out_797));
CLKBUFX1 gbuf_q_797(.A(q_in_797), .Y(text_o[14]));
CLKBUFX1 gbuf_qn_797(.A(qn_in_797), .Y(n12880));
CLKBUFX1 gbuf_d_798(.A(n3680), .Y(d_out_798));
CLKBUFX1 gbuf_q_798(.A(q_in_798), .Y(text_o[13]));
CLKBUFX1 gbuf_qn_798(.A(qn_in_798), .Y(n12878));
CLKBUFX1 gbuf_d_799(.A(n3681), .Y(d_out_799));
CLKBUFX1 gbuf_q_799(.A(q_in_799), .Y(text_o[12]));
CLKBUFX1 gbuf_qn_799(.A(qn_in_799), .Y(n12876));
CLKBUFX1 gbuf_d_800(.A(n3682), .Y(d_out_800));
CLKBUFX1 gbuf_q_800(.A(q_in_800), .Y(text_o[11]));
CLKBUFX1 gbuf_qn_800(.A(qn_in_800), .Y(n12874));
CLKBUFX1 gbuf_d_801(.A(n3683), .Y(d_out_801));
CLKBUFX1 gbuf_q_801(.A(q_in_801), .Y(text_o[10]));
CLKBUFX1 gbuf_qn_801(.A(qn_in_801), .Y(n12872));
CLKBUFX1 gbuf_d_802(.A(n3684), .Y(d_out_802));
CLKBUFX1 gbuf_q_802(.A(q_in_802), .Y(text_o[9]));
CLKBUFX1 gbuf_qn_802(.A(qn_in_802), .Y(n12870));
CLKBUFX1 gbuf_d_803(.A(n3685), .Y(d_out_803));
CLKBUFX1 gbuf_q_803(.A(q_in_803), .Y(text_o[8]));
CLKBUFX1 gbuf_qn_803(.A(qn_in_803), .Y(n12868));
CLKBUFX1 gbuf_d_804(.A(n3686), .Y(d_out_804));
CLKBUFX1 gbuf_q_804(.A(q_in_804), .Y(text_o[7]));
CLKBUFX1 gbuf_qn_804(.A(qn_in_804), .Y(n12866));
CLKBUFX1 gbuf_d_805(.A(n3687), .Y(d_out_805));
CLKBUFX1 gbuf_q_805(.A(q_in_805), .Y(text_o[6]));
CLKBUFX1 gbuf_qn_805(.A(qn_in_805), .Y(n12864));
CLKBUFX1 gbuf_d_806(.A(n3688), .Y(d_out_806));
CLKBUFX1 gbuf_q_806(.A(q_in_806), .Y(text_o[5]));
CLKBUFX1 gbuf_qn_806(.A(qn_in_806), .Y(n12862));
CLKBUFX1 gbuf_d_807(.A(n3689), .Y(d_out_807));
CLKBUFX1 gbuf_q_807(.A(q_in_807), .Y(text_o[4]));
CLKBUFX1 gbuf_qn_807(.A(qn_in_807), .Y(n12860));
CLKBUFX1 gbuf_d_808(.A(n3690), .Y(d_out_808));
CLKBUFX1 gbuf_q_808(.A(q_in_808), .Y(text_o[3]));
CLKBUFX1 gbuf_qn_808(.A(qn_in_808), .Y(n12858));
CLKBUFX1 gbuf_d_809(.A(n3691), .Y(d_out_809));
CLKBUFX1 gbuf_q_809(.A(q_in_809), .Y(text_o[2]));
CLKBUFX1 gbuf_qn_809(.A(qn_in_809), .Y(n12856));
CLKBUFX1 gbuf_d_810(.A(n3692), .Y(d_out_810));
CLKBUFX1 gbuf_q_810(.A(q_in_810), .Y(text_o[1]));
CLKBUFX1 gbuf_qn_810(.A(qn_in_810), .Y(n12854));
CLKBUFX1 gbuf_d_811(.A(n3693), .Y(d_out_811));
CLKBUFX1 gbuf_q_811(.A(q_in_811), .Y(text_o[0]));
CLKBUFX1 gbuf_qn_811(.A(qn_in_811), .Y(n12852));
NAND2_X2 U4142 ( .A1(n9302), .A2(n9303), .ZN(n4532) );
NAND2_X2 U4144 ( .A1(n14933), .A2(n9304), .ZN(n9302) );
OR3_X2 U4149 ( .A1(cmd_w_i), .A2(n8326), .A3(n13395), .ZN(n9311) );
NAND2_X2 U4152 ( .A1(n9309), .A2(cmd_o[1]), .ZN(n9314) );
NAND2_X2 U4157 ( .A1(n13315), .A2(n15424), .ZN(n9317) );
XOR2_X2 U4163 ( .A(n9326), .B(n9327), .Z(n9325) );
XNOR2_X2 U4164 ( .A(n15411), .B(n8323), .ZN(n9327) );
XNOR2_X2 U4165 ( .A(n15419), .B(n12978), .ZN(n9326) );
XOR2_X2 U4170 ( .A(n9333), .B(n9334), .Z(n9332) );
XNOR2_X2 U4171 ( .A(n14963), .B(n8322), .ZN(n9334) );
XNOR2_X2 U4172 ( .A(n14971), .B(n12976), .ZN(n9333) );
XOR2_X2 U4177 ( .A(n9339), .B(n9340), .Z(n9338) );
XNOR2_X2 U4178 ( .A(n14977), .B(n8320), .ZN(n9340) );
XNOR2_X2 U4179 ( .A(n14985), .B(n12974), .ZN(n9339) );
XOR2_X2 U4184 ( .A(n9345), .B(n9346), .Z(n9344) );
XNOR2_X2 U4185 ( .A(n14991), .B(n8318), .ZN(n9346) );
XNOR2_X2 U4186 ( .A(n14999), .B(n12972), .ZN(n9345) );
XOR2_X2 U4191 ( .A(n9351), .B(n9352), .Z(n9350) );
XNOR2_X2 U4192 ( .A(n15005), .B(n8316), .ZN(n9352) );
XNOR2_X2 U4193 ( .A(n15013), .B(n12970), .ZN(n9351) );
XOR2_X2 U4198 ( .A(n9357), .B(n9358), .Z(n9356) );
XNOR2_X2 U4199 ( .A(n15019), .B(n8314), .ZN(n9358) );
XNOR2_X2 U4200 ( .A(n15027), .B(n12968), .ZN(n9357) );
XOR2_X2 U4205 ( .A(n9363), .B(n9364), .Z(n9362) );
XNOR2_X2 U4206 ( .A(n15033), .B(n8312), .ZN(n9364) );
XNOR2_X2 U4207 ( .A(n15041), .B(n12966), .ZN(n9363) );
XOR2_X2 U4212 ( .A(n9369), .B(n9370), .Z(n9368) );
XNOR2_X2 U4213 ( .A(n15047), .B(n8310), .ZN(n9370) );
XNOR2_X2 U4214 ( .A(n15055), .B(n12964), .ZN(n9369) );
XOR2_X2 U4219 ( .A(n9375), .B(n9376), .Z(n9374) );
XNOR2_X2 U4220 ( .A(n15061), .B(n8308), .ZN(n9376) );
XNOR2_X2 U4221 ( .A(n15069), .B(n12962), .ZN(n9375) );
XOR2_X2 U4226 ( .A(n9381), .B(n9382), .Z(n9380) );
XNOR2_X2 U4227 ( .A(n15075), .B(n8306), .ZN(n9382) );
XNOR2_X2 U4228 ( .A(n15083), .B(n12960), .ZN(n9381) );
XOR2_X2 U4233 ( .A(n9387), .B(n9388), .Z(n9386) );
XNOR2_X2 U4234 ( .A(n15089), .B(n8304), .ZN(n9388) );
XNOR2_X2 U4235 ( .A(n15097), .B(n12958), .ZN(n9387) );
XOR2_X2 U4240 ( .A(n9393), .B(n9394), .Z(n9392) );
XNOR2_X2 U4241 ( .A(n15103), .B(n8302), .ZN(n9394) );
XNOR2_X2 U4242 ( .A(n15111), .B(n12956), .ZN(n9393) );
XOR2_X2 U4247 ( .A(n9399), .B(n9400), .Z(n9398) );
XNOR2_X2 U4248 ( .A(n15117), .B(n8300), .ZN(n9400) );
XNOR2_X2 U4249 ( .A(n15125), .B(n12954), .ZN(n9399) );
XOR2_X2 U4254 ( .A(n9405), .B(n9406), .Z(n9404) );
XNOR2_X2 U4255 ( .A(n15131), .B(n8298), .ZN(n9406) );
XNOR2_X2 U4256 ( .A(n15139), .B(n12952), .ZN(n9405) );
XOR2_X2 U4261 ( .A(n9411), .B(n9412), .Z(n9410) );
XNOR2_X2 U4262 ( .A(n15145), .B(n8296), .ZN(n9412) );
XNOR2_X2 U4263 ( .A(n15153), .B(n12950), .ZN(n9411) );
XOR2_X2 U4268 ( .A(n9417), .B(n9418), .Z(n9416) );
XNOR2_X2 U4269 ( .A(n15159), .B(n8294), .ZN(n9418) );
XNOR2_X2 U4270 ( .A(n15167), .B(n12948), .ZN(n9417) );
XOR2_X2 U4275 ( .A(n9423), .B(n9424), .Z(n9422) );
XNOR2_X2 U4276 ( .A(n15173), .B(n8292), .ZN(n9424) );
XNOR2_X2 U4277 ( .A(n15181), .B(n12946), .ZN(n9423) );
XOR2_X2 U4282 ( .A(n9429), .B(n9430), .Z(n9428) );
XNOR2_X2 U4283 ( .A(n15187), .B(n8290), .ZN(n9430) );
XNOR2_X2 U4284 ( .A(n15195), .B(n12944), .ZN(n9429) );
NAND2_X2 U4288 ( .A1(n13315), .A2(n9434), .ZN(n9432) );
XOR2_X2 U4289 ( .A(n9435), .B(n9436), .Z(n9434) );
XNOR2_X2 U4290 ( .A(n15201), .B(n8288), .ZN(n9436) );
XNOR2_X2 U4291 ( .A(n15209), .B(n12942), .ZN(n9435) );
NAND2_X2 U4295 ( .A1(n13315), .A2(n9440), .ZN(n9438) );
XOR2_X2 U4296 ( .A(n9441), .B(n9442), .Z(n9440) );
XNOR2_X2 U4297 ( .A(n15216), .B(n8286), .ZN(n9442) );
XNOR2_X2 U4298 ( .A(n15224), .B(n12940), .ZN(n9441) );
NAND2_X2 U4302 ( .A1(n13314), .A2(n9446), .ZN(n9444) );
XOR2_X2 U4303 ( .A(n9447), .B(n9448), .Z(n9446) );
XNOR2_X2 U4304 ( .A(n15231), .B(n8284), .ZN(n9448) );
XNOR2_X2 U4305 ( .A(n15239), .B(n12938), .ZN(n9447) );
NAND2_X2 U4309 ( .A1(n13314), .A2(n9452), .ZN(n9450) );
XOR2_X2 U4310 ( .A(n9453), .B(n9454), .Z(n9452) );
XNOR2_X2 U4311 ( .A(n15246), .B(n8282), .ZN(n9454) );
XNOR2_X2 U4312 ( .A(n15254), .B(n12936), .ZN(n9453) );
NAND2_X2 U4316 ( .A1(n13314), .A2(n9458), .ZN(n9456) );
XOR2_X2 U4317 ( .A(n9459), .B(n9460), .Z(n9458) );
XNOR2_X2 U4318 ( .A(n15261), .B(n8280), .ZN(n9460) );
XNOR2_X2 U4319 ( .A(n15269), .B(n12934), .ZN(n9459) );
NAND2_X2 U4323 ( .A1(n13314), .A2(n9464), .ZN(n9462) );
XOR2_X2 U4324 ( .A(n9465), .B(n9466), .Z(n9464) );
XNOR2_X2 U4325 ( .A(n15276), .B(n8278), .ZN(n9466) );
XNOR2_X2 U4326 ( .A(n15284), .B(n12932), .ZN(n9465) );
NAND2_X2 U4330 ( .A1(n13314), .A2(n9470), .ZN(n9468) );
XOR2_X2 U4331 ( .A(n9471), .B(n9472), .Z(n9470) );
XNOR2_X2 U4332 ( .A(n15291), .B(n8276), .ZN(n9472) );
XNOR2_X2 U4333 ( .A(n15299), .B(n12930), .ZN(n9471) );
NAND2_X2 U4337 ( .A1(n13314), .A2(n9476), .ZN(n9474) );
XOR2_X2 U4338 ( .A(n9477), .B(n9478), .Z(n9476) );
XNOR2_X2 U4339 ( .A(n15306), .B(n8274), .ZN(n9478) );
XNOR2_X2 U4340 ( .A(n15314), .B(n12928), .ZN(n9477) );
NAND2_X2 U4344 ( .A1(n13314), .A2(n9482), .ZN(n9480) );
XOR2_X2 U4345 ( .A(n9483), .B(n9484), .Z(n9482) );
XNOR2_X2 U4346 ( .A(n15321), .B(n8272), .ZN(n9484) );
XNOR2_X2 U4347 ( .A(n15329), .B(n12926), .ZN(n9483) );
NAND2_X2 U4351 ( .A1(n13314), .A2(n9488), .ZN(n9486) );
XOR2_X2 U4352 ( .A(n9489), .B(n9490), .Z(n9488) );
XNOR2_X2 U4353 ( .A(n15336), .B(n8270), .ZN(n9490) );
XNOR2_X2 U4354 ( .A(n15344), .B(n12924), .ZN(n9489) );
NAND2_X2 U4358 ( .A1(n13314), .A2(n9494), .ZN(n9492) );
XOR2_X2 U4359 ( .A(n9495), .B(n9496), .Z(n9494) );
XNOR2_X2 U4360 ( .A(n15351), .B(n8268), .ZN(n9496) );
XNOR2_X2 U4361 ( .A(n15359), .B(n12922), .ZN(n9495) );
NAND2_X2 U4365 ( .A1(n13314), .A2(n9500), .ZN(n9498) );
XOR2_X2 U4366 ( .A(n9501), .B(n9502), .Z(n9500) );
XNOR2_X2 U4367 ( .A(n15366), .B(n8266), .ZN(n9502) );
XNOR2_X2 U4368 ( .A(n15374), .B(n12920), .ZN(n9501) );
NAND2_X2 U4372 ( .A1(n13314), .A2(n9506), .ZN(n9504) );
XOR2_X2 U4373 ( .A(n9507), .B(n9508), .Z(n9506) );
XNOR2_X2 U4374 ( .A(n15381), .B(n8264), .ZN(n9508) );
XNOR2_X2 U4375 ( .A(n15389), .B(n12918), .ZN(n9507) );
NAND2_X2 U4379 ( .A1(n13313), .A2(n9512), .ZN(n9510) );
XOR2_X2 U4380 ( .A(n9513), .B(n9514), .Z(n9512) );
XNOR2_X2 U4381 ( .A(n15396), .B(n8262), .ZN(n9514) );
XNOR2_X2 U4382 ( .A(n15404), .B(n12916), .ZN(n9513) );
NAND2_X2 U4460 ( .A1(n13313), .A2(Wt[18]), .ZN(n9577) );
NAND2_X2 U4462 ( .A1(n13268), .A2(n13045), .ZN(n9575) );
NAND2_X2 U4464 ( .A1(n13313), .A2(Wt[19]), .ZN(n9580) );
NAND2_X2 U4466 ( .A1(n13268), .A2(n13044), .ZN(n9578) );
NAND2_X2 U4468 ( .A1(n13313), .A2(Wt[20]), .ZN(n9583) );
NAND2_X2 U4470 ( .A1(n13268), .A2(n13043), .ZN(n9581) );
NAND2_X2 U4472 ( .A1(n13313), .A2(Wt[21]), .ZN(n9586) );
NAND2_X2 U4474 ( .A1(n13267), .A2(n13042), .ZN(n9584) );
NAND2_X2 U4476 ( .A1(n13313), .A2(Wt[22]), .ZN(n9589) );
NAND2_X2 U4478 ( .A1(n13267), .A2(n13041), .ZN(n9587) );
NAND2_X2 U4480 ( .A1(n13313), .A2(Wt[23]), .ZN(n9592) );
NAND2_X2 U4482 ( .A1(n13267), .A2(n13040), .ZN(n9590) );
NAND2_X2 U4484 ( .A1(n13313), .A2(Wt[24]), .ZN(n9595) );
NAND2_X2 U4486 ( .A1(n13267), .A2(n13039), .ZN(n9593) );
NAND2_X2 U4488 ( .A1(n13313), .A2(Wt[25]), .ZN(n9598) );
NAND2_X2 U4490 ( .A1(n13267), .A2(n13038), .ZN(n9596) );
NAND2_X2 U4492 ( .A1(n13313), .A2(Wt[26]), .ZN(n9601) );
NAND2_X2 U4494 ( .A1(n13267), .A2(n13037), .ZN(n9599) );
NAND2_X2 U4496 ( .A1(n13313), .A2(Wt[27]), .ZN(n9604) );
NAND2_X2 U4498 ( .A1(n13267), .A2(n13036), .ZN(n9602) );
NAND2_X2 U4500 ( .A1(n13312), .A2(Wt[28]), .ZN(n9607) );
NAND2_X2 U4502 ( .A1(n13267), .A2(n13035), .ZN(n9605) );
NAND2_X2 U4504 ( .A1(n13312), .A2(Wt[29]), .ZN(n9610) );
NAND2_X2 U4506 ( .A1(n13267), .A2(n13034), .ZN(n9608) );
NAND2_X2 U4508 ( .A1(n13312), .A2(Wt[30]), .ZN(n9613) );
NAND2_X2 U4510 ( .A1(n13267), .A2(n13033), .ZN(n9611) );
NAND2_X2 U4512 ( .A1(n13312), .A2(Wt[31]), .ZN(n9616) );
NAND2_X2 U4515 ( .A1(n13267), .A2(n13032), .ZN(n9614) );
NAND2_X2 U4519 ( .A1(n13312), .A2(n14951), .ZN(n9623) );
NAND2_X2 U4521 ( .A1(n13391), .A2(n13063), .ZN(n9621) );
NAND2_X2 U4523 ( .A1(n13312), .A2(n14934), .ZN(n9628) );
NAND2_X2 U4525 ( .A1(n13391), .A2(n13062), .ZN(n9626) );
NAND2_X2 U4527 ( .A1(n13312), .A2(n14935), .ZN(n9631) );
NAND2_X2 U4529 ( .A1(n13391), .A2(n13061), .ZN(n9629) );
NAND2_X2 U4531 ( .A1(n13312), .A2(n14936), .ZN(n9634) );
NAND2_X2 U4533 ( .A1(n13391), .A2(n13060), .ZN(n9632) );
NAND2_X2 U4535 ( .A1(n13312), .A2(n14937), .ZN(n9637) );
NAND2_X2 U4537 ( .A1(n13391), .A2(n13059), .ZN(n9635) );
NAND2_X2 U4539 ( .A1(n13312), .A2(n14938), .ZN(n9640) );
NAND2_X2 U4541 ( .A1(n13391), .A2(n13058), .ZN(n9638) );
NAND2_X2 U4543 ( .A1(n13312), .A2(n14939), .ZN(n9643) );
NAND2_X2 U4545 ( .A1(n13391), .A2(n13057), .ZN(n9641) );
NAND2_X2 U4547 ( .A1(n13311), .A2(n14940), .ZN(n9646) );
NAND2_X2 U4549 ( .A1(n13391), .A2(n13056), .ZN(n9644) );
NAND2_X2 U4551 ( .A1(n13311), .A2(n14941), .ZN(n9649) );
NAND2_X2 U4553 ( .A1(n13391), .A2(n13055), .ZN(n9647) );
NAND2_X2 U4555 ( .A1(n13311), .A2(n14942), .ZN(n9652) );
NAND2_X2 U4557 ( .A1(n13391), .A2(n13054), .ZN(n9650) );
NAND2_X2 U4559 ( .A1(n13311), .A2(n14943), .ZN(n9655) );
NAND2_X2 U4561 ( .A1(n13390), .A2(n13053), .ZN(n9653) );
NAND2_X2 U4563 ( .A1(n13311), .A2(n14944), .ZN(n9658) );
NAND2_X2 U4565 ( .A1(n13390), .A2(n13052), .ZN(n9656) );
NAND2_X2 U4567 ( .A1(n13311), .A2(n14945), .ZN(n9661) );
NAND2_X2 U4569 ( .A1(n13390), .A2(n13051), .ZN(n9659) );
NAND2_X2 U4571 ( .A1(n13311), .A2(n14946), .ZN(n9664) );
NAND2_X2 U4573 ( .A1(n13390), .A2(n13050), .ZN(n9662) );
NAND2_X2 U4575 ( .A1(n13311), .A2(n14947), .ZN(n9667) );
NAND2_X2 U4577 ( .A1(n13390), .A2(n13049), .ZN(n9665) );
NAND2_X2 U4579 ( .A1(n13311), .A2(n14948), .ZN(n9670) );
NAND2_X2 U4581 ( .A1(n13390), .A2(n13048), .ZN(n9668) );
NAND2_X2 U4583 ( .A1(n13311), .A2(n14949), .ZN(n9673) );
NAND2_X2 U4585 ( .A1(n13390), .A2(n13047), .ZN(n9671) );
NAND2_X2 U4587 ( .A1(n13311), .A2(n14950), .ZN(n9676) );
NAND2_X2 U4589 ( .A1(n13390), .A2(n13046), .ZN(n9674) );
NAND2_X2 U4591 ( .A1(n13310), .A2(n15210), .ZN(n9679) );
NAND2_X2 U4593 ( .A1(n13390), .A2(n13045), .ZN(n9677) );
NAND2_X2 U4595 ( .A1(n13310), .A2(n15225), .ZN(n9682) );
NAND2_X2 U4597 ( .A1(n13390), .A2(n13044), .ZN(n9680) );
NAND2_X2 U4599 ( .A1(n13310), .A2(n15240), .ZN(n9685) );
NAND2_X2 U4601 ( .A1(n13390), .A2(n13043), .ZN(n9683) );
NAND2_X2 U4603 ( .A1(n13310), .A2(n15255), .ZN(n9688) );
NAND2_X2 U4605 ( .A1(n13389), .A2(n13042), .ZN(n9686) );
NAND2_X2 U4607 ( .A1(n13310), .A2(n15270), .ZN(n9691) );
NAND2_X2 U4609 ( .A1(n13389), .A2(n13041), .ZN(n9689) );
NAND2_X2 U4611 ( .A1(n13310), .A2(n15285), .ZN(n9694) );
NAND2_X2 U4613 ( .A1(n13389), .A2(n13040), .ZN(n9692) );
NAND2_X2 U4615 ( .A1(n13310), .A2(n15300), .ZN(n9697) );
NAND2_X2 U4617 ( .A1(n13389), .A2(n13039), .ZN(n9695) );
NAND2_X2 U4619 ( .A1(n13310), .A2(n15315), .ZN(n9700) );
NAND2_X2 U4621 ( .A1(n13389), .A2(n13038), .ZN(n9698) );
NAND2_X2 U4623 ( .A1(n13310), .A2(n15330), .ZN(n9703) );
NAND2_X2 U4625 ( .A1(n13389), .A2(n13037), .ZN(n9701) );
NAND2_X2 U4627 ( .A1(n13310), .A2(n15345), .ZN(n9706) );
NAND2_X2 U4629 ( .A1(n13389), .A2(n13036), .ZN(n9704) );
NAND2_X2 U4631 ( .A1(n13310), .A2(n15360), .ZN(n9709) );
NAND2_X2 U4633 ( .A1(n13389), .A2(n13035), .ZN(n9707) );
NAND2_X2 U4635 ( .A1(n13309), .A2(n15375), .ZN(n9712) );
NAND2_X2 U4637 ( .A1(n13389), .A2(n13034), .ZN(n9710) );
NAND2_X2 U4639 ( .A1(n13309), .A2(n15390), .ZN(n9715) );
NAND2_X2 U4641 ( .A1(n13389), .A2(n13033), .ZN(n9713) );
NAND2_X2 U4643 ( .A1(n13309), .A2(n15405), .ZN(n9718) );
NAND2_X2 U4646 ( .A1(n13389), .A2(n13032), .ZN(n9716) );
NAND2_X2 U4650 ( .A1(n13309), .A2(n15420), .ZN(n9723) );
NAND2_X2 U4652 ( .A1(n13388), .A2(n13063), .ZN(n9721) );
NAND2_X2 U4654 ( .A1(n13309), .A2(n14972), .ZN(n9728) );
NAND2_X2 U4656 ( .A1(n13388), .A2(n13062), .ZN(n9726) );
NAND2_X2 U4658 ( .A1(n13309), .A2(n14986), .ZN(n9731) );
NAND2_X2 U4660 ( .A1(n13388), .A2(n13061), .ZN(n9729) );
NAND2_X2 U4662 ( .A1(n13309), .A2(n15000), .ZN(n9734) );
NAND2_X2 U4664 ( .A1(n13388), .A2(n13060), .ZN(n9732) );
NAND2_X2 U4666 ( .A1(n13309), .A2(n15014), .ZN(n9737) );
NAND2_X2 U4668 ( .A1(n13388), .A2(n13059), .ZN(n9735) );
NAND2_X2 U4670 ( .A1(n13309), .A2(n15028), .ZN(n9740) );
NAND2_X2 U4672 ( .A1(n13388), .A2(n13058), .ZN(n9738) );
NAND2_X2 U4674 ( .A1(n13309), .A2(n15042), .ZN(n9743) );
NAND2_X2 U4676 ( .A1(n13388), .A2(n13057), .ZN(n9741) );
NAND2_X2 U4678 ( .A1(n13309), .A2(n15056), .ZN(n9746) );
NAND2_X2 U4680 ( .A1(n13388), .A2(n13056), .ZN(n9744) );
NAND2_X2 U4682 ( .A1(n13308), .A2(n15070), .ZN(n9749) );
NAND2_X2 U4684 ( .A1(n13388), .A2(n13055), .ZN(n9747) );
NAND2_X2 U4686 ( .A1(n13308), .A2(n15084), .ZN(n9752) );
NAND2_X2 U4688 ( .A1(n13388), .A2(n13054), .ZN(n9750) );
NAND2_X2 U4690 ( .A1(n13308), .A2(n15098), .ZN(n9755) );
NAND2_X2 U4692 ( .A1(n13387), .A2(n13053), .ZN(n9753) );
NAND2_X2 U4694 ( .A1(n13308), .A2(n15112), .ZN(n9758) );
NAND2_X2 U4696 ( .A1(n13387), .A2(n13052), .ZN(n9756) );
NAND2_X2 U4698 ( .A1(n13308), .A2(n15126), .ZN(n9761) );
NAND2_X2 U4700 ( .A1(n13387), .A2(n13051), .ZN(n9759) );
NAND2_X2 U4702 ( .A1(n13308), .A2(n15140), .ZN(n9764) );
NAND2_X2 U4704 ( .A1(n13387), .A2(n13050), .ZN(n9762) );
NAND2_X2 U4706 ( .A1(n13308), .A2(n15154), .ZN(n9767) );
NAND2_X2 U4708 ( .A1(n13387), .A2(n13049), .ZN(n9765) );
NAND2_X2 U4710 ( .A1(n13308), .A2(n15168), .ZN(n9770) );
NAND2_X2 U4712 ( .A1(n13387), .A2(n13048), .ZN(n9768) );
NAND2_X2 U4714 ( .A1(n13308), .A2(n15182), .ZN(n9773) );
NAND2_X2 U4716 ( .A1(n13387), .A2(n13047), .ZN(n9771) );
NAND2_X2 U4718 ( .A1(n13308), .A2(n15196), .ZN(n9776) );
NAND2_X2 U4720 ( .A1(n13387), .A2(n13046), .ZN(n9774) );
NAND2_X2 U4722 ( .A1(n13308), .A2(n15211), .ZN(n9779) );
NAND2_X2 U4724 ( .A1(n13387), .A2(n13045), .ZN(n9777) );
NAND2_X2 U4726 ( .A1(n13307), .A2(n15226), .ZN(n9782) );
NAND2_X2 U4728 ( .A1(n13387), .A2(n13044), .ZN(n9780) );
NAND2_X2 U4730 ( .A1(n13307), .A2(n15241), .ZN(n9785) );
NAND2_X2 U4732 ( .A1(n13387), .A2(n13043), .ZN(n9783) );
NAND2_X2 U4734 ( .A1(n13307), .A2(n15256), .ZN(n9788) );
NAND2_X2 U4736 ( .A1(n13386), .A2(n13042), .ZN(n9786) );
NAND2_X2 U4738 ( .A1(n13307), .A2(n15271), .ZN(n9791) );
NAND2_X2 U4740 ( .A1(n13386), .A2(n13041), .ZN(n9789) );
NAND2_X2 U4742 ( .A1(n13307), .A2(n15286), .ZN(n9794) );
NAND2_X2 U4744 ( .A1(n13386), .A2(n13040), .ZN(n9792) );
NAND2_X2 U4746 ( .A1(n13307), .A2(n15301), .ZN(n9797) );
NAND2_X2 U4748 ( .A1(n13386), .A2(n13039), .ZN(n9795) );
NAND2_X2 U4750 ( .A1(n13307), .A2(n15316), .ZN(n9800) );
NAND2_X2 U4752 ( .A1(n13386), .A2(n13038), .ZN(n9798) );
NAND2_X2 U4754 ( .A1(n13307), .A2(n15331), .ZN(n9803) );
NAND2_X2 U4756 ( .A1(n13386), .A2(n13037), .ZN(n9801) );
NAND2_X2 U4758 ( .A1(n13307), .A2(n15346), .ZN(n9806) );
NAND2_X2 U4760 ( .A1(n13386), .A2(n13036), .ZN(n9804) );
NAND2_X2 U4762 ( .A1(n13307), .A2(n15361), .ZN(n9809) );
NAND2_X2 U4764 ( .A1(n13386), .A2(n13035), .ZN(n9807) );
NAND2_X2 U4766 ( .A1(n13307), .A2(n15376), .ZN(n9812) );
NAND2_X2 U4768 ( .A1(n13386), .A2(n13034), .ZN(n9810) );
NAND2_X2 U4770 ( .A1(n13306), .A2(n15391), .ZN(n9815) );
NAND2_X2 U4772 ( .A1(n13386), .A2(n13033), .ZN(n9813) );
NAND2_X2 U4774 ( .A1(n13306), .A2(n15406), .ZN(n9818) );
NAND2_X2 U4777 ( .A1(n13386), .A2(n13032), .ZN(n9816) );
NAND2_X2 U4780 ( .A1(n13306), .A2(n15421), .ZN(n9822) );
NAND2_X2 U4782 ( .A1(n13385), .A2(n13063), .ZN(n9820) );
NAND2_X2 U4784 ( .A1(n13306), .A2(n14973), .ZN(n9827) );
NAND2_X2 U4786 ( .A1(n13385), .A2(n13062), .ZN(n9825) );
NAND2_X2 U4788 ( .A1(n13306), .A2(n14987), .ZN(n9830) );
NAND2_X2 U4790 ( .A1(n13385), .A2(n13061), .ZN(n9828) );
NAND2_X2 U4792 ( .A1(n13306), .A2(n15001), .ZN(n9833) );
NAND2_X2 U4794 ( .A1(n13385), .A2(n13060), .ZN(n9831) );
NAND2_X2 U4796 ( .A1(n13306), .A2(n15015), .ZN(n9836) );
NAND2_X2 U4798 ( .A1(n13385), .A2(n13059), .ZN(n9834) );
NAND2_X2 U4800 ( .A1(n13306), .A2(n15029), .ZN(n9839) );
NAND2_X2 U4802 ( .A1(n13385), .A2(n13058), .ZN(n9837) );
NAND2_X2 U4804 ( .A1(n13306), .A2(n15043), .ZN(n9842) );
NAND2_X2 U4806 ( .A1(n13385), .A2(n13057), .ZN(n9840) );
NAND2_X2 U4808 ( .A1(n13306), .A2(n15057), .ZN(n9845) );
NAND2_X2 U4810 ( .A1(n13385), .A2(n13056), .ZN(n9843) );
NAND2_X2 U4812 ( .A1(n13306), .A2(n15071), .ZN(n9848) );
NAND2_X2 U4814 ( .A1(n13385), .A2(n13055), .ZN(n9846) );
NAND2_X2 U4816 ( .A1(n13305), .A2(n15085), .ZN(n9851) );
NAND2_X2 U4818 ( .A1(n13385), .A2(n13054), .ZN(n9849) );
NAND2_X2 U4820 ( .A1(n13305), .A2(n15099), .ZN(n9854) );
NAND2_X2 U4822 ( .A1(n13384), .A2(n13053), .ZN(n9852) );
NAND2_X2 U4824 ( .A1(n13305), .A2(n15113), .ZN(n9857) );
NAND2_X2 U4826 ( .A1(n13384), .A2(n13052), .ZN(n9855) );
NAND2_X2 U4828 ( .A1(n13305), .A2(n15127), .ZN(n9860) );
NAND2_X2 U4830 ( .A1(n13384), .A2(n13051), .ZN(n9858) );
NAND2_X2 U4832 ( .A1(n13305), .A2(n15141), .ZN(n9863) );
NAND2_X2 U4834 ( .A1(n13384), .A2(n13050), .ZN(n9861) );
NAND2_X2 U4836 ( .A1(n13305), .A2(n15155), .ZN(n9866) );
NAND2_X2 U4838 ( .A1(n13384), .A2(n13049), .ZN(n9864) );
NAND2_X2 U4840 ( .A1(n13305), .A2(n15169), .ZN(n9869) );
NAND2_X2 U4842 ( .A1(n13384), .A2(n13048), .ZN(n9867) );
NAND2_X2 U4844 ( .A1(n13305), .A2(n15183), .ZN(n9872) );
NAND2_X2 U4846 ( .A1(n13384), .A2(n13047), .ZN(n9870) );
NAND2_X2 U4848 ( .A1(n13305), .A2(n15197), .ZN(n9875) );
NAND2_X2 U4850 ( .A1(n13384), .A2(n13046), .ZN(n9873) );
NAND2_X2 U4852 ( .A1(n13305), .A2(n15212), .ZN(n9878) );
NAND2_X2 U4854 ( .A1(n13384), .A2(n13045), .ZN(n9876) );
NAND2_X2 U4856 ( .A1(n13305), .A2(n15227), .ZN(n9881) );
NAND2_X2 U4858 ( .A1(n13384), .A2(n13044), .ZN(n9879) );
NAND2_X2 U4860 ( .A1(n13304), .A2(n15242), .ZN(n9884) );
NAND2_X2 U4862 ( .A1(n13384), .A2(n13043), .ZN(n9882) );
NAND2_X2 U4864 ( .A1(n13304), .A2(n15257), .ZN(n9887) );
NAND2_X2 U4866 ( .A1(n13383), .A2(n13042), .ZN(n9885) );
NAND2_X2 U4868 ( .A1(n13304), .A2(n15272), .ZN(n9890) );
NAND2_X2 U4870 ( .A1(n13383), .A2(n13041), .ZN(n9888) );
NAND2_X2 U4872 ( .A1(n13304), .A2(n15287), .ZN(n9893) );
NAND2_X2 U4874 ( .A1(n13383), .A2(n13040), .ZN(n9891) );
NAND2_X2 U4876 ( .A1(n13304), .A2(n15302), .ZN(n9896) );
NAND2_X2 U4878 ( .A1(n13383), .A2(n13039), .ZN(n9894) );
NAND2_X2 U4880 ( .A1(n13304), .A2(n15317), .ZN(n9899) );
NAND2_X2 U4882 ( .A1(n13383), .A2(n13038), .ZN(n9897) );
NAND2_X2 U4884 ( .A1(n13304), .A2(n15332), .ZN(n9902) );
NAND2_X2 U4886 ( .A1(n13383), .A2(n13037), .ZN(n9900) );
NAND2_X2 U4888 ( .A1(n13304), .A2(n15347), .ZN(n9905) );
NAND2_X2 U4890 ( .A1(n13383), .A2(n13036), .ZN(n9903) );
NAND2_X2 U4892 ( .A1(n13304), .A2(n15362), .ZN(n9908) );
NAND2_X2 U4894 ( .A1(n13383), .A2(n13035), .ZN(n9906) );
NAND2_X2 U4896 ( .A1(n13304), .A2(n15377), .ZN(n9911) );
NAND2_X2 U4898 ( .A1(n13383), .A2(n13034), .ZN(n9909) );
NAND2_X2 U4900 ( .A1(n13304), .A2(n15392), .ZN(n9914) );
NAND2_X2 U4902 ( .A1(n13383), .A2(n13033), .ZN(n9912) );
NAND2_X2 U4904 ( .A1(n13303), .A2(n15407), .ZN(n9917) );
NAND2_X2 U4908 ( .A1(n13383), .A2(n13032), .ZN(n9915) );
NAND2_X2 U4911 ( .A1(n13303), .A2(n15422), .ZN(n9923) );
NAND2_X2 U4913 ( .A1(n13380), .A2(n13063), .ZN(n9921) );
NAND2_X2 U4915 ( .A1(n13303), .A2(n14974), .ZN(n9928) );
NAND2_X2 U4917 ( .A1(n13380), .A2(n13062), .ZN(n9926) );
NAND2_X2 U4919 ( .A1(n13303), .A2(n14988), .ZN(n9931) );
NAND2_X2 U4921 ( .A1(n13380), .A2(n13061), .ZN(n9929) );
NAND2_X2 U4923 ( .A1(n13303), .A2(n15002), .ZN(n9934) );
NAND2_X2 U4925 ( .A1(n13380), .A2(n13060), .ZN(n9932) );
NAND2_X2 U4927 ( .A1(n13303), .A2(n15016), .ZN(n9937) );
NAND2_X2 U4929 ( .A1(n13380), .A2(n13059), .ZN(n9935) );
NAND2_X2 U4931 ( .A1(n13303), .A2(n15030), .ZN(n9940) );
NAND2_X2 U4933 ( .A1(n13380), .A2(n13058), .ZN(n9938) );
NAND2_X2 U4935 ( .A1(n13303), .A2(n15044), .ZN(n9943) );
NAND2_X2 U4937 ( .A1(n13380), .A2(n13057), .ZN(n9941) );
NAND2_X2 U4939 ( .A1(n13303), .A2(n15058), .ZN(n9946) );
NAND2_X2 U4941 ( .A1(n13380), .A2(n13056), .ZN(n9944) );
NAND2_X2 U4943 ( .A1(n13303), .A2(n15072), .ZN(n9949) );
NAND2_X2 U4945 ( .A1(n13380), .A2(n13055), .ZN(n9947) );
NAND2_X2 U4947 ( .A1(n13303), .A2(n15086), .ZN(n9952) );
NAND2_X2 U4949 ( .A1(n13380), .A2(n13054), .ZN(n9950) );
NAND2_X2 U4951 ( .A1(n13302), .A2(n15100), .ZN(n9955) );
NAND2_X2 U4953 ( .A1(n13380), .A2(n13053), .ZN(n9953) );
NAND2_X2 U4955 ( .A1(n13302), .A2(n15114), .ZN(n9958) );
NAND2_X2 U4957 ( .A1(n13381), .A2(n13052), .ZN(n9956) );
NAND2_X2 U4959 ( .A1(n13302), .A2(n15128), .ZN(n9961) );
NAND2_X2 U4961 ( .A1(n13381), .A2(n13051), .ZN(n9959) );
NAND2_X2 U4963 ( .A1(n13302), .A2(n15142), .ZN(n9964) );
NAND2_X2 U4965 ( .A1(n13381), .A2(n13050), .ZN(n9962) );
NAND2_X2 U4967 ( .A1(n13302), .A2(n15156), .ZN(n9967) );
NAND2_X2 U4969 ( .A1(n13381), .A2(n13049), .ZN(n9965) );
NAND2_X2 U4971 ( .A1(n13302), .A2(n15170), .ZN(n9970) );
NAND2_X2 U4973 ( .A1(n13381), .A2(n13048), .ZN(n9968) );
NAND2_X2 U4975 ( .A1(n13302), .A2(n15184), .ZN(n9973) );
NAND2_X2 U4977 ( .A1(n13381), .A2(n13047), .ZN(n9971) );
NAND2_X2 U4979 ( .A1(n13302), .A2(n15198), .ZN(n9976) );
NAND2_X2 U4981 ( .A1(n13381), .A2(n13046), .ZN(n9974) );
NAND2_X2 U4983 ( .A1(n13302), .A2(n15213), .ZN(n9979) );
NAND2_X2 U4985 ( .A1(n13381), .A2(n13045), .ZN(n9977) );
NAND2_X2 U4987 ( .A1(n13302), .A2(n15228), .ZN(n9982) );
NAND2_X2 U4989 ( .A1(n13381), .A2(n13044), .ZN(n9980) );
NAND2_X2 U4991 ( .A1(n13302), .A2(n15243), .ZN(n9985) );
NAND2_X2 U4993 ( .A1(n13381), .A2(n13043), .ZN(n9983) );
NAND2_X2 U4995 ( .A1(n13301), .A2(n15258), .ZN(n9988) );
NAND2_X2 U4997 ( .A1(n13381), .A2(n13042), .ZN(n9986) );
NAND2_X2 U4999 ( .A1(n13301), .A2(n15273), .ZN(n9991) );
NAND2_X2 U5001 ( .A1(n13382), .A2(n13041), .ZN(n9989) );
NAND2_X2 U5003 ( .A1(n13301), .A2(n15288), .ZN(n9994) );
NAND2_X2 U5005 ( .A1(n13382), .A2(n13040), .ZN(n9992) );
NAND2_X2 U5007 ( .A1(n13301), .A2(n15303), .ZN(n9997) );
NAND2_X2 U5009 ( .A1(n13382), .A2(n13039), .ZN(n9995) );
NAND2_X2 U5011 ( .A1(n13301), .A2(n15318), .ZN(n10000) );
NAND2_X2 U5013 ( .A1(n13382), .A2(n13038), .ZN(n9998) );
NAND2_X2 U5015 ( .A1(n13301), .A2(n15333), .ZN(n10003) );
NAND2_X2 U5017 ( .A1(n13382), .A2(n13037), .ZN(n10001) );
NAND2_X2 U5019 ( .A1(n13301), .A2(n15348), .ZN(n10006) );
NAND2_X2 U5021 ( .A1(n13382), .A2(n13036), .ZN(n10004) );
NAND2_X2 U5023 ( .A1(n13301), .A2(n15363), .ZN(n10009) );
NAND2_X2 U5025 ( .A1(n13382), .A2(n13035), .ZN(n10007) );
NAND2_X2 U5027 ( .A1(n13301), .A2(n15378), .ZN(n10012) );
NAND2_X2 U5029 ( .A1(n13382), .A2(n13034), .ZN(n10010) );
NAND2_X2 U5031 ( .A1(n13301), .A2(n15393), .ZN(n10015) );
NAND2_X2 U5033 ( .A1(n13382), .A2(n13033), .ZN(n10013) );
NAND2_X2 U5035 ( .A1(n13301), .A2(n15408), .ZN(n10018) );
NAND2_X2 U5038 ( .A1(n13382), .A2(n13032), .ZN(n10016) );
NAND2_X2 U5042 ( .A1(n13300), .A2(n15423), .ZN(n10022) );
NAND2_X2 U5044 ( .A1(n13377), .A2(n13063), .ZN(n10020) );
NAND2_X2 U5046 ( .A1(n13300), .A2(n14975), .ZN(n10027) );
NAND2_X2 U5048 ( .A1(n13377), .A2(n13062), .ZN(n10025) );
NAND2_X2 U5050 ( .A1(n13300), .A2(n14989), .ZN(n10030) );
NAND2_X2 U5052 ( .A1(n13377), .A2(n13061), .ZN(n10028) );
NAND2_X2 U5054 ( .A1(n13300), .A2(n15003), .ZN(n10033) );
NAND2_X2 U5056 ( .A1(n13377), .A2(n13060), .ZN(n10031) );
NAND2_X2 U5058 ( .A1(n13300), .A2(n15017), .ZN(n10036) );
NAND2_X2 U5060 ( .A1(n13377), .A2(n13059), .ZN(n10034) );
NAND2_X2 U5062 ( .A1(n13300), .A2(n15031), .ZN(n10039) );
NAND2_X2 U5064 ( .A1(n13377), .A2(n13058), .ZN(n10037) );
NAND2_X2 U5066 ( .A1(n13300), .A2(n15045), .ZN(n10042) );
NAND2_X2 U5068 ( .A1(n13377), .A2(n13057), .ZN(n10040) );
NAND2_X2 U5070 ( .A1(n13300), .A2(n15059), .ZN(n10045) );
NAND2_X2 U5072 ( .A1(n13377), .A2(n13056), .ZN(n10043) );
NAND2_X2 U5074 ( .A1(n13300), .A2(n15073), .ZN(n10048) );
NAND2_X2 U5076 ( .A1(n13377), .A2(n13055), .ZN(n10046) );
NAND2_X2 U5078 ( .A1(n13300), .A2(n15087), .ZN(n10051) );
NAND2_X2 U5080 ( .A1(n13377), .A2(n13054), .ZN(n10049) );
NAND2_X2 U5082 ( .A1(n13300), .A2(n15101), .ZN(n10054) );
NAND2_X2 U5084 ( .A1(n13377), .A2(n13053), .ZN(n10052) );
NAND2_X2 U5086 ( .A1(n13299), .A2(n15115), .ZN(n10057) );
NAND2_X2 U5088 ( .A1(n13378), .A2(n13052), .ZN(n10055) );
NAND2_X2 U5090 ( .A1(n13299), .A2(n15129), .ZN(n10060) );
NAND2_X2 U5092 ( .A1(n13378), .A2(n13051), .ZN(n10058) );
NAND2_X2 U5094 ( .A1(n13299), .A2(n15143), .ZN(n10063) );
NAND2_X2 U5096 ( .A1(n13378), .A2(n13050), .ZN(n10061) );
NAND2_X2 U5098 ( .A1(n13299), .A2(n15157), .ZN(n10066) );
NAND2_X2 U5100 ( .A1(n13378), .A2(n13049), .ZN(n10064) );
NAND2_X2 U5102 ( .A1(n13299), .A2(n15171), .ZN(n10069) );
NAND2_X2 U5104 ( .A1(n13378), .A2(n13048), .ZN(n10067) );
NAND2_X2 U5106 ( .A1(n13299), .A2(n15185), .ZN(n10072) );
NAND2_X2 U5108 ( .A1(n13378), .A2(n13047), .ZN(n10070) );
NAND2_X2 U5110 ( .A1(n13299), .A2(n15199), .ZN(n10075) );
NAND2_X2 U5112 ( .A1(n13378), .A2(n13046), .ZN(n10073) );
NAND2_X2 U5114 ( .A1(n13299), .A2(n15214), .ZN(n10078) );
NAND2_X2 U5116 ( .A1(n13378), .A2(n13045), .ZN(n10076) );
NAND2_X2 U5118 ( .A1(n13299), .A2(n15229), .ZN(n10081) );
NAND2_X2 U5120 ( .A1(n13378), .A2(n13044), .ZN(n10079) );
NAND2_X2 U5122 ( .A1(n13299), .A2(n15244), .ZN(n10084) );
NAND2_X2 U5124 ( .A1(n13378), .A2(n13043), .ZN(n10082) );
NAND2_X2 U5126 ( .A1(n13299), .A2(n15259), .ZN(n10087) );
NAND2_X2 U5128 ( .A1(n13378), .A2(n13042), .ZN(n10085) );
NAND2_X2 U5130 ( .A1(n13298), .A2(n15274), .ZN(n10090) );
NAND2_X2 U5132 ( .A1(n13379), .A2(n13041), .ZN(n10088) );
NAND2_X2 U5134 ( .A1(n13298), .A2(n15289), .ZN(n10093) );
NAND2_X2 U5136 ( .A1(n13379), .A2(n13040), .ZN(n10091) );
NAND2_X2 U5138 ( .A1(n13298), .A2(n15304), .ZN(n10096) );
NAND2_X2 U5140 ( .A1(n13379), .A2(n13039), .ZN(n10094) );
NAND2_X2 U5142 ( .A1(n13298), .A2(n15319), .ZN(n10099) );
NAND2_X2 U5144 ( .A1(n13379), .A2(n13038), .ZN(n10097) );
NAND2_X2 U5146 ( .A1(n13298), .A2(n15334), .ZN(n10102) );
NAND2_X2 U5148 ( .A1(n13379), .A2(n13037), .ZN(n10100) );
NAND2_X2 U5150 ( .A1(n13298), .A2(n15349), .ZN(n10105) );
NAND2_X2 U5152 ( .A1(n13379), .A2(n13036), .ZN(n10103) );
NAND2_X2 U5154 ( .A1(n13298), .A2(n15364), .ZN(n10108) );
NAND2_X2 U5156 ( .A1(n13379), .A2(n13035), .ZN(n10106) );
NAND2_X2 U5158 ( .A1(n13298), .A2(n15379), .ZN(n10111) );
NAND2_X2 U5160 ( .A1(n13379), .A2(n13034), .ZN(n10109) );
NAND2_X2 U5162 ( .A1(n13298), .A2(n15394), .ZN(n10114) );
NAND2_X2 U5164 ( .A1(n13379), .A2(n13033), .ZN(n10112) );
NAND2_X2 U5166 ( .A1(n13298), .A2(n15409), .ZN(n10117) );
NAND2_X2 U5169 ( .A1(n13379), .A2(n13032), .ZN(n10115) );
NAND2_X2 U5173 ( .A1(n13298), .A2(n14976), .ZN(n10121) );
NAND2_X2 U5175 ( .A1(n13062), .A2(n13392), .ZN(n10119) );
NAND2_X2 U5177 ( .A1(n13297), .A2(n14990), .ZN(n10124) );
NAND2_X2 U5179 ( .A1(n13061), .A2(n13392), .ZN(n10122) );
NAND2_X2 U5181 ( .A1(n13297), .A2(n15004), .ZN(n10127) );
NAND2_X2 U5183 ( .A1(n13060), .A2(n13392), .ZN(n10125) );
NAND2_X2 U5185 ( .A1(n13297), .A2(n15018), .ZN(n10130) );
NAND2_X2 U5187 ( .A1(n13059), .A2(n13392), .ZN(n10128) );
NAND2_X2 U5189 ( .A1(n13297), .A2(n15032), .ZN(n10133) );
NAND2_X2 U5191 ( .A1(n13058), .A2(n13392), .ZN(n10131) );
NAND2_X2 U5193 ( .A1(n13297), .A2(n15046), .ZN(n10136) );
NAND2_X2 U5195 ( .A1(n13057), .A2(n13392), .ZN(n10134) );
NAND2_X2 U5197 ( .A1(n13297), .A2(n15060), .ZN(n10139) );
NAND2_X2 U5199 ( .A1(n13056), .A2(n13392), .ZN(n10137) );
NAND2_X2 U5201 ( .A1(n13297), .A2(n15074), .ZN(n10142) );
NAND2_X2 U5203 ( .A1(n13055), .A2(n13392), .ZN(n10140) );
NAND2_X2 U5205 ( .A1(n13297), .A2(n15088), .ZN(n10145) );
NAND2_X2 U5207 ( .A1(n13054), .A2(n13392), .ZN(n10143) );
NAND2_X2 U5209 ( .A1(n13297), .A2(n15102), .ZN(n10148) );
NAND2_X2 U5211 ( .A1(n13053), .A2(n13392), .ZN(n10146) );
NAND2_X2 U5213 ( .A1(n13297), .A2(n15116), .ZN(n10151) );
NAND2_X2 U5215 ( .A1(n13052), .A2(n13393), .ZN(n10149) );
NAND2_X2 U5217 ( .A1(n13297), .A2(n15130), .ZN(n10154) );
NAND2_X2 U5219 ( .A1(n13051), .A2(n13393), .ZN(n10152) );
NAND2_X2 U5221 ( .A1(n13296), .A2(n15144), .ZN(n10157) );
NAND2_X2 U5223 ( .A1(n13050), .A2(n13393), .ZN(n10155) );
NAND2_X2 U5225 ( .A1(n13296), .A2(n15158), .ZN(n10160) );
NAND2_X2 U5227 ( .A1(n13049), .A2(n13393), .ZN(n10158) );
NAND2_X2 U5229 ( .A1(n13296), .A2(n15172), .ZN(n10163) );
NAND2_X2 U5231 ( .A1(n13048), .A2(n13393), .ZN(n10161) );
NAND2_X2 U5233 ( .A1(n13296), .A2(n15186), .ZN(n10166) );
NAND2_X2 U5235 ( .A1(n13047), .A2(n13393), .ZN(n10164) );
NAND2_X2 U5237 ( .A1(n13296), .A2(n15200), .ZN(n10169) );
NAND2_X2 U5239 ( .A1(n13046), .A2(n13393), .ZN(n10167) );
NAND2_X2 U5241 ( .A1(n13296), .A2(n15215), .ZN(n10172) );
NAND2_X2 U5243 ( .A1(n13045), .A2(n13393), .ZN(n10170) );
NAND2_X2 U5245 ( .A1(n13296), .A2(n15230), .ZN(n10175) );
NAND2_X2 U5247 ( .A1(n13044), .A2(n13393), .ZN(n10173) );
NAND2_X2 U5249 ( .A1(n13296), .A2(n15245), .ZN(n10178) );
NAND2_X2 U5251 ( .A1(n13043), .A2(n13393), .ZN(n10176) );
NAND2_X2 U5253 ( .A1(n13296), .A2(n15260), .ZN(n10181) );
NAND2_X2 U5255 ( .A1(n13042), .A2(n13393), .ZN(n10179) );
NAND2_X2 U5257 ( .A1(n13296), .A2(n15275), .ZN(n10184) );
NAND2_X2 U5259 ( .A1(n13041), .A2(n13394), .ZN(n10182) );
NAND2_X2 U5261 ( .A1(n13296), .A2(n15290), .ZN(n10187) );
NAND2_X2 U5263 ( .A1(n13040), .A2(n13394), .ZN(n10185) );
NAND2_X2 U5265 ( .A1(n13295), .A2(n15305), .ZN(n10190) );
NAND2_X2 U5267 ( .A1(n13039), .A2(n13394), .ZN(n10188) );
NAND2_X2 U5269 ( .A1(n13295), .A2(n15320), .ZN(n10193) );
NAND2_X2 U5271 ( .A1(n13038), .A2(n13394), .ZN(n10191) );
NAND2_X2 U5273 ( .A1(n13295), .A2(n15335), .ZN(n10196) );
NAND2_X2 U5275 ( .A1(n13037), .A2(n13394), .ZN(n10194) );
NAND2_X2 U5277 ( .A1(n13295), .A2(n15350), .ZN(n10199) );
NAND2_X2 U5279 ( .A1(n13036), .A2(n13394), .ZN(n10197) );
NAND2_X2 U5281 ( .A1(n13295), .A2(n15365), .ZN(n10202) );
NAND2_X2 U5283 ( .A1(n13035), .A2(n13394), .ZN(n10200) );
NAND2_X2 U5285 ( .A1(n13295), .A2(n15380), .ZN(n10205) );
NAND2_X2 U5287 ( .A1(n13034), .A2(n13394), .ZN(n10203) );
NAND2_X2 U5289 ( .A1(n13295), .A2(n15395), .ZN(n10208) );
NAND2_X2 U5291 ( .A1(n13033), .A2(n13394), .ZN(n10206) );
NAND2_X2 U5293 ( .A1(n13295), .A2(n15410), .ZN(n10211) );
NAND2_X2 U5296 ( .A1(n13032), .A2(n13394), .ZN(n10209) );
NAND2_X2 U5299 ( .A1(n13295), .A2(n14963), .ZN(n10215) );
NAND2_X2 U5301 ( .A1(n13376), .A2(n13063), .ZN(n10213) );
NAND2_X2 U5303 ( .A1(n13295), .A2(n14977), .ZN(n10220) );
NAND2_X2 U5305 ( .A1(n13376), .A2(n13062), .ZN(n10218) );
NAND2_X2 U5307 ( .A1(n13295), .A2(n14991), .ZN(n10223) );
NAND2_X2 U5309 ( .A1(n13376), .A2(n13061), .ZN(n10221) );
NAND2_X2 U5311 ( .A1(n13294), .A2(n15005), .ZN(n10226) );
NAND2_X2 U5313 ( .A1(n13376), .A2(n13060), .ZN(n10224) );
NAND2_X2 U5315 ( .A1(n13294), .A2(n15019), .ZN(n10229) );
NAND2_X2 U5317 ( .A1(n13376), .A2(n13059), .ZN(n10227) );
NAND2_X2 U5319 ( .A1(n13294), .A2(n15033), .ZN(n10232) );
NAND2_X2 U5321 ( .A1(n13376), .A2(n13058), .ZN(n10230) );
NAND2_X2 U5323 ( .A1(n13294), .A2(n15047), .ZN(n10235) );
NAND2_X2 U5325 ( .A1(n13376), .A2(n13057), .ZN(n10233) );
NAND2_X2 U5327 ( .A1(n13294), .A2(n15061), .ZN(n10238) );
NAND2_X2 U5329 ( .A1(n13376), .A2(n13056), .ZN(n10236) );
NAND2_X2 U5331 ( .A1(n13294), .A2(n15075), .ZN(n10241) );
NAND2_X2 U5333 ( .A1(n13376), .A2(n13055), .ZN(n10239) );
NAND2_X2 U5335 ( .A1(n13294), .A2(n15089), .ZN(n10244) );
NAND2_X2 U5337 ( .A1(n13376), .A2(n13054), .ZN(n10242) );
NAND2_X2 U5339 ( .A1(n13294), .A2(n15103), .ZN(n10247) );
NAND2_X2 U5341 ( .A1(n13375), .A2(n13053), .ZN(n10245) );
NAND2_X2 U5343 ( .A1(n13294), .A2(n15117), .ZN(n10250) );
NAND2_X2 U5345 ( .A1(n13375), .A2(n13052), .ZN(n10248) );
NAND2_X2 U5347 ( .A1(n13294), .A2(n15131), .ZN(n10253) );
NAND2_X2 U5349 ( .A1(n13375), .A2(n13051), .ZN(n10251) );
NAND2_X2 U5351 ( .A1(n13294), .A2(n15145), .ZN(n10256) );
NAND2_X2 U5353 ( .A1(n13375), .A2(n13050), .ZN(n10254) );
NAND2_X2 U5355 ( .A1(n13293), .A2(n15159), .ZN(n10259) );
NAND2_X2 U5357 ( .A1(n13375), .A2(n13049), .ZN(n10257) );
NAND2_X2 U5359 ( .A1(n13293), .A2(n15173), .ZN(n10262) );
NAND2_X2 U5361 ( .A1(n13375), .A2(n13048), .ZN(n10260) );
NAND2_X2 U5363 ( .A1(n13293), .A2(n15187), .ZN(n10265) );
NAND2_X2 U5365 ( .A1(n13375), .A2(n13047), .ZN(n10263) );
NAND2_X2 U5367 ( .A1(n13293), .A2(n15201), .ZN(n10268) );
NAND2_X2 U5369 ( .A1(n13375), .A2(n13046), .ZN(n10266) );
NAND2_X2 U5371 ( .A1(n13293), .A2(n15216), .ZN(n10271) );
NAND2_X2 U5373 ( .A1(n13375), .A2(n13045), .ZN(n10269) );
NAND2_X2 U5375 ( .A1(n13293), .A2(n15231), .ZN(n10274) );
NAND2_X2 U5377 ( .A1(n13375), .A2(n13044), .ZN(n10272) );
NAND2_X2 U5379 ( .A1(n13293), .A2(n15246), .ZN(n10277) );
NAND2_X2 U5381 ( .A1(n13375), .A2(n13043), .ZN(n10275) );
NAND2_X2 U5383 ( .A1(n13293), .A2(n15261), .ZN(n10280) );
NAND2_X2 U5385 ( .A1(n13374), .A2(n13042), .ZN(n10278) );
NAND2_X2 U5387 ( .A1(n13293), .A2(n15276), .ZN(n10283) );
NAND2_X2 U5389 ( .A1(n13374), .A2(n13041), .ZN(n10281) );
NAND2_X2 U5391 ( .A1(n13293), .A2(n15291), .ZN(n10286) );
NAND2_X2 U5393 ( .A1(n13374), .A2(n13040), .ZN(n10284) );
NAND2_X2 U5395 ( .A1(n13293), .A2(n15306), .ZN(n10289) );
NAND2_X2 U5397 ( .A1(n13374), .A2(n13039), .ZN(n10287) );
NAND2_X2 U5399 ( .A1(n13292), .A2(n15321), .ZN(n10292) );
NAND2_X2 U5401 ( .A1(n13374), .A2(n13038), .ZN(n10290) );
NAND2_X2 U5403 ( .A1(n13292), .A2(n15336), .ZN(n10295) );
NAND2_X2 U5405 ( .A1(n13374), .A2(n13037), .ZN(n10293) );
NAND2_X2 U5407 ( .A1(n13292), .A2(n15351), .ZN(n10298) );
NAND2_X2 U5409 ( .A1(n13374), .A2(n13036), .ZN(n10296) );
NAND2_X2 U5411 ( .A1(n13292), .A2(n15366), .ZN(n10301) );
NAND2_X2 U5413 ( .A1(n13374), .A2(n13035), .ZN(n10299) );
NAND2_X2 U5415 ( .A1(n13292), .A2(n15381), .ZN(n10304) );
NAND2_X2 U5417 ( .A1(n13374), .A2(n13034), .ZN(n10302) );
NAND2_X2 U5419 ( .A1(n13292), .A2(n15396), .ZN(n10307) );
NAND2_X2 U5421 ( .A1(n13374), .A2(n13033), .ZN(n10305) );
NAND2_X2 U5423 ( .A1(n13292), .A2(n15411), .ZN(n10310) );
NAND2_X2 U5427 ( .A1(n13374), .A2(n13032), .ZN(n10308) );
NAND2_X2 U5430 ( .A1(n13292), .A2(n14964), .ZN(n10315) );
NAND2_X2 U5432 ( .A1(n13371), .A2(n13063), .ZN(n10313) );
NAND2_X2 U5434 ( .A1(n13292), .A2(n14978), .ZN(n10320) );
NAND2_X2 U5436 ( .A1(n13371), .A2(n13062), .ZN(n10318) );
NAND2_X2 U5438 ( .A1(n13292), .A2(n14992), .ZN(n10323) );
NAND2_X2 U5440 ( .A1(n13371), .A2(n13061), .ZN(n10321) );
NAND2_X2 U5442 ( .A1(n13292), .A2(n15006), .ZN(n10326) );
NAND2_X2 U5444 ( .A1(n13371), .A2(n13060), .ZN(n10324) );
NAND2_X2 U5446 ( .A1(n13291), .A2(n15020), .ZN(n10329) );
NAND2_X2 U5448 ( .A1(n13371), .A2(n13059), .ZN(n10327) );
NAND2_X2 U5450 ( .A1(n13291), .A2(n15034), .ZN(n10332) );
NAND2_X2 U5452 ( .A1(n13371), .A2(n13058), .ZN(n10330) );
NAND2_X2 U5454 ( .A1(n13291), .A2(n15048), .ZN(n10335) );
NAND2_X2 U5456 ( .A1(n13371), .A2(n13057), .ZN(n10333) );
NAND2_X2 U5458 ( .A1(n13291), .A2(n15062), .ZN(n10338) );
NAND2_X2 U5460 ( .A1(n13371), .A2(n13056), .ZN(n10336) );
NAND2_X2 U5462 ( .A1(n13291), .A2(n15076), .ZN(n10341) );
NAND2_X2 U5464 ( .A1(n13371), .A2(n13055), .ZN(n10339) );
NAND2_X2 U5466 ( .A1(n13291), .A2(n15090), .ZN(n10344) );
NAND2_X2 U5468 ( .A1(n13371), .A2(n13054), .ZN(n10342) );
NAND2_X2 U5470 ( .A1(n13291), .A2(n15104), .ZN(n10347) );
NAND2_X2 U5472 ( .A1(n13371), .A2(n13053), .ZN(n10345) );
NAND2_X2 U5474 ( .A1(n13291), .A2(n15118), .ZN(n10350) );
NAND2_X2 U5476 ( .A1(n13372), .A2(n13052), .ZN(n10348) );
NAND2_X2 U5478 ( .A1(n13291), .A2(n15132), .ZN(n10353) );
NAND2_X2 U5480 ( .A1(n13372), .A2(n13051), .ZN(n10351) );
NAND2_X2 U5482 ( .A1(n13291), .A2(n15146), .ZN(n10356) );
NAND2_X2 U5484 ( .A1(n13372), .A2(n13050), .ZN(n10354) );
NAND2_X2 U5486 ( .A1(n13291), .A2(n15160), .ZN(n10359) );
NAND2_X2 U5488 ( .A1(n13372), .A2(n13049), .ZN(n10357) );
NAND2_X2 U5490 ( .A1(n13290), .A2(n15174), .ZN(n10362) );
NAND2_X2 U5492 ( .A1(n13372), .A2(n13048), .ZN(n10360) );
NAND2_X2 U5494 ( .A1(n13290), .A2(n15188), .ZN(n10365) );
NAND2_X2 U5496 ( .A1(n13372), .A2(n13047), .ZN(n10363) );
NAND2_X2 U5498 ( .A1(n13290), .A2(n15202), .ZN(n10368) );
NAND2_X2 U5500 ( .A1(n13372), .A2(n13046), .ZN(n10366) );
NAND2_X2 U5502 ( .A1(n13290), .A2(n15217), .ZN(n10371) );
NAND2_X2 U5504 ( .A1(n13372), .A2(n13045), .ZN(n10369) );
NAND2_X2 U5506 ( .A1(n13290), .A2(n15232), .ZN(n10374) );
NAND2_X2 U5508 ( .A1(n13372), .A2(n13044), .ZN(n10372) );
NAND2_X2 U5510 ( .A1(n13290), .A2(n15247), .ZN(n10377) );
NAND2_X2 U5512 ( .A1(n13372), .A2(n13043), .ZN(n10375) );
NAND2_X2 U5514 ( .A1(n13290), .A2(n15262), .ZN(n10380) );
NAND2_X2 U5516 ( .A1(n13372), .A2(n13042), .ZN(n10378) );
NAND2_X2 U5518 ( .A1(n13290), .A2(n15277), .ZN(n10383) );
NAND2_X2 U5520 ( .A1(n13373), .A2(n13041), .ZN(n10381) );
NAND2_X2 U5522 ( .A1(n13290), .A2(n15292), .ZN(n10386) );
NAND2_X2 U5524 ( .A1(n13373), .A2(n13040), .ZN(n10384) );
NAND2_X2 U5526 ( .A1(n13290), .A2(n15307), .ZN(n10389) );
NAND2_X2 U5528 ( .A1(n13373), .A2(n13039), .ZN(n10387) );
NAND2_X2 U5530 ( .A1(n13290), .A2(n15322), .ZN(n10392) );
NAND2_X2 U5532 ( .A1(n13373), .A2(n13038), .ZN(n10390) );
NAND2_X2 U5534 ( .A1(n13289), .A2(n15337), .ZN(n10395) );
NAND2_X2 U5536 ( .A1(n13373), .A2(n13037), .ZN(n10393) );
NAND2_X2 U5538 ( .A1(n13289), .A2(n15352), .ZN(n10398) );
NAND2_X2 U5540 ( .A1(n13373), .A2(n13036), .ZN(n10396) );
NAND2_X2 U5542 ( .A1(n13289), .A2(n15367), .ZN(n10401) );
NAND2_X2 U5544 ( .A1(n13373), .A2(n13035), .ZN(n10399) );
NAND2_X2 U5546 ( .A1(n13289), .A2(n15382), .ZN(n10404) );
NAND2_X2 U5548 ( .A1(n13373), .A2(n13034), .ZN(n10402) );
NAND2_X2 U5550 ( .A1(n13289), .A2(n15397), .ZN(n10407) );
NAND2_X2 U5552 ( .A1(n13373), .A2(n13033), .ZN(n10405) );
NAND2_X2 U5554 ( .A1(n13289), .A2(n15412), .ZN(n10410) );
NAND2_X2 U5557 ( .A1(n13373), .A2(n13032), .ZN(n10408) );
NAND2_X2 U5561 ( .A1(n13289), .A2(n14965), .ZN(n10414) );
NAND2_X2 U5563 ( .A1(n13368), .A2(n13063), .ZN(n10412) );
NAND2_X2 U5565 ( .A1(n13289), .A2(n14979), .ZN(n10419) );
NAND2_X2 U5567 ( .A1(n13368), .A2(n13062), .ZN(n10417) );
NAND2_X2 U5569 ( .A1(n13289), .A2(n14993), .ZN(n10422) );
NAND2_X2 U5571 ( .A1(n13368), .A2(n13061), .ZN(n10420) );
NAND2_X2 U5573 ( .A1(n13289), .A2(n15007), .ZN(n10425) );
NAND2_X2 U5575 ( .A1(n13368), .A2(n13060), .ZN(n10423) );
NAND2_X2 U5577 ( .A1(n13289), .A2(n15021), .ZN(n10428) );
NAND2_X2 U5579 ( .A1(n13368), .A2(n13059), .ZN(n10426) );
NAND2_X2 U5581 ( .A1(n13288), .A2(n15035), .ZN(n10431) );
NAND2_X2 U5583 ( .A1(n13368), .A2(n13058), .ZN(n10429) );
NAND2_X2 U5585 ( .A1(n13288), .A2(n15049), .ZN(n10434) );
NAND2_X2 U5587 ( .A1(n13368), .A2(n13057), .ZN(n10432) );
NAND2_X2 U5589 ( .A1(n13288), .A2(n15063), .ZN(n10437) );
NAND2_X2 U5591 ( .A1(n13368), .A2(n13056), .ZN(n10435) );
NAND2_X2 U5593 ( .A1(n13288), .A2(n15077), .ZN(n10440) );
NAND2_X2 U5595 ( .A1(n13368), .A2(n13055), .ZN(n10438) );
NAND2_X2 U5597 ( .A1(n13288), .A2(n15091), .ZN(n10443) );
NAND2_X2 U5599 ( .A1(n13368), .A2(n13054), .ZN(n10441) );
NAND2_X2 U5601 ( .A1(n13288), .A2(n15105), .ZN(n10446) );
NAND2_X2 U5603 ( .A1(n13368), .A2(n13053), .ZN(n10444) );
NAND2_X2 U5605 ( .A1(n13288), .A2(n15119), .ZN(n10449) );
NAND2_X2 U5607 ( .A1(n13369), .A2(n13052), .ZN(n10447) );
NAND2_X2 U5609 ( .A1(n13288), .A2(n15133), .ZN(n10452) );
NAND2_X2 U5611 ( .A1(n13369), .A2(n13051), .ZN(n10450) );
NAND2_X2 U5613 ( .A1(n13288), .A2(n15147), .ZN(n10455) );
NAND2_X2 U5615 ( .A1(n13369), .A2(n13050), .ZN(n10453) );
NAND2_X2 U5617 ( .A1(n13288), .A2(n15161), .ZN(n10458) );
NAND2_X2 U5619 ( .A1(n13369), .A2(n13049), .ZN(n10456) );
NAND2_X2 U5621 ( .A1(n13288), .A2(n15175), .ZN(n10461) );
NAND2_X2 U5623 ( .A1(n13369), .A2(n13048), .ZN(n10459) );
NAND2_X2 U5625 ( .A1(n13287), .A2(n15189), .ZN(n10464) );
NAND2_X2 U5627 ( .A1(n13369), .A2(n13047), .ZN(n10462) );
NAND2_X2 U5629 ( .A1(n13287), .A2(n15203), .ZN(n10467) );
NAND2_X2 U5631 ( .A1(n13369), .A2(n13046), .ZN(n10465) );
NAND2_X2 U5633 ( .A1(n13287), .A2(n15218), .ZN(n10470) );
NAND2_X2 U5635 ( .A1(n13369), .A2(n13045), .ZN(n10468) );
NAND2_X2 U5637 ( .A1(n13287), .A2(n15233), .ZN(n10473) );
NAND2_X2 U5639 ( .A1(n13369), .A2(n13044), .ZN(n10471) );
NAND2_X2 U5641 ( .A1(n13287), .A2(n15248), .ZN(n10476) );
NAND2_X2 U5643 ( .A1(n13369), .A2(n13043), .ZN(n10474) );
NAND2_X2 U5645 ( .A1(n13287), .A2(n15263), .ZN(n10479) );
NAND2_X2 U5647 ( .A1(n13369), .A2(n13042), .ZN(n10477) );
NAND2_X2 U5649 ( .A1(n13287), .A2(n15278), .ZN(n10482) );
NAND2_X2 U5651 ( .A1(n13370), .A2(n13041), .ZN(n10480) );
NAND2_X2 U5653 ( .A1(n13287), .A2(n15293), .ZN(n10485) );
NAND2_X2 U5655 ( .A1(n13370), .A2(n13040), .ZN(n10483) );
NAND2_X2 U5657 ( .A1(n13287), .A2(n15308), .ZN(n10488) );
NAND2_X2 U5659 ( .A1(n13370), .A2(n13039), .ZN(n10486) );
NAND2_X2 U5661 ( .A1(n13287), .A2(n15323), .ZN(n10491) );
NAND2_X2 U5663 ( .A1(n13370), .A2(n13038), .ZN(n10489) );
NAND2_X2 U5665 ( .A1(n13287), .A2(n15338), .ZN(n10494) );
NAND2_X2 U5667 ( .A1(n13370), .A2(n13037), .ZN(n10492) );
NAND2_X2 U5669 ( .A1(n13286), .A2(n15353), .ZN(n10497) );
NAND2_X2 U5671 ( .A1(n13370), .A2(n13036), .ZN(n10495) );
NAND2_X2 U5673 ( .A1(n13286), .A2(n15368), .ZN(n10500) );
NAND2_X2 U5675 ( .A1(n13370), .A2(n13035), .ZN(n10498) );
NAND2_X2 U5677 ( .A1(n13286), .A2(n15383), .ZN(n10503) );
NAND2_X2 U5679 ( .A1(n13370), .A2(n13034), .ZN(n10501) );
NAND2_X2 U5681 ( .A1(n13286), .A2(n15398), .ZN(n10506) );
NAND2_X2 U5683 ( .A1(n13370), .A2(n13033), .ZN(n10504) );
NAND2_X2 U5685 ( .A1(n13286), .A2(n15413), .ZN(n10509) );
NAND2_X2 U5688 ( .A1(n13370), .A2(n13032), .ZN(n10507) );
NAND2_X2 U5692 ( .A1(n13286), .A2(n14966), .ZN(n10513) );
NAND2_X2 U5694 ( .A1(n13365), .A2(n13063), .ZN(n10511) );
NAND2_X2 U5696 ( .A1(n13286), .A2(n14980), .ZN(n10518) );
NAND2_X2 U5698 ( .A1(n13365), .A2(n13062), .ZN(n10516) );
NAND2_X2 U5700 ( .A1(n13286), .A2(n14994), .ZN(n10521) );
NAND2_X2 U5702 ( .A1(n13365), .A2(n13061), .ZN(n10519) );
NAND2_X2 U5704 ( .A1(n13286), .A2(n15008), .ZN(n10524) );
NAND2_X2 U5706 ( .A1(n13365), .A2(n13060), .ZN(n10522) );
NAND2_X2 U5708 ( .A1(n13286), .A2(n15022), .ZN(n10527) );
NAND2_X2 U5710 ( .A1(n13365), .A2(n13059), .ZN(n10525) );
NAND2_X2 U5712 ( .A1(n13286), .A2(n15036), .ZN(n10530) );
NAND2_X2 U5714 ( .A1(n13365), .A2(n13058), .ZN(n10528) );
NAND2_X2 U5716 ( .A1(n13285), .A2(n15050), .ZN(n10533) );
NAND2_X2 U5718 ( .A1(n13365), .A2(n13057), .ZN(n10531) );
NAND2_X2 U5720 ( .A1(n13285), .A2(n15064), .ZN(n10536) );
NAND2_X2 U5722 ( .A1(n13365), .A2(n13056), .ZN(n10534) );
NAND2_X2 U5724 ( .A1(n13285), .A2(n15078), .ZN(n10539) );
NAND2_X2 U5726 ( .A1(n13365), .A2(n13055), .ZN(n10537) );
NAND2_X2 U5728 ( .A1(n13285), .A2(n15092), .ZN(n10542) );
NAND2_X2 U5730 ( .A1(n13365), .A2(n13054), .ZN(n10540) );
NAND2_X2 U5732 ( .A1(n13285), .A2(n15106), .ZN(n10545) );
NAND2_X2 U5734 ( .A1(n13365), .A2(n13053), .ZN(n10543) );
NAND2_X2 U5736 ( .A1(n13285), .A2(n15120), .ZN(n10548) );
NAND2_X2 U5738 ( .A1(n13366), .A2(n13052), .ZN(n10546) );
NAND2_X2 U5740 ( .A1(n13285), .A2(n15134), .ZN(n10551) );
NAND2_X2 U5742 ( .A1(n13366), .A2(n13051), .ZN(n10549) );
NAND2_X2 U5744 ( .A1(n13285), .A2(n15148), .ZN(n10554) );
NAND2_X2 U5746 ( .A1(n13366), .A2(n13050), .ZN(n10552) );
NAND2_X2 U5748 ( .A1(n13285), .A2(n15162), .ZN(n10557) );
NAND2_X2 U5750 ( .A1(n13366), .A2(n13049), .ZN(n10555) );
NAND2_X2 U5752 ( .A1(n13285), .A2(n15176), .ZN(n10560) );
NAND2_X2 U5754 ( .A1(n13366), .A2(n13048), .ZN(n10558) );
NAND2_X2 U5756 ( .A1(n13285), .A2(n15190), .ZN(n10563) );
NAND2_X2 U5758 ( .A1(n13366), .A2(n13047), .ZN(n10561) );
NAND2_X2 U5760 ( .A1(n13284), .A2(n15204), .ZN(n10566) );
NAND2_X2 U5762 ( .A1(n13366), .A2(n13046), .ZN(n10564) );
NAND2_X2 U5764 ( .A1(n13284), .A2(n15219), .ZN(n10569) );
NAND2_X2 U5766 ( .A1(n13366), .A2(n13045), .ZN(n10567) );
NAND2_X2 U5768 ( .A1(n13284), .A2(n15234), .ZN(n10572) );
NAND2_X2 U5770 ( .A1(n13366), .A2(n13044), .ZN(n10570) );
NAND2_X2 U5772 ( .A1(n13284), .A2(n15249), .ZN(n10575) );
NAND2_X2 U5774 ( .A1(n13366), .A2(n13043), .ZN(n10573) );
NAND2_X2 U5776 ( .A1(n13284), .A2(n15264), .ZN(n10578) );
NAND2_X2 U5778 ( .A1(n13366), .A2(n13042), .ZN(n10576) );
NAND2_X2 U5780 ( .A1(n13284), .A2(n15279), .ZN(n10581) );
NAND2_X2 U5782 ( .A1(n13367), .A2(n13041), .ZN(n10579) );
NAND2_X2 U5784 ( .A1(n13284), .A2(n15294), .ZN(n10584) );
NAND2_X2 U5786 ( .A1(n13367), .A2(n13040), .ZN(n10582) );
NAND2_X2 U5788 ( .A1(n13284), .A2(n15309), .ZN(n10587) );
NAND2_X2 U5790 ( .A1(n13367), .A2(n13039), .ZN(n10585) );
NAND2_X2 U5792 ( .A1(n13284), .A2(n15324), .ZN(n10590) );
NAND2_X2 U5794 ( .A1(n13367), .A2(n13038), .ZN(n10588) );
NAND2_X2 U5796 ( .A1(n13284), .A2(n15339), .ZN(n10593) );
NAND2_X2 U5798 ( .A1(n13367), .A2(n13037), .ZN(n10591) );
NAND2_X2 U5800 ( .A1(n13284), .A2(n15354), .ZN(n10596) );
NAND2_X2 U5802 ( .A1(n13367), .A2(n13036), .ZN(n10594) );
NAND2_X2 U5804 ( .A1(n13283), .A2(n15369), .ZN(n10599) );
NAND2_X2 U5806 ( .A1(n13367), .A2(n13035), .ZN(n10597) );
NAND2_X2 U5808 ( .A1(n13283), .A2(n15384), .ZN(n10602) );
NAND2_X2 U5810 ( .A1(n13367), .A2(n13034), .ZN(n10600) );
NAND2_X2 U5812 ( .A1(n13283), .A2(n15399), .ZN(n10605) );
NAND2_X2 U5814 ( .A1(n13367), .A2(n13033), .ZN(n10603) );
NAND2_X2 U5816 ( .A1(n13283), .A2(n15414), .ZN(n10608) );
NAND2_X2 U5819 ( .A1(n13367), .A2(n13032), .ZN(n10606) );
NAND2_X2 U5822 ( .A1(n13283), .A2(n14967), .ZN(n10612) );
NAND2_X2 U5824 ( .A1(n13364), .A2(n13063), .ZN(n10610) );
NAND2_X2 U5826 ( .A1(n13283), .A2(n14981), .ZN(n10617) );
NAND2_X2 U5828 ( .A1(n13364), .A2(n13062), .ZN(n10615) );
NAND2_X2 U5830 ( .A1(n13283), .A2(n14995), .ZN(n10620) );
NAND2_X2 U5832 ( .A1(n13364), .A2(n13061), .ZN(n10618) );
NAND2_X2 U5834 ( .A1(n13283), .A2(n15009), .ZN(n10623) );
NAND2_X2 U5836 ( .A1(n13364), .A2(n13060), .ZN(n10621) );
NAND2_X2 U5838 ( .A1(n13283), .A2(n15023), .ZN(n10626) );
NAND2_X2 U5840 ( .A1(n13364), .A2(n13059), .ZN(n10624) );
NAND2_X2 U5842 ( .A1(n13283), .A2(n15037), .ZN(n10629) );
NAND2_X2 U5844 ( .A1(n13364), .A2(n13058), .ZN(n10627) );
NAND2_X2 U5846 ( .A1(n13283), .A2(n15051), .ZN(n10632) );
NAND2_X2 U5848 ( .A1(n13364), .A2(n13057), .ZN(n10630) );
NAND2_X2 U5850 ( .A1(n13282), .A2(n15065), .ZN(n10635) );
NAND2_X2 U5852 ( .A1(n13364), .A2(n13056), .ZN(n10633) );
NAND2_X2 U5854 ( .A1(n13282), .A2(n15079), .ZN(n10638) );
NAND2_X2 U5856 ( .A1(n13364), .A2(n13055), .ZN(n10636) );
NAND2_X2 U5858 ( .A1(n13282), .A2(n15093), .ZN(n10641) );
NAND2_X2 U5860 ( .A1(n13364), .A2(n13054), .ZN(n10639) );
NAND2_X2 U5862 ( .A1(n13282), .A2(n15107), .ZN(n10644) );
NAND2_X2 U5864 ( .A1(n13363), .A2(n13053), .ZN(n10642) );
NAND2_X2 U5866 ( .A1(n13282), .A2(n15121), .ZN(n10647) );
NAND2_X2 U5868 ( .A1(n13363), .A2(n13052), .ZN(n10645) );
NAND2_X2 U5870 ( .A1(n13282), .A2(n15135), .ZN(n10650) );
NAND2_X2 U5872 ( .A1(n13363), .A2(n13051), .ZN(n10648) );
NAND2_X2 U5874 ( .A1(n13282), .A2(n15149), .ZN(n10653) );
NAND2_X2 U5876 ( .A1(n13363), .A2(n13050), .ZN(n10651) );
NAND2_X2 U5878 ( .A1(n13282), .A2(n15163), .ZN(n10656) );
NAND2_X2 U5880 ( .A1(n13363), .A2(n13049), .ZN(n10654) );
NAND2_X2 U5882 ( .A1(n13282), .A2(n15177), .ZN(n10659) );
NAND2_X2 U5884 ( .A1(n13363), .A2(n13048), .ZN(n10657) );
NAND2_X2 U5886 ( .A1(n13282), .A2(n15191), .ZN(n10662) );
NAND2_X2 U5888 ( .A1(n13363), .A2(n13047), .ZN(n10660) );
NAND2_X2 U5890 ( .A1(n13282), .A2(n15205), .ZN(n10665) );
NAND2_X2 U5892 ( .A1(n13363), .A2(n13046), .ZN(n10663) );
NAND2_X2 U5894 ( .A1(n13281), .A2(n15220), .ZN(n10668) );
NAND2_X2 U5896 ( .A1(n13363), .A2(n13045), .ZN(n10666) );
NAND2_X2 U5898 ( .A1(n13281), .A2(n15235), .ZN(n10671) );
NAND2_X2 U5900 ( .A1(n13363), .A2(n13044), .ZN(n10669) );
NAND2_X2 U5902 ( .A1(n13281), .A2(n15250), .ZN(n10674) );
NAND2_X2 U5904 ( .A1(n13363), .A2(n13043), .ZN(n10672) );
NAND2_X2 U5906 ( .A1(n13281), .A2(n15265), .ZN(n10677) );
NAND2_X2 U5908 ( .A1(n13362), .A2(n13042), .ZN(n10675) );
NAND2_X2 U5910 ( .A1(n13281), .A2(n15280), .ZN(n10680) );
NAND2_X2 U5912 ( .A1(n13362), .A2(n13041), .ZN(n10678) );
NAND2_X2 U5914 ( .A1(n13281), .A2(n15295), .ZN(n10683) );
NAND2_X2 U5916 ( .A1(n13362), .A2(n13040), .ZN(n10681) );
NAND2_X2 U5918 ( .A1(n13281), .A2(n15310), .ZN(n10686) );
NAND2_X2 U5920 ( .A1(n13362), .A2(n13039), .ZN(n10684) );
NAND2_X2 U5922 ( .A1(n13281), .A2(n15325), .ZN(n10689) );
NAND2_X2 U5924 ( .A1(n13362), .A2(n13038), .ZN(n10687) );
NAND2_X2 U5926 ( .A1(n13281), .A2(n15340), .ZN(n10692) );
NAND2_X2 U5928 ( .A1(n13362), .A2(n13037), .ZN(n10690) );
NAND2_X2 U5930 ( .A1(n13281), .A2(n15355), .ZN(n10695) );
NAND2_X2 U5932 ( .A1(n13362), .A2(n13036), .ZN(n10693) );
NAND2_X2 U5934 ( .A1(n13281), .A2(n15370), .ZN(n10698) );
NAND2_X2 U5936 ( .A1(n13362), .A2(n13035), .ZN(n10696) );
NAND2_X2 U5938 ( .A1(n13280), .A2(n15385), .ZN(n10701) );
NAND2_X2 U5940 ( .A1(n13362), .A2(n13034), .ZN(n10699) );
NAND2_X2 U5942 ( .A1(n13280), .A2(n15400), .ZN(n10704) );
NAND2_X2 U5944 ( .A1(n13362), .A2(n13033), .ZN(n10702) );
NAND2_X2 U5946 ( .A1(n13280), .A2(n15415), .ZN(n10707) );
NAND2_X2 U5950 ( .A1(n13362), .A2(n13032), .ZN(n10705) );
NAND2_X2 U5953 ( .A1(n13280), .A2(n14968), .ZN(n10713) );
NAND2_X2 U5955 ( .A1(n13361), .A2(n13063), .ZN(n10711) );
NAND2_X2 U5957 ( .A1(n13280), .A2(n14982), .ZN(n10718) );
NAND2_X2 U5959 ( .A1(n13361), .A2(n13062), .ZN(n10716) );
NAND2_X2 U5961 ( .A1(n13280), .A2(n14996), .ZN(n10721) );
NAND2_X2 U5963 ( .A1(n13361), .A2(n13061), .ZN(n10719) );
NAND2_X2 U5965 ( .A1(n13280), .A2(n15010), .ZN(n10724) );
NAND2_X2 U5967 ( .A1(n13361), .A2(n13060), .ZN(n10722) );
NAND2_X2 U5969 ( .A1(n13280), .A2(n15024), .ZN(n10727) );
NAND2_X2 U5971 ( .A1(n13361), .A2(n13059), .ZN(n10725) );
NAND2_X2 U5973 ( .A1(n13280), .A2(n15038), .ZN(n10730) );
NAND2_X2 U5975 ( .A1(n13361), .A2(n13058), .ZN(n10728) );
NAND2_X2 U5977 ( .A1(n13280), .A2(n15052), .ZN(n10733) );
NAND2_X2 U5979 ( .A1(n13361), .A2(n13057), .ZN(n10731) );
NAND2_X2 U5981 ( .A1(n13280), .A2(n15066), .ZN(n10736) );
NAND2_X2 U5983 ( .A1(n13361), .A2(n13056), .ZN(n10734) );
NAND2_X2 U5985 ( .A1(n13279), .A2(n15080), .ZN(n10739) );
NAND2_X2 U5987 ( .A1(n13361), .A2(n13055), .ZN(n10737) );
NAND2_X2 U5989 ( .A1(n13279), .A2(n15094), .ZN(n10742) );
NAND2_X2 U5991 ( .A1(n13361), .A2(n13054), .ZN(n10740) );
NAND2_X2 U5993 ( .A1(n13279), .A2(n15108), .ZN(n10745) );
NAND2_X2 U5995 ( .A1(n13360), .A2(n13053), .ZN(n10743) );
NAND2_X2 U5997 ( .A1(n13279), .A2(n15122), .ZN(n10748) );
NAND2_X2 U5999 ( .A1(n13360), .A2(n13052), .ZN(n10746) );
NAND2_X2 U6001 ( .A1(n13279), .A2(n15136), .ZN(n10751) );
NAND2_X2 U6003 ( .A1(n13360), .A2(n13051), .ZN(n10749) );
NAND2_X2 U6005 ( .A1(n13279), .A2(n15150), .ZN(n10754) );
NAND2_X2 U6007 ( .A1(n13360), .A2(n13050), .ZN(n10752) );
NAND2_X2 U6009 ( .A1(n13279), .A2(n15164), .ZN(n10757) );
NAND2_X2 U6011 ( .A1(n13360), .A2(n13049), .ZN(n10755) );
NAND2_X2 U6013 ( .A1(n13279), .A2(n15178), .ZN(n10760) );
NAND2_X2 U6015 ( .A1(n13360), .A2(n13048), .ZN(n10758) );
NAND2_X2 U6017 ( .A1(n13279), .A2(n15192), .ZN(n10763) );
NAND2_X2 U6019 ( .A1(n13360), .A2(n13047), .ZN(n10761) );
NAND2_X2 U6021 ( .A1(n13279), .A2(n15206), .ZN(n10766) );
NAND2_X2 U6023 ( .A1(n13360), .A2(n13046), .ZN(n10764) );
NAND2_X2 U6025 ( .A1(n13279), .A2(n15221), .ZN(n10769) );
NAND2_X2 U6027 ( .A1(n13360), .A2(n13045), .ZN(n10767) );
NAND2_X2 U6029 ( .A1(n13278), .A2(n15236), .ZN(n10772) );
NAND2_X2 U6031 ( .A1(n13360), .A2(n13044), .ZN(n10770) );
NAND2_X2 U6033 ( .A1(n13278), .A2(n15251), .ZN(n10775) );
NAND2_X2 U6035 ( .A1(n13360), .A2(n13043), .ZN(n10773) );
NAND2_X2 U6037 ( .A1(n13278), .A2(n15266), .ZN(n10778) );
NAND2_X2 U6039 ( .A1(n13359), .A2(n13042), .ZN(n10776) );
NAND2_X2 U6041 ( .A1(n13278), .A2(n15281), .ZN(n10781) );
NAND2_X2 U6043 ( .A1(n13359), .A2(n13041), .ZN(n10779) );
NAND2_X2 U6045 ( .A1(n13278), .A2(n15296), .ZN(n10784) );
NAND2_X2 U6047 ( .A1(n13359), .A2(n13040), .ZN(n10782) );
NAND2_X2 U6049 ( .A1(n13278), .A2(n15311), .ZN(n10787) );
NAND2_X2 U6051 ( .A1(n13359), .A2(n13039), .ZN(n10785) );
NAND2_X2 U6053 ( .A1(n13278), .A2(n15326), .ZN(n10790) );
NAND2_X2 U6055 ( .A1(n13359), .A2(n13038), .ZN(n10788) );
NAND2_X2 U6057 ( .A1(n13278), .A2(n15341), .ZN(n10793) );
NAND2_X2 U6059 ( .A1(n13359), .A2(n13037), .ZN(n10791) );
NAND2_X2 U6061 ( .A1(n13278), .A2(n15356), .ZN(n10796) );
NAND2_X2 U6063 ( .A1(n13359), .A2(n13036), .ZN(n10794) );
NAND2_X2 U6065 ( .A1(n13278), .A2(n15371), .ZN(n10799) );
NAND2_X2 U6067 ( .A1(n13359), .A2(n13035), .ZN(n10797) );
NAND2_X2 U6069 ( .A1(n13278), .A2(n15386), .ZN(n10802) );
NAND2_X2 U6071 ( .A1(n13359), .A2(n13034), .ZN(n10800) );
NAND2_X2 U6073 ( .A1(n13277), .A2(n15401), .ZN(n10805) );
NAND2_X2 U6075 ( .A1(n13359), .A2(n13033), .ZN(n10803) );
NAND2_X2 U6077 ( .A1(n13277), .A2(n15416), .ZN(n10808) );
NAND2_X2 U6081 ( .A1(n13359), .A2(n13032), .ZN(n10806) );
NAND2_X2 U6084 ( .A1(n13277), .A2(n14969), .ZN(n10812) );
NAND2_X2 U6086 ( .A1(n13358), .A2(n13063), .ZN(n10810) );
NAND2_X2 U6088 ( .A1(n13277), .A2(n14983), .ZN(n10817) );
NAND2_X2 U6090 ( .A1(n13358), .A2(n13062), .ZN(n10815) );
NAND2_X2 U6092 ( .A1(n13277), .A2(n14997), .ZN(n10820) );
NAND2_X2 U6094 ( .A1(n13358), .A2(n13061), .ZN(n10818) );
NAND2_X2 U6096 ( .A1(n13277), .A2(n15011), .ZN(n10823) );
NAND2_X2 U6098 ( .A1(n13358), .A2(n13060), .ZN(n10821) );
NAND2_X2 U6100 ( .A1(n13277), .A2(n15025), .ZN(n10826) );
NAND2_X2 U6102 ( .A1(n13358), .A2(n13059), .ZN(n10824) );
NAND2_X2 U6104 ( .A1(n13277), .A2(n15039), .ZN(n10829) );
NAND2_X2 U6106 ( .A1(n13358), .A2(n13058), .ZN(n10827) );
NAND2_X2 U6108 ( .A1(n13277), .A2(n15053), .ZN(n10832) );
NAND2_X2 U6110 ( .A1(n13358), .A2(n13057), .ZN(n10830) );
NAND2_X2 U6112 ( .A1(n13277), .A2(n15067), .ZN(n10835) );
NAND2_X2 U6114 ( .A1(n13358), .A2(n13056), .ZN(n10833) );
NAND2_X2 U6116 ( .A1(n13277), .A2(n15081), .ZN(n10838) );
NAND2_X2 U6118 ( .A1(n13358), .A2(n13055), .ZN(n10836) );
NAND2_X2 U6120 ( .A1(n13276), .A2(n15095), .ZN(n10841) );
NAND2_X2 U6122 ( .A1(n13358), .A2(n13054), .ZN(n10839) );
NAND2_X2 U6124 ( .A1(n13276), .A2(n15109), .ZN(n10844) );
NAND2_X2 U6126 ( .A1(n13357), .A2(n13053), .ZN(n10842) );
NAND2_X2 U6128 ( .A1(n13276), .A2(n15123), .ZN(n10847) );
NAND2_X2 U6130 ( .A1(n13357), .A2(n13052), .ZN(n10845) );
NAND2_X2 U6132 ( .A1(n13276), .A2(n15137), .ZN(n10850) );
NAND2_X2 U6134 ( .A1(n13357), .A2(n13051), .ZN(n10848) );
NAND2_X2 U6136 ( .A1(n13276), .A2(n15151), .ZN(n10853) );
NAND2_X2 U6138 ( .A1(n13357), .A2(n13050), .ZN(n10851) );
NAND2_X2 U6140 ( .A1(n13276), .A2(n15165), .ZN(n10856) );
NAND2_X2 U6142 ( .A1(n13357), .A2(n13049), .ZN(n10854) );
NAND2_X2 U6144 ( .A1(n13276), .A2(n15179), .ZN(n10859) );
NAND2_X2 U6146 ( .A1(n13357), .A2(n13048), .ZN(n10857) );
NAND2_X2 U6148 ( .A1(n13276), .A2(n15193), .ZN(n10862) );
NAND2_X2 U6150 ( .A1(n13357), .A2(n13047), .ZN(n10860) );
NAND2_X2 U6152 ( .A1(n13276), .A2(n15207), .ZN(n10865) );
NAND2_X2 U6154 ( .A1(n13357), .A2(n13046), .ZN(n10863) );
NAND2_X2 U6156 ( .A1(n13276), .A2(n15222), .ZN(n10868) );
NAND2_X2 U6158 ( .A1(n13357), .A2(n13045), .ZN(n10866) );
NAND2_X2 U6160 ( .A1(n13276), .A2(n15237), .ZN(n10871) );
NAND2_X2 U6162 ( .A1(n13357), .A2(n13044), .ZN(n10869) );
NAND2_X2 U6164 ( .A1(n13275), .A2(n15252), .ZN(n10874) );
NAND2_X2 U6166 ( .A1(n13357), .A2(n13043), .ZN(n10872) );
NAND2_X2 U6168 ( .A1(n13275), .A2(n15267), .ZN(n10877) );
NAND2_X2 U6170 ( .A1(n13356), .A2(n13042), .ZN(n10875) );
NAND2_X2 U6172 ( .A1(n13275), .A2(n15282), .ZN(n10880) );
NAND2_X2 U6174 ( .A1(n13356), .A2(n13041), .ZN(n10878) );
NAND2_X2 U6176 ( .A1(n13275), .A2(n15297), .ZN(n10883) );
NAND2_X2 U6178 ( .A1(n13356), .A2(n13040), .ZN(n10881) );
NAND2_X2 U6180 ( .A1(n13275), .A2(n15312), .ZN(n10886) );
NAND2_X2 U6182 ( .A1(n13356), .A2(n13039), .ZN(n10884) );
NAND2_X2 U6184 ( .A1(n13275), .A2(n15327), .ZN(n10889) );
NAND2_X2 U6186 ( .A1(n13356), .A2(n13038), .ZN(n10887) );
NAND2_X2 U6188 ( .A1(n13275), .A2(n15342), .ZN(n10892) );
NAND2_X2 U6190 ( .A1(n13356), .A2(n13037), .ZN(n10890) );
NAND2_X2 U6192 ( .A1(n13275), .A2(n15357), .ZN(n10895) );
NAND2_X2 U6194 ( .A1(n13356), .A2(n13036), .ZN(n10893) );
NAND2_X2 U6196 ( .A1(n13275), .A2(n15372), .ZN(n10898) );
NAND2_X2 U6198 ( .A1(n13356), .A2(n13035), .ZN(n10896) );
NAND2_X2 U6200 ( .A1(n13275), .A2(n15387), .ZN(n10901) );
NAND2_X2 U6202 ( .A1(n13356), .A2(n13034), .ZN(n10899) );
NAND2_X2 U6204 ( .A1(n13275), .A2(n15402), .ZN(n10904) );
NAND2_X2 U6206 ( .A1(n13356), .A2(n13033), .ZN(n10902) );
NAND2_X2 U6208 ( .A1(n13274), .A2(n15417), .ZN(n10907) );
NAND2_X2 U6212 ( .A1(n13356), .A2(n13032), .ZN(n10905) );
NAND2_X2 U6217 ( .A1(n13274), .A2(n14970), .ZN(n10910) );
NAND2_X2 U6218 ( .A1(n13353), .A2(n13063), .ZN(n10909) );
NAND2_X2 U6221 ( .A1(n13274), .A2(n14984), .ZN(n10915) );
NAND2_X2 U6222 ( .A1(n13353), .A2(n13062), .ZN(n10914) );
NAND2_X2 U6225 ( .A1(n13274), .A2(n14998), .ZN(n10918) );
NAND2_X2 U6226 ( .A1(n13353), .A2(n13061), .ZN(n10917) );
NAND2_X2 U6229 ( .A1(n13274), .A2(n15012), .ZN(n10921) );
NAND2_X2 U6230 ( .A1(n13353), .A2(n13060), .ZN(n10920) );
NAND2_X2 U6233 ( .A1(n13274), .A2(n15026), .ZN(n10924) );
NAND2_X2 U6234 ( .A1(n13353), .A2(n13059), .ZN(n10923) );
NAND2_X2 U6237 ( .A1(n13274), .A2(n15040), .ZN(n10927) );
NAND2_X2 U6238 ( .A1(n13353), .A2(n13058), .ZN(n10926) );
NAND2_X2 U6241 ( .A1(n13274), .A2(n15054), .ZN(n10930) );
NAND2_X2 U6242 ( .A1(n13353), .A2(n13057), .ZN(n10929) );
NAND2_X2 U6245 ( .A1(n13274), .A2(n15068), .ZN(n10933) );
NAND2_X2 U6246 ( .A1(n13353), .A2(n13056), .ZN(n10932) );
NAND2_X2 U6249 ( .A1(n13274), .A2(n15082), .ZN(n10936) );
NAND2_X2 U6250 ( .A1(n13353), .A2(n13055), .ZN(n10935) );
NAND2_X2 U6253 ( .A1(n13274), .A2(n15096), .ZN(n10939) );
NAND2_X2 U6254 ( .A1(n13353), .A2(n13054), .ZN(n10938) );
NAND2_X2 U6257 ( .A1(n13273), .A2(n15110), .ZN(n10942) );
NAND2_X2 U6258 ( .A1(n13353), .A2(n13053), .ZN(n10941) );
NAND2_X2 U6261 ( .A1(n13273), .A2(n15124), .ZN(n10945) );
NAND2_X2 U6262 ( .A1(n13354), .A2(n13052), .ZN(n10944) );
NAND2_X2 U6265 ( .A1(n13273), .A2(n15138), .ZN(n10948) );
NAND2_X2 U6266 ( .A1(n13354), .A2(n13051), .ZN(n10947) );
NAND2_X2 U6269 ( .A1(n13273), .A2(n15152), .ZN(n10951) );
NAND2_X2 U6270 ( .A1(n13354), .A2(n13050), .ZN(n10950) );
NAND2_X2 U6273 ( .A1(n13273), .A2(n15166), .ZN(n10954) );
NAND2_X2 U6274 ( .A1(n13354), .A2(n13049), .ZN(n10953) );
NAND2_X2 U6277 ( .A1(n13273), .A2(n15180), .ZN(n10957) );
NAND2_X2 U6278 ( .A1(n13354), .A2(n13048), .ZN(n10956) );
NAND2_X2 U6281 ( .A1(n13273), .A2(n15194), .ZN(n10960) );
NAND2_X2 U6282 ( .A1(n13354), .A2(n13047), .ZN(n10959) );
NAND2_X2 U6285 ( .A1(n13273), .A2(n15208), .ZN(n10963) );
NAND2_X2 U6286 ( .A1(n13354), .A2(n13046), .ZN(n10962) );
NAND2_X2 U6289 ( .A1(n13273), .A2(n15223), .ZN(n10966) );
NAND2_X2 U6290 ( .A1(n13354), .A2(n13045), .ZN(n10965) );
NAND2_X2 U6293 ( .A1(n13273), .A2(n15238), .ZN(n10969) );
NAND2_X2 U6294 ( .A1(n13354), .A2(n13044), .ZN(n10968) );
NAND2_X2 U6297 ( .A1(n13273), .A2(n15253), .ZN(n10972) );
NAND2_X2 U6298 ( .A1(n13354), .A2(n13043), .ZN(n10971) );
NAND2_X2 U6301 ( .A1(n13272), .A2(n15268), .ZN(n10975) );
NAND2_X2 U6302 ( .A1(n13354), .A2(n13042), .ZN(n10974) );
NAND2_X2 U6305 ( .A1(n13272), .A2(n15283), .ZN(n10978) );
NAND2_X2 U6306 ( .A1(n13355), .A2(n13041), .ZN(n10977) );
NAND2_X2 U6309 ( .A1(n13272), .A2(n15298), .ZN(n10981) );
NAND2_X2 U6310 ( .A1(n13355), .A2(n13040), .ZN(n10980) );
NAND2_X2 U6313 ( .A1(n13272), .A2(n15313), .ZN(n10984) );
NAND2_X2 U6314 ( .A1(n13355), .A2(n13039), .ZN(n10983) );
NAND2_X2 U6317 ( .A1(n13272), .A2(n15328), .ZN(n10987) );
NAND2_X2 U6318 ( .A1(n13355), .A2(n13038), .ZN(n10986) );
NAND2_X2 U6321 ( .A1(n13272), .A2(n15343), .ZN(n10990) );
NAND2_X2 U6322 ( .A1(n13355), .A2(n13037), .ZN(n10989) );
NAND2_X2 U6325 ( .A1(n13272), .A2(n15358), .ZN(n10993) );
NAND2_X2 U6326 ( .A1(n13355), .A2(n13036), .ZN(n10992) );
NAND2_X2 U6329 ( .A1(n13272), .A2(n15373), .ZN(n10996) );
NAND2_X2 U6330 ( .A1(n13355), .A2(n13035), .ZN(n10995) );
NAND2_X2 U6333 ( .A1(n13272), .A2(n15388), .ZN(n10999) );
NAND2_X2 U6334 ( .A1(n13355), .A2(n13034), .ZN(n10998) );
NAND2_X2 U6337 ( .A1(n13272), .A2(n15403), .ZN(n11002) );
NAND2_X2 U6338 ( .A1(n13355), .A2(n13033), .ZN(n11001) );
NAND2_X2 U6341 ( .A1(n13272), .A2(n15418), .ZN(n11005) );
NAND2_X2 U6343 ( .A1(n13355), .A2(n13032), .ZN(n11004) );
NAND2_X2 U7493 ( .A1(n11835), .A2(n11836), .ZN(n3696) );
NAND2_X2 U7495 ( .A1(read_counter[0]), .A2(n14954), .ZN(n11835) );
NAND2_X2 U7496 ( .A1(n11838), .A2(n11839), .ZN(n3695) );
NAND4_X2 U7503 ( .A1(n347), .A2(n11845), .A3(n11846), .A4(n14953), .ZN(n11837) );
NAND2_X2 U7505 ( .A1(n14955), .A2(n15425), .ZN(n11843) );
NAND4_X2 U7674 ( .A1(n11999), .A2(n12000), .A3(n12001), .A4(n12002), .ZN(n3672) );
NAND4_X2 U7682 ( .A1(n12006), .A2(n12007), .A3(n12008), .A4(n12009), .ZN(n3671) );
NAND4_X2 U7690 ( .A1(n12013), .A2(n12014), .A3(n12015), .A4(n12016), .ZN(n3670) );
NAND4_X2 U7698 ( .A1(n12020), .A2(n12021), .A3(n12022), .A4(n12023), .ZN(n3669) );
NAND4_X2 U7706 ( .A1(n12027), .A2(n12028), .A3(n12029), .A4(n12030), .ZN(n3668) );
NAND4_X2 U7714 ( .A1(n12034), .A2(n12035), .A3(n12036), .A4(n12037), .ZN(n3667) );
NAND4_X2 U7722 ( .A1(n12041), .A2(n12042), .A3(n12043), .A4(n12044), .ZN(n3666) );
NAND4_X2 U7730 ( .A1(n12048), .A2(n12049), .A3(n12050), .A4(n12051), .ZN(n3665) );
NAND4_X2 U7738 ( .A1(n12055), .A2(n12056), .A3(n12057), .A4(n12058), .ZN(n3664) );
NAND4_X2 U7746 ( .A1(n12062), .A2(n12063), .A3(n12064), .A4(n12065), .ZN(n3663) );
NAND4_X2 U7754 ( .A1(n12069), .A2(n12070), .A3(n12071), .A4(n12072), .ZN(n3662) );
NAND2_X2 U7760 ( .A1(read_counter[2]), .A2(n14956), .ZN(n11846) );
CLKBUFX1 gbuf_d_812(.A(N1717), .Y(d_out_812));
CLKBUFX1 gbuf_q_812(.A(q_in_812), .Y(round[3]));
CLKBUFX1 gbuf_qn_812(.A(qn_in_812), .Y(n14061));
CLKBUFX1 gbuf_d_813(.A(N1719), .Y(d_out_813));
CLKBUFX1 gbuf_q_813(.A(q_in_813), .Y(round[5]));
CLKBUFX1 gbuf_qn_813(.A(qn_in_813), .Y(n13973));
CLKBUFX1 gbuf_d_814(.A(n3990), .Y(d_out_814));
CLKBUFX1 gbuf_q_814(.A(q_in_814), .Y(n14394));
CLKBUFX1 gbuf_qn_814(.A(qn_in_814), .Y(n12903));
CLKBUFX1 gbuf_d_815(.A(n3992), .Y(d_out_815));
CLKBUFX1 gbuf_q_815(.A(q_in_815), .Y(n14400));
CLKBUFX1 gbuf_qn_815(.A(qn_in_815), .Y(n12899));
CLKBUFX1 gbuf_d_816(.A(n3991), .Y(d_out_816));
CLKBUFX1 gbuf_q_816(.A(q_in_816), .Y(n14397));
CLKBUFX1 gbuf_qn_816(.A(qn_in_816), .Y(n12901));
CLKBUFX1 gbuf_d_817(.A(n3995), .Y(d_out_817));
CLKBUFX1 gbuf_q_817(.A(q_in_817), .Y(n14408));
CLKBUFX1 gbuf_qn_817(.A(qn_in_817), .Y(n12893));
CLKBUFX1 gbuf_d_818(.A(N1716), .Y(d_out_818));
CLKBUFX1 gbuf_q_818(.A(q_in_818), .Y(n12988));
CLKBUFX1 gbuf_qn_818(.A(qn_in_818), .Y(n13116));
CLKBUFX1 gbuf_d_819(.A(N1715), .Y(d_out_819));
CLKBUFX1 gbuf_q_819(.A(q_in_819), .Y(round[1]));
CLKBUFX1 gbuf_qn_819(.A(qn_in_819), .Y(n14066));
CLKBUFX1 gbuf_d_820(.A(n3987), .Y(d_out_820));
CLKBUFX1 gbuf_q_820(.A(q_in_820), .Y(n14385));
CLKBUFX1 gbuf_qn_820(.A(qn_in_820), .Y(n12909));
CLKBUFX1 gbuf_d_821(.A(N1718), .Y(d_out_821));
CLKBUFX1 gbuf_q_821(.A(q_in_821), .Y(n12985));
CLKBUFX1 gbuf_qn_821(.A(qn_in_821), .Y(n13110));
CLKBUFX1 gbuf_d_822(.A(n3986), .Y(d_out_822));
CLKBUFX1 gbuf_q_822(.A(q_in_822), .Y(n14382));
CLKBUFX1 gbuf_qn_822(.A(qn_in_822), .Y(n12911));
CLKBUFX1 gbuf_d_823(.A(n3989), .Y(d_out_823));
CLKBUFX1 gbuf_q_823(.A(q_in_823), .Y(n14391));
CLKBUFX1 gbuf_qn_823(.A(qn_in_823), .Y(n12905));
CLKBUFX1 gbuf_d_824(.A(n3985), .Y(d_out_824));
CLKBUFX1 gbuf_q_824(.A(q_in_824), .Y(n14464));
CLKBUFX1 gbuf_qn_824(.A(qn_in_824), .Y(n12913));
CLKBUFX1 gbuf_d_825(.A(n3988), .Y(d_out_825));
CLKBUFX1 gbuf_q_825(.A(q_in_825), .Y(n14388));
CLKBUFX1 gbuf_qn_825(.A(qn_in_825), .Y(n12907));
CLKBUFX1 gbuf_d_826(.A(n3951), .Y(d_out_826));
CLKBUFX1 gbuf_q_826(.A(q_in_826), .Y(next_C[31]));
CLKBUFX1 gbuf_qn_826(.A(qn_in_826), .Y(n14743));
CLKBUFX1 gbuf_d_827(.A(n3947), .Y(d_out_827));
CLKBUFX1 gbuf_q_827(.A(q_in_827), .Y(next_C[3]));
CLKBUFX1 gbuf_qn_827(.A(qn_in_827), .Y(n13080));
CLKBUFX1 gbuf_d_828(.A(n4532), .Y(d_out_828));
CLKBUFX1 gbuf_q_828(.A(q_in_828), .Y(n14735));
CLKBUFX1 gbuf_qn_828(.A(qn_in_828), .Y(n8326));
CLKBUFX1 gbuf_d_829(.A(n13068), .Y(d_out_829));
CLKBUFX1 gbuf_q_829(.A(q_in_829), .Y(cmd_o[3]));
CLKBUFX1 gbuf_d_830(.A(n8328), .Y(d_out_830));
CLKBUFX1 gbuf_q_830(.A(q_in_830), .Y(Kt[28]));
CLKBUFX1 gbuf_d_831(.A(n14962), .Y(d_out_831));
CLKBUFX1 gbuf_q_831(.A(q_in_831), .Y(Kt[29]));
CLKBUFX1 gbuf_d_832(.A(n14962), .Y(d_out_832));
CLKBUFX1 gbuf_q_832(.A(q_in_832), .Y(Kt[9]));
CLKBUFX1 gbuf_d_833(.A(n14962), .Y(d_out_833));
CLKBUFX1 gbuf_q_833(.A(q_in_833), .Y(Kt[5]));
CLKBUFX1 gbuf_d_834(.A(N2583), .Y(d_out_834));
CLKBUFX1 gbuf_q_834(.A(q_in_834), .Y(Kt[23]));
CLKBUFX1 gbuf_d_835(.A(N2583), .Y(d_out_835));
CLKBUFX1 gbuf_q_835(.A(q_in_835), .Y(Kt[0]));
CLKBUFX1 gbuf_d_836(.A(n3696), .Y(d_out_836));
CLKBUFX1 gbuf_q_836(.A(q_in_836), .Y(read_counter[0]));
CLKBUFX1 gbuf_qn_836(.A(qn_in_836), .Y(n14952));
CLKBUFX1 gbuf_d_837(.A(n3695), .Y(d_out_837));
CLKBUFX1 gbuf_q_837(.A(q_in_837), .Y(read_counter[1]));
CLKBUFX1 gbuf_d_838(.A(n3694), .Y(d_out_838));
CLKBUFX1 gbuf_q_838(.A(q_in_838), .Y(read_counter[2]));
CLKBUFX1 gbuf_d_839(.A(n14932), .Y(d_out_839));
CLKBUFX1 gbuf_q_839(.A(q_in_839), .Y(Kt[21]));
CLKBUFX1 gbuf_d_840(.A(n14932), .Y(d_out_840));
CLKBUFX1 gbuf_q_840(.A(q_in_840), .Y(Kt[1]));
CLKBUFX1 gbuf_d_841(.A(N2595), .Y(d_out_841));
CLKBUFX1 gbuf_q_841(.A(q_in_841), .Y(Kt[22]));
CLKBUFX1 gbuf_d_842(.A(N2590), .Y(d_out_842));
CLKBUFX1 gbuf_q_842(.A(q_in_842), .Y(Kt[30]));
CLKBUFX1 gbuf_d_843(.A(N2590), .Y(d_out_843));
CLKBUFX1 gbuf_q_843(.A(q_in_843), .Y(Kt[14]));
CLKBUFX1 gbuf_d_844(.A(N2590), .Y(d_out_844));
CLKBUFX1 gbuf_q_844(.A(q_in_844), .Y(Kt[8]));
CLKBUFX1 gbuf_d_845(.A(n14931), .Y(d_out_845));
CLKBUFX1 gbuf_q_845(.A(q_in_845), .Y(Kt[24]));
CLKBUFX1 gbuf_d_846(.A(n14931), .Y(d_out_846));
CLKBUFX1 gbuf_q_846(.A(q_in_846), .Y(Kt[10]));
CLKBUFX1 gbuf_d_847(.A(n14961), .Y(d_out_847));
CLKBUFX1 gbuf_q_847(.A(q_in_847), .Y(Kt[12]));
CLKBUFX1 gbuf_d_848(.A(n14961), .Y(d_out_848));
CLKBUFX1 gbuf_q_848(.A(q_in_848), .Y(Kt[3]));
CLKBUFX1 gbuf_d_849(.A(N2589), .Y(d_out_849));
CLKBUFX1 gbuf_q_849(.A(q_in_849), .Y(Kt[27]));
CLKBUFX1 gbuf_d_850(.A(N2589), .Y(d_out_850));
CLKBUFX1 gbuf_q_850(.A(q_in_850), .Y(Kt[25]));
CLKBUFX1 gbuf_d_851(.A(N2589), .Y(d_out_851));
CLKBUFX1 gbuf_q_851(.A(q_in_851), .Y(Kt[7]));
CLKBUFX1 gbuf_d_852(.A(N2585), .Y(d_out_852));
CLKBUFX1 gbuf_q_852(.A(q_in_852), .Y(Kt[31]));
CLKBUFX1 gbuf_d_853(.A(N2585), .Y(d_out_853));
CLKBUFX1 gbuf_q_853(.A(q_in_853), .Y(Kt[6]));
CLKBUFX1 gbuf_d_854(.A(N2585), .Y(d_out_854));
CLKBUFX1 gbuf_q_854(.A(q_in_854), .Y(Kt[2]));
CLKBUFX1 gbuf_d_855(.A(n8330), .Y(d_out_855));
CLKBUFX1 gbuf_q_855(.A(q_in_855), .Y(Kt[26]));
CLKBUFX1 gbuf_d_856(.A(n8330), .Y(d_out_856));
CLKBUFX1 gbuf_q_856(.A(q_in_856), .Y(Kt[20]));
CLKBUFX1 gbuf_d_857(.A(n8330), .Y(d_out_857));
CLKBUFX1 gbuf_q_857(.A(q_in_857), .Y(Kt[19]));
CLKBUFX1 gbuf_d_858(.A(n8330), .Y(d_out_858));
CLKBUFX1 gbuf_q_858(.A(q_in_858), .Y(Kt[16]));
CLKBUFX1 gbuf_d_859(.A(n14960), .Y(d_out_859));
CLKBUFX1 gbuf_q_859(.A(q_in_859), .Y(Kt[15]));
CLKBUFX1 gbuf_d_860(.A(N2587), .Y(d_out_860));
CLKBUFX1 gbuf_q_860(.A(q_in_860), .Y(Kt[17]));
CLKBUFX1 gbuf_d_861(.A(N2587), .Y(d_out_861));
CLKBUFX1 gbuf_q_861(.A(q_in_861), .Y(Kt[4]));
CLKBUFX1 gbuf_d_862(.A(N2592), .Y(d_out_862));
CLKBUFX1 gbuf_q_862(.A(q_in_862), .Y(Kt[13]));
CLKBUFX1 gbuf_d_863(.A(N2592), .Y(d_out_863));
CLKBUFX1 gbuf_q_863(.A(q_in_863), .Y(Kt[11]));
CLKBUFX1 gbuf_d_864(.A(n3762), .Y(d_out_864));
CLKBUFX1 gbuf_q_864(.A(q_in_864), .Y(H4[30]));
CLKBUFX1 gbuf_d_865(.A(n3767), .Y(d_out_865));
CLKBUFX1 gbuf_q_865(.A(q_in_865), .Y(H4[25]));
CLKBUFX1 gbuf_d_866(.A(n3768), .Y(d_out_866));
CLKBUFX1 gbuf_q_866(.A(q_in_866), .Y(H4[24]));
CLKBUFX1 gbuf_d_867(.A(n3856), .Y(d_out_867));
CLKBUFX1 gbuf_q_867(.A(q_in_867), .Y(H3[0]));
CLKBUFX1 gbuf_d_868(.A(n3849), .Y(d_out_868));
CLKBUFX1 gbuf_q_868(.A(q_in_868), .Y(H3[7]));
CLKBUFX1 gbuf_d_869(.A(n3853), .Y(d_out_869));
CLKBUFX1 gbuf_q_869(.A(q_in_869), .Y(H3[3]));
CLKBUFX1 gbuf_d_870(.A(n3984), .Y(d_out_870));
CLKBUFX1 gbuf_q_870(.A(q_in_870), .Y(H0[0]));
CLKBUFX1 gbuf_d_871(.A(n3761), .Y(d_out_871));
CLKBUFX1 gbuf_q_871(.A(q_in_871), .Y(H4[31]));
CLKBUFX1 gbuf_d_872(.A(n3835), .Y(d_out_872));
CLKBUFX1 gbuf_q_872(.A(q_in_872), .Y(H3[21]));
CLKBUFX1 gbuf_d_873(.A(n3839), .Y(d_out_873));
CLKBUFX1 gbuf_q_873(.A(q_in_873), .Y(H3[17]));
CLKBUFX1 gbuf_d_874(.A(n3842), .Y(d_out_874));
CLKBUFX1 gbuf_q_874(.A(q_in_874), .Y(H3[14]));
CLKBUFX1 gbuf_d_875(.A(n3844), .Y(d_out_875));
CLKBUFX1 gbuf_q_875(.A(q_in_875), .Y(H3[12]));
CLKBUFX1 gbuf_d_876(.A(n3846), .Y(d_out_876));
CLKBUFX1 gbuf_q_876(.A(q_in_876), .Y(H3[10]));
CLKBUFX1 gbuf_d_877(.A(n3850), .Y(d_out_877));
CLKBUFX1 gbuf_q_877(.A(q_in_877), .Y(H3[6]));
CLKBUFX1 gbuf_d_878(.A(n3851), .Y(d_out_878));
CLKBUFX1 gbuf_q_878(.A(q_in_878), .Y(H3[5]));
CLKBUFX1 gbuf_d_879(.A(n3852), .Y(d_out_879));
CLKBUFX1 gbuf_q_879(.A(q_in_879), .Y(H3[4]));
CLKBUFX1 gbuf_d_880(.A(n3854), .Y(d_out_880));
CLKBUFX1 gbuf_q_880(.A(q_in_880), .Y(H3[2]));
CLKBUFX1 gbuf_d_881(.A(n3828), .Y(d_out_881));
CLKBUFX1 gbuf_q_881(.A(q_in_881), .Y(H3[28]));
CLKBUFX1 gbuf_d_882(.A(n3836), .Y(d_out_882));
CLKBUFX1 gbuf_q_882(.A(q_in_882), .Y(H3[20]));
CLKBUFX1 gbuf_d_883(.A(n3749), .Y(d_out_883));
CLKBUFX1 gbuf_q_883(.A(q_in_883), .Y(H2[11]));
CLKBUFX1 gbuf_d_884(.A(n3750), .Y(d_out_884));
CLKBUFX1 gbuf_q_884(.A(q_in_884), .Y(H2[10]));
CLKBUFX1 gbuf_d_885(.A(n3753), .Y(d_out_885));
CLKBUFX1 gbuf_q_885(.A(q_in_885), .Y(H2[7]));
CLKBUFX1 gbuf_d_886(.A(n3754), .Y(d_out_886));
CLKBUFX1 gbuf_q_886(.A(q_in_886), .Y(H2[6]));
CLKBUFX1 gbuf_d_887(.A(n3755), .Y(d_out_887));
CLKBUFX1 gbuf_q_887(.A(q_in_887), .Y(H2[5]));
CLKBUFX1 gbuf_d_888(.A(n3756), .Y(d_out_888));
CLKBUFX1 gbuf_q_888(.A(q_in_888), .Y(H2[4]));
CLKBUFX1 gbuf_d_889(.A(n3757), .Y(d_out_889));
CLKBUFX1 gbuf_q_889(.A(q_in_889), .Y(H2[3]));
CLKBUFX1 gbuf_d_890(.A(n3758), .Y(d_out_890));
CLKBUFX1 gbuf_q_890(.A(q_in_890), .Y(H2[2]));
CLKBUFX1 gbuf_d_891(.A(n3759), .Y(d_out_891));
CLKBUFX1 gbuf_q_891(.A(q_in_891), .Y(H2[1]));
CLKBUFX1 gbuf_d_892(.A(n3769), .Y(d_out_892));
CLKBUFX1 gbuf_q_892(.A(q_in_892), .Y(H4[23]));
CLKBUFX1 gbuf_d_893(.A(n13031), .Y(d_out_893));
CLKBUFX1 gbuf_q_893(.A(q_in_893), .Y(cmd_o[2]));
CLKBUFX1 gbuf_qn_893(.A(qn_in_893), .Y(n341));
CLKBUFX1 gbuf_d_894(.A(n3929), .Y(d_out_894));
CLKBUFX1 gbuf_q_894(.A(q_in_894), .Y(next_C[21]));
CLKBUFX1 gbuf_qn_894(.A(qn_in_894), .Y(n14680));
CLKBUFX1 gbuf_d_895(.A(n3879), .Y(d_out_895));
CLKBUFX1 gbuf_q_895(.A(q_in_895), .Y(n14797));
CLKBUFX1 gbuf_d_896(.A(n3919), .Y(d_out_896));
CLKBUFX1 gbuf_q_896(.A(q_in_896), .Y(SHA1_result[65]));
CLKBUFX1 gbuf_qn_896(.A(qn_in_896), .Y(n474));
CLKBUFX1 gbuf_d_897(.A(n4007), .Y(d_out_897));
CLKBUFX1 gbuf_q_897(.A(q_in_897), .Y(n14443));
CLKBUFX1 gbuf_qn_897(.A(qn_in_897), .Y(n12869));
CLKBUFX1 gbuf_d_898(.A(n4004), .Y(d_out_898));
CLKBUFX1 gbuf_q_898(.A(q_in_898), .Y(n14434));
CLKBUFX1 gbuf_qn_898(.A(qn_in_898), .Y(n12875));
CLKBUFX1 gbuf_d_899(.A(n4005), .Y(d_out_899));
CLKBUFX1 gbuf_q_899(.A(q_in_899), .Y(n14437));
CLKBUFX1 gbuf_qn_899(.A(qn_in_899), .Y(n12873));
CLKBUFX1 gbuf_d_900(.A(n4000), .Y(d_out_900));
CLKBUFX1 gbuf_q_900(.A(q_in_900), .Y(n14422));
CLKBUFX1 gbuf_qn_900(.A(qn_in_900), .Y(n12883));
CLKBUFX1 gbuf_d_901(.A(n3997), .Y(d_out_901));
CLKBUFX1 gbuf_q_901(.A(q_in_901), .Y(n14413));
CLKBUFX1 gbuf_qn_901(.A(qn_in_901), .Y(n12889));
CLKBUFX1 gbuf_d_902(.A(n4003), .Y(d_out_902));
CLKBUFX1 gbuf_q_902(.A(q_in_902), .Y(n14431));
CLKBUFX1 gbuf_qn_902(.A(qn_in_902), .Y(n12877));
CLKBUFX1 gbuf_d_903(.A(n4001), .Y(d_out_903));
CLKBUFX1 gbuf_q_903(.A(q_in_903), .Y(n14425));
CLKBUFX1 gbuf_qn_903(.A(qn_in_903), .Y(n12881));
CLKBUFX1 gbuf_d_904(.A(n4002), .Y(d_out_904));
CLKBUFX1 gbuf_q_904(.A(q_in_904), .Y(n14428));
CLKBUFX1 gbuf_qn_904(.A(qn_in_904), .Y(n12879));
CLKBUFX1 gbuf_d_905(.A(n3999), .Y(d_out_905));
CLKBUFX1 gbuf_q_905(.A(q_in_905), .Y(n14419));
CLKBUFX1 gbuf_qn_905(.A(qn_in_905), .Y(n12885));
CLKBUFX1 gbuf_d_906(.A(n3998), .Y(d_out_906));
CLKBUFX1 gbuf_q_906(.A(q_in_906), .Y(n14416));
CLKBUFX1 gbuf_qn_906(.A(qn_in_906), .Y(n12887));
CLKBUFX1 gbuf_d_907(.A(n3994), .Y(d_out_907));
CLKBUFX1 gbuf_q_907(.A(q_in_907), .Y(n14405));
CLKBUFX1 gbuf_qn_907(.A(qn_in_907), .Y(n12895));
CLKBUFX1 gbuf_d_908(.A(n3933), .Y(d_out_908));
CLKBUFX1 gbuf_q_908(.A(q_in_908), .Y(next_C[17]));
CLKBUFX1 gbuf_qn_908(.A(qn_in_908), .Y(n14861));
CLKBUFX1 gbuf_d_909(.A(n3949), .Y(d_out_909));
CLKBUFX1 gbuf_q_909(.A(q_in_909), .Y(next_C[1]));
CLKBUFX1 gbuf_qn_909(.A(qn_in_909), .Y(n14757));
CLKBUFX1 gbuf_d_910(.A(n3993), .Y(d_out_910));
CLKBUFX1 gbuf_q_910(.A(q_in_910), .Y(SHA1_result_151));
CLKBUFX1 gbuf_qn_910(.A(qn_in_910), .Y(n12897));
NAND3_X1 U8972 ( .A1(n14315), .A2(n14334), .A3(n13081), .ZN(n14316) );
INV_X2 U8973 ( .A(n14334), .ZN(n14360) );
INV_X4 U8974 ( .A(n14069), .ZN(n14350) );
NAND2_X2 U8975 ( .A1(next_C[12]), .A2(n13117), .ZN(n14218) );
INV_X16 U8976 ( .A(n13117), .ZN(n13163) );
NAND3_X2 U8977 ( .A1(n13591), .A2(n13590), .A3(n13589), .ZN(n3997) );
BUF_X32 U8978 ( .A(next_A[25]), .Z(n12982) );
NAND2_X1 U8979 ( .A1(n14330), .A2(n14312), .ZN(n14317) );
NAND3_X2 U8980 ( .A1(n13966), .A2(n13967), .A3(n14688), .ZN(n13078) );
INV_X4 U8981 ( .A(n13087), .ZN(n12980) );
NAND2_X2 U8982 ( .A1(n13146), .A2(n13971), .ZN(n14071) );
NAND2_X1 U8983 ( .A1(next_A[23]), .A2(n13207), .ZN(n13543) );
BUF_X32 U8984 ( .A(next_A[24]), .Z(n12981) );
BUF_X32 U8985 ( .A(next_A[30]), .Z(n12983) );
INV_X16 U8986 ( .A(n14174), .ZN(n13147) );
NAND3_X2 U8987 ( .A1(n14370), .A2(n13099), .A3(n13160), .ZN(n14374) );
NAND3_X2 U8988 ( .A1(n14372), .A2(n13084), .A3(n14371), .ZN(n14373) );
BUF_X32 U8989 ( .A(next_A[28]), .Z(n12984) );
NAND3_X4 U8990 ( .A1(n14327), .A2(n14328), .A3(n14329), .ZN(SHA1_ft_BCD[4]));
INV_X1 U8991 ( .A(n13092), .ZN(n14365) );
NOR2_X4 U8992 ( .A1(n474), .A2(n13092), .ZN(n14357) );
INV_X4 U8993 ( .A(n12985), .ZN(n12986) );
INV_X16 U8994 ( .A(n13113), .ZN(n14067) );
NOR3_X4 U8995 ( .A1(n14300), .A2(n14302), .A3(n14301), .ZN(n14303) );
NAND4_X4 U8996 ( .A1(n14303), .A2(n14306), .A3(n14304), .A4(n14305), .ZN(SHA1_ft_BCD[6]) );
MUX2_X2 U8997 ( .A(n14330), .B(n13142), .S(n13019), .Z(n14294) );
MUX2_X2 U8998 ( .A(n14331), .B(n13142), .S(n13015), .Z(n14326) );
NAND3_X1 U8999 ( .A1(n14332), .A2(SHA1_result[67]), .A3(n14331), .ZN(n14339));
INV_X8 U9000 ( .A(n13165), .ZN(n13162) );
NAND3_X4 U9001 ( .A1(n14234), .A2(n14233), .A3(n14232), .ZN(SHA1_ft_BCD[13]));
NAND2_X2 U9002 ( .A1(next_C[7]), .A2(n14342), .ZN(n14269) );
NAND3_X2 U9003 ( .A1(n14348), .A2(n13099), .A3(n14343), .ZN(n14347) );
NAND2_X1 U9004 ( .A1(next_C[6]), .A2(n14342), .ZN(n14280) );
NAND2_X1 U9005 ( .A1(next_C[2]), .A2(n14342), .ZN(n14322) );
INV_X1 U9006 ( .A(n14342), .ZN(n14343) );
INV_X8 U9007 ( .A(n13146), .ZN(n14065) );
NAND3_X2 U9008 ( .A1(n14220), .A2(SHA1_result[78]), .A3(n13163), .ZN(n14223));
INV_X4 U9009 ( .A(n13110), .ZN(n13146) );
NAND3_X2 U9010 ( .A1(n13542), .A2(n13543), .A3(n13541), .ZN(n3993) );
NAND2_X2 U9011 ( .A1(N875), .A2(n13212), .ZN(n13542) );
INV_X2 U9012 ( .A(n13116), .ZN(n13145) );
NAND2_X4 U9013 ( .A1(n14074), .A2(n13130), .ZN(n14198) );
INV_X8 U9014 ( .A(n14321), .ZN(n14330) );
INV_X16 U9015 ( .A(n14330), .ZN(n13117) );
AND2_X2 U9016 ( .A1(n14284), .A2(n14280), .ZN(n12987) );
NAND2_X4 U9017 ( .A1(n14266), .A2(n14071), .ZN(n14072) );
INV_X4 U9018 ( .A(n12988), .ZN(n12989) );
NAND3_X2 U9019 ( .A1(n13493), .A2(n13494), .A3(n13495), .ZN(n3989) );
NAND2_X2 U9020 ( .A1(N879), .A2(n13212), .ZN(n13493) );
INV_X16 U9021 ( .A(n13157), .ZN(n13160) );
NAND3_X2 U9022 ( .A1(n14198), .A2(n14273), .A3(n14350), .ZN(n14278) );
INV_X4 U9023 ( .A(n13098), .ZN(n13091) );
NOR3_X2 U9024 ( .A1(n437), .A2(next_C[4]), .A3(n13160), .ZN(n14300) );
NAND2_X2 U9025 ( .A1(n14186), .A2(n14185), .ZN(SHA1_ft_BCD[18]) );
INV_X4 U9026 ( .A(n14263), .ZN(n14255) );
INV_X4 U9027 ( .A(n13090), .ZN(n13097) );
NOR2_X2 U9028 ( .A1(n13147), .A2(n14258), .ZN(n14261) );
NOR3_X2 U9029 ( .A1(n14257), .A2(n433), .A3(n14256), .ZN(n14260) );
NOR3_X2 U9030 ( .A1(n14337), .A2(n14336), .A3(n14335), .ZN(n14338) );
NOR3_X2 U9031 ( .A1(n13160), .A2(next_C[1]), .A3(n440), .ZN(n14335) );
NOR3_X2 U9032 ( .A1(n14371), .A2(n14333), .A3(SHA1_result[67]), .ZN(n14337));
NAND4_X2 U9033 ( .A1(n14067), .A2(n14065), .A3(n13116), .A4(n14066), .ZN(n14068) );
NAND2_X2 U9034 ( .A1(n14349), .A2(n14309), .ZN(n14318) );
INV_X2 U9035 ( .A(n13147), .ZN(n13096) );
NAND2_X2 U9036 ( .A1(n14376), .A2(SHA1_result[32]), .ZN(n14377) );
INV_X4 U9037 ( .A(n442), .ZN(n14742) );
NAND3_X2 U9038 ( .A1(n13482), .A2(n13483), .A3(n13481), .ZN(n3988) );
NAND2_X2 U9039 ( .A1(N880), .A2(n13213), .ZN(n13482) );
NAND2_X1 U9040 ( .A1(next_C[31]), .A2(n13224), .ZN(n14533) );
NAND2_X1 U9041 ( .A1(n13197), .A2(next_C[31]), .ZN(n14529) );
NAND2_X1 U9042 ( .A1(n13200), .A2(next_C[31]), .ZN(n14599) );
INV_X16 U9043 ( .A(n13157), .ZN(n13161) );
INV_X16 U9044 ( .A(n13115), .ZN(n13157) );
OR2_X4 U9045 ( .A1(rst_i), .A2(n13805), .ZN(n12990) );
NAND3_X2 U9046 ( .A1(n13434), .A2(n13998), .A3(n12995), .ZN(n12991) );
NAND2_X2 U9047 ( .A1(n11114), .A2(cmd_o[2]), .ZN(n12992) );
AND2_X4 U9048 ( .A1(n11114), .A2(n341), .ZN(n12993) );
NAND2_X2 U9049 ( .A1(n13178), .A2(n13069), .ZN(n12994) );
AND2_X4 U9050 ( .A1(n13121), .A2(n14953), .ZN(n12995) );
NAND2_X2 U9051 ( .A1(n13438), .A2(n13437), .ZN(n12996) );
NAND3_X2 U9052 ( .A1(n13435), .A2(n14953), .A3(n13437), .ZN(n12997) );
AND2_X4 U9053 ( .A1(n13437), .A2(n14959), .ZN(n12998) );
AND2_X4 U9054 ( .A1(n14691), .A2(n13129), .ZN(n12999) );
NAND2_X1 U9055 ( .A1(n13178), .A2(n14688), .ZN(n14601) );
OR2_X4 U9056 ( .A1(n14732), .A2(n14731), .ZN(n13017) );
AND2_X4 U9057 ( .A1(n14691), .A2(n14953), .ZN(n13024) );
AND2_X4 U9058 ( .A1(n13129), .A2(n13398), .ZN(n13025) );
AND4_X4 U9059 ( .A1(n14699), .A2(n14719), .A3(n14729), .A4(n13401), .ZN(n13026) );
AND2_X4 U9060 ( .A1(n14726), .A2(n13413), .ZN(n13027) );
AND2_X4 U9061 ( .A1(n14704), .A2(n14953), .ZN(n13028) );
AND2_X4 U9062 ( .A1(n14002), .A2(n14953), .ZN(n13029) );
NAND3_X4 U9063 ( .A1(n13614), .A2(n13615), .A3(n13613), .ZN(n3999) );
NAND2_X4 U9064 ( .A1(N869), .A2(n13211), .ZN(n13614) );
NAND2_X1 U9065 ( .A1(n9301), .A2(cmd_o[3]), .ZN(n9308) );
INV_X1 U9066 ( .A(n13030), .ZN(n13031) );
INV_X32 U9067 ( .A(n4533), .ZN(n13030) );
NAND2_X1 U9068 ( .A1(n9299), .A2(n9300), .ZN(n4533) );
NAND2_X1 U9069 ( .A1(cmd_i[2]), .A2(n9301), .ZN(n9299) );
CLKBUF_X2 U9070 ( .A(text_i[31]), .Z(n13032) );
NAND2_X1 U9071 ( .A1(n13032), .A2(n13320), .ZN(n9509) );
CLKBUF_X2 U9072 ( .A(text_i[30]), .Z(n13033) );
NAND2_X1 U9073 ( .A1(n13033), .A2(n13320), .ZN(n9503) );
CLKBUF_X2 U9074 ( .A(text_i[29]), .Z(n13034) );
NAND2_X1 U9075 ( .A1(n13034), .A2(n13320), .ZN(n9497) );
CLKBUF_X2 U9076 ( .A(text_i[28]), .Z(n13035) );
NAND2_X1 U9077 ( .A1(n13035), .A2(n13320), .ZN(n9491) );
CLKBUF_X2 U9078 ( .A(text_i[27]), .Z(n13036) );
NAND2_X1 U9079 ( .A1(n13036), .A2(n13320), .ZN(n9485) );
CLKBUF_X2 U9080 ( .A(text_i[26]), .Z(n13037) );
NAND2_X1 U9081 ( .A1(n13037), .A2(n13320), .ZN(n9479) );
CLKBUF_X2 U9082 ( .A(text_i[25]), .Z(n13038) );
NAND2_X1 U9083 ( .A1(n13038), .A2(n13320), .ZN(n9473) );
CLKBUF_X2 U9084 ( .A(text_i[24]), .Z(n13039) );
NAND2_X1 U9085 ( .A1(n13039), .A2(n13320), .ZN(n9467) );
CLKBUF_X2 U9086 ( .A(text_i[23]), .Z(n13040) );
NAND2_X1 U9087 ( .A1(n13040), .A2(n13320), .ZN(n9461) );
CLKBUF_X2 U9088 ( .A(text_i[22]), .Z(n13041) );
NAND2_X1 U9089 ( .A1(n13041), .A2(n13320), .ZN(n9455) );
CLKBUF_X2 U9090 ( .A(text_i[21]), .Z(n13042) );
NAND2_X1 U9091 ( .A1(n13042), .A2(n13319), .ZN(n9449) );
CLKBUF_X2 U9092 ( .A(text_i[20]), .Z(n13043) );
NAND2_X1 U9093 ( .A1(n13043), .A2(n13319), .ZN(n9443) );
CLKBUF_X2 U9094 ( .A(text_i[19]), .Z(n13044) );
NAND2_X1 U9095 ( .A1(n13044), .A2(n13319), .ZN(n9437) );
CLKBUF_X2 U9096 ( .A(text_i[18]), .Z(n13045) );
NAND2_X1 U9097 ( .A1(n13045), .A2(n13319), .ZN(n9431) );
CLKBUF_X2 U9098 ( .A(text_i[17]), .Z(n13046) );
NAND2_X1 U9099 ( .A1(n13318), .A2(n13046), .ZN(n14005) );
CLKBUF_X2 U9100 ( .A(text_i[16]), .Z(n13047) );
NAND2_X1 U9101 ( .A1(n13318), .A2(n13047), .ZN(n14008) );
CLKBUF_X2 U9102 ( .A(text_i[15]), .Z(n13048) );
NAND2_X1 U9103 ( .A1(n13318), .A2(n13048), .ZN(n14011) );
CLKBUF_X2 U9104 ( .A(text_i[14]), .Z(n13049) );
NAND2_X1 U9105 ( .A1(n13318), .A2(n13049), .ZN(n14014) );
CLKBUF_X2 U9106 ( .A(text_i[13]), .Z(n13050) );
NAND2_X1 U9107 ( .A1(n13318), .A2(n13050), .ZN(n14017) );
CLKBUF_X2 U9108 ( .A(text_i[12]), .Z(n13051) );
NAND2_X1 U9109 ( .A1(n13318), .A2(n13051), .ZN(n14020) );
CLKBUF_X2 U9110 ( .A(text_i[11]), .Z(n13052) );
NAND2_X1 U9111 ( .A1(n13318), .A2(n13052), .ZN(n14023) );
CLKBUF_X2 U9112 ( .A(text_i[10]), .Z(n13053) );
NAND2_X1 U9113 ( .A1(n13318), .A2(n13053), .ZN(n14026) );
CLKBUF_X2 U9114 ( .A(text_i[9]), .Z(n13054) );
NAND2_X1 U9115 ( .A1(n13318), .A2(n13054), .ZN(n14029) );
CLKBUF_X2 U9116 ( .A(text_i[8]), .Z(n13055) );
NAND2_X1 U9117 ( .A1(n13318), .A2(n13055), .ZN(n14032) );
CLKBUF_X2 U9118 ( .A(text_i[7]), .Z(n13056) );
NAND2_X1 U9119 ( .A1(n13318), .A2(n13056), .ZN(n14035) );
CLKBUF_X2 U9120 ( .A(text_i[6]), .Z(n13057) );
NAND2_X1 U9121 ( .A1(n13319), .A2(n13057), .ZN(n14038) );
CLKBUF_X2 U9122 ( .A(text_i[5]), .Z(n13058) );
NAND2_X1 U9123 ( .A1(n13319), .A2(n13058), .ZN(n14041) );
CLKBUF_X2 U9124 ( .A(text_i[4]), .Z(n13059) );
NAND2_X1 U9125 ( .A1(n13319), .A2(n13059), .ZN(n14044) );
CLKBUF_X2 U9126 ( .A(text_i[3]), .Z(n13060) );
NAND2_X1 U9127 ( .A1(n13319), .A2(n13060), .ZN(n14047) );
CLKBUF_X2 U9128 ( .A(text_i[2]), .Z(n13061) );
NAND2_X1 U9129 ( .A1(n13319), .A2(n13061), .ZN(n14050) );
CLKBUF_X2 U9130 ( .A(text_i[1]), .Z(n13062) );
NAND2_X1 U9131 ( .A1(n13319), .A2(n13062), .ZN(n14053) );
CLKBUF_X2 U9132 ( .A(text_i[0]), .Z(n13063) );
NAND2_X1 U9133 ( .A1(n13063), .A2(n13392), .ZN(n9315) );
INV_X1 U9134 ( .A(n13064), .ZN(n13065) );
INV_X32 U9135 ( .A(n4530), .ZN(n13064) );
NAND2_X1 U9136 ( .A1(n9310), .A2(n9311), .ZN(n4530) );
NAND2_X1 U9137 ( .A1(cmd_i[0]), .A2(n9301), .ZN(n9310) );
INV_X1 U9138 ( .A(n13066), .ZN(n13067) );
INV_X32 U9139 ( .A(n4529), .ZN(n13066) );
NAND2_X1 U9140 ( .A1(n9313), .A2(n9314), .ZN(n4529) );
NAND2_X1 U9141 ( .A1(cmd_i[1]), .A2(n9301), .ZN(n9313) );
BUF_X8 U9142 ( .A(n4531), .Z(n13068) );
NAND2_X1 U9143 ( .A1(n14958), .A2(n9308), .ZN(n4531) );
NOR3_X1 U9144 ( .A1(n8326), .A2(rst_i), .A3(cmd_w_i), .ZN(n9309) );
NAND4_X2 U9145 ( .A1(n13529), .A2(n13530), .A3(n14601), .A4(n13531), .ZN(n3992) );
NAND2_X2 U9146 ( .A1(N878), .A2(n13178), .ZN(n13505) );
NAND4_X2 U9147 ( .A1(n13505), .A2(n13507), .A3(n14601), .A4(n13506), .ZN(n3990) );
NOR2_X2 U9148 ( .A1(n13097), .A2(n13163), .ZN(n14254) );
NAND3_X1 U9149 ( .A1(n465), .A2(n14368), .A3(n14263), .ZN(n14264) );
NAND2_X1 U9150 ( .A1(n13968), .A2(n14688), .ZN(n13970) );
NAND2_X1 U9151 ( .A1(n13069), .A2(n12986), .ZN(n13429) );
INV_X1 U9152 ( .A(n14071), .ZN(n13070) );
INV_X4 U9153 ( .A(n13070), .ZN(n13071) );
INV_X2 U9154 ( .A(n14350), .ZN(n13072) );
INV_X4 U9155 ( .A(n13072), .ZN(n13073) );
INV_X16 U9156 ( .A(n13160), .ZN(n13158) );
INV_X8 U9157 ( .A(n13160), .ZN(n13159) );
NOR3_X2 U9158 ( .A1(n13161), .A2(n442), .A3(next_C[31]), .ZN(n14362) );
INV_X1 U9159 ( .A(n14368), .ZN(n13074) );
INV_X8 U9160 ( .A(n14064), .ZN(n14213) );
NAND2_X4 U9161 ( .A1(n14198), .A2(n14273), .ZN(n14064) );
NAND2_X4 U9162 ( .A1(round[3]), .A2(n13077), .ZN(n13966) );
INV_X2 U9163 ( .A(n14351), .ZN(n13099) );
NAND2_X2 U9164 ( .A1(n14266), .A2(n14071), .ZN(n13075) );
INV_X4 U9165 ( .A(next_A[16]), .ZN(n13107) );
INV_X8 U9166 ( .A(n13077), .ZN(n13076) );
INV_X4 U9167 ( .A(n13973), .ZN(n13077) );
NAND2_X2 U9168 ( .A1(n13103), .A2(n14198), .ZN(n14369) );
NAND2_X1 U9169 ( .A1(next_A[12]), .A2(n13206), .ZN(n13675) );
NAND3_X2 U9170 ( .A1(n14297), .A2(n14296), .A3(n14295), .ZN(SHA1_ft_BCD[7]));
INV_X8 U9171 ( .A(n14356), .ZN(n14349) );
MUX2_X2 U9172 ( .A(n14351), .B(n13142), .S(n13079), .Z(n14274) );
INV_X4 U9173 ( .A(n13080), .ZN(n13081) );
INV_X4 U9174 ( .A(n14369), .ZN(n14351) );
NAND3_X4 U9175 ( .A1(n14353), .A2(n14354), .A3(n14355), .ZN(SHA1_ft_BCD[2]));
NAND2_X4 U9176 ( .A1(n14352), .A2(SHA1_result[34]), .ZN(n14353) );
INV_X1 U9177 ( .A(n13142), .ZN(n13082) );
BUF_X4 U9178 ( .A(n14375), .Z(n13142) );
NAND2_X2 U9179 ( .A1(n14279), .A2(n14267), .ZN(n14356) );
INV_X8 U9180 ( .A(n13143), .ZN(n14331) );
MUX2_X2 U9181 ( .A(n14351), .B(n13142), .S(n13083), .Z(n14352) );
NAND2_X4 U9182 ( .A1(n14279), .A2(n14278), .ZN(n14344) );
MUX2_X2 U9183 ( .A(n14351), .B(n13142), .S(n13084), .Z(n14376) );
AND3_X4 U9184 ( .A1(n13114), .A2(n13973), .A3(n14061), .ZN(n14060) );
NAND3_X2 U9185 ( .A1(n14197), .A2(n14196), .A3(n14195), .ZN(SHA1_ft_BCD[17]));
BUF_X32 U9186 ( .A(next_A[18]), .Z(n13085) );
NAND2_X1 U9187 ( .A1(n13085), .A2(n13207), .ZN(n13601) );
NAND2_X1 U9188 ( .A1(next_A[7]), .A2(n13206), .ZN(n13735) );
NAND2_X1 U9189 ( .A1(next_A[9]), .A2(n13206), .ZN(n13709) );
NOR2_X1 U9190 ( .A1(n13411), .A2(n12989), .ZN(n13412) );
INV_X1 U9191 ( .A(round[3]), .ZN(n13086) );
INV_X4 U9192 ( .A(n13086), .ZN(n13087) );
NAND3_X2 U9193 ( .A1(n14060), .A2(n14066), .A3(n14067), .ZN(n13088) );
INV_X4 U9194 ( .A(n13107), .ZN(n13108) );
BUF_X32 U9195 ( .A(next_A[14]), .Z(n13089) );
NAND3_X1 U9196 ( .A1(n12999), .A2(n13069), .A3(n13076), .ZN(n13426) );
NAND2_X4 U9197 ( .A1(n13091), .A2(n13157), .ZN(n13090) );
XNOR2_X2 U9198 ( .A(next_C[31]), .B(n14742), .ZN(n13092) );
INV_X4 U9199 ( .A(round[1]), .ZN(n13093) );
NOR2_X1 U9200 ( .A1(n14065), .A2(n14061), .ZN(n13130) );
BUF_X32 U9201 ( .A(next_A[21]), .Z(n13094) );
NAND2_X1 U9202 ( .A1(n12982), .A2(n13208), .ZN(n13517) );
BUF_X32 U9203 ( .A(next_A[13]), .Z(n13095) );
NAND4_X4 U9204 ( .A1(n14225), .A2(n14224), .A3(n14223), .A4(n14222), .ZN(SHA1_ft_BCD[14]) );
BUF_X32 U9205 ( .A(next_A[20]), .Z(n13106) );
NAND2_X2 U9206 ( .A1(n14169), .A2(n14168), .ZN(SHA1_ft_BCD[20]) );
NOR2_X1 U9207 ( .A1(n13076), .A2(n13419), .ZN(n13415) );
NAND2_X1 U9208 ( .A1(n13076), .A2(n12986), .ZN(n13402) );
NAND2_X4 U9209 ( .A1(n14068), .A2(n14688), .ZN(n14069) );
BUF_X32 U9210 ( .A(next_A[17]), .Z(n13100) );
INV_X4 U9211 ( .A(n13974), .ZN(n13101) );
INV_X4 U9212 ( .A(n13114), .ZN(n13144) );
NAND3_X2 U9213 ( .A1(n14060), .A2(n14066), .A3(n14067), .ZN(n13102) );
AND2_X2 U9214 ( .A1(n13078), .A2(n14350), .ZN(n13103) );
NAND2_X4 U9215 ( .A1(n14213), .A2(n13073), .ZN(n13143) );
NAND3_X1 U9216 ( .A1(n14322), .A2(n14344), .A3(n14320), .ZN(n14325) );
BUF_X32 U9217 ( .A(next_A[27]), .Z(n13104) );
NAND3_X1 U9218 ( .A1(next_C[12]), .A2(n13158), .A3(SHA1_result[78]), .ZN(n14224) );
NAND2_X1 U9219 ( .A1(next_C[15]), .A2(n13158), .ZN(n14191) );
NOR4_X4 U9220 ( .A1(n14262), .A2(n14261), .A3(n14260), .A4(n14259), .ZN(n14265) );
NAND2_X1 U9221 ( .A1(n13207), .A2(n13089), .ZN(n13651) );
NAND2_X1 U9222 ( .A1(n13222), .A2(n14391), .ZN(n13494) );
INV_X8 U9223 ( .A(n14073), .ZN(n14279) );
BUF_X32 U9224 ( .A(next_A[19]), .Z(n13105) );
NAND2_X1 U9225 ( .A1(n13105), .A2(n13207), .ZN(n13591) );
NAND2_X4 U9226 ( .A1(n14072), .A2(n13088), .ZN(n14375) );
NAND2_X4 U9227 ( .A1(n13102), .A2(n14072), .ZN(n14073) );
BUF_X32 U9228 ( .A(next_A[15]), .Z(n13109) );
BUF_X32 U9229 ( .A(next_A[10]), .Z(n13111) );
NAND2_X1 U9230 ( .A1(n13207), .A2(n13109), .ZN(n13639) );
INV_X4 U9231 ( .A(n13112), .ZN(n13113) );
NAND3_X1 U9232 ( .A1(n14281), .A2(n14371), .A3(n14280), .ZN(n14282) );
NAND2_X1 U9233 ( .A1(n12984), .A2(n13208), .ZN(n13483) );
INV_X8 U9234 ( .A(n13165), .ZN(n13164) );
INV_X8 U9235 ( .A(n14331), .ZN(n13165) );
NAND2_X1 U9236 ( .A1(n14174), .A2(n14165), .ZN(n14166) );
NAND2_X1 U9237 ( .A1(n14174), .A2(n14157), .ZN(n14158) );
NAND2_X1 U9238 ( .A1(n14174), .A2(n14149), .ZN(n14150) );
NAND2_X1 U9239 ( .A1(n14174), .A2(n14173), .ZN(n14175) );
NAND3_X2 U9240 ( .A1(n474), .A2(n14365), .A3(n14368), .ZN(n14366) );
NAND3_X2 U9241 ( .A1(n14198), .A2(n13078), .A3(n14350), .ZN(n14267) );
NAND4_X4 U9242 ( .A1(n14319), .A2(n14318), .A3(n14317), .A4(n14316), .ZN(n14930) );
NAND3_X1 U9243 ( .A1(round[0]), .A2(n13398), .A3(n13093), .ZN(n14693) );
NAND2_X1 U9244 ( .A1(n13104), .A2(n13208), .ZN(n13495) );
NAND2_X1 U9245 ( .A1(n13111), .A2(n13206), .ZN(n13699) );
NAND2_X1 U9246 ( .A1(n12981), .A2(n13207), .ZN(n13531) );
NAND2_X1 U9247 ( .A1(n13100), .A2(n13207), .ZN(n13615) );
INV_X4 U9248 ( .A(n14375), .ZN(n13115) );
NAND2_X1 U9249 ( .A1(n13095), .A2(n13207), .ZN(n13661) );
NAND2_X4 U9250 ( .A1(n13145), .A2(n14062), .ZN(n14063) );
NAND2_X4 U9251 ( .A1(n14067), .A2(n14066), .ZN(n14062) );
NAND2_X2 U9252 ( .A1(n13077), .A2(n13146), .ZN(n13967) );
INV_X16 U9253 ( .A(n14371), .ZN(n14174) );
NAND2_X4 U9254 ( .A1(n14213), .A2(n13073), .ZN(n14321) );
NAND2_X1 U9255 ( .A1(next_A[29]), .A2(n13208), .ZN(n13471) );
NAND2_X2 U9256 ( .A1(n12987), .A2(n13117), .ZN(n14283) );
NOR2_X1 U9257 ( .A1(n13082), .A2(n13014), .ZN(n14100) );
NOR2_X1 U9258 ( .A1(n13082), .A2(n13007), .ZN(n14084) );
NOR2_X1 U9259 ( .A1(n13082), .A2(n13013), .ZN(n14092) );
NOR2_X1 U9260 ( .A1(n13082), .A2(n13002), .ZN(n14076) );
NAND3_X1 U9261 ( .A1(cmd_o[1]), .A2(n12999), .A3(n14688), .ZN(n14689) );
NAND3_X1 U9262 ( .A1(n13101), .A2(n14953), .A3(n13969), .ZN(n13983) );
INV_X1 U9263 ( .A(n13078), .ZN(n13974) );
INV_X4 U9264 ( .A(n13182), .ZN(n13184) );
INV_X4 U9265 ( .A(n13182), .ZN(n13183) );
INV_X4 U9266 ( .A(n12991), .ZN(n13206) );
INV_X4 U9267 ( .A(n13430), .ZN(n13179) );
INV_X4 U9268 ( .A(n13430), .ZN(n13180) );
INV_X4 U9269 ( .A(n12991), .ZN(n13204) );
INV_X4 U9270 ( .A(n12991), .ZN(n13202) );
INV_X4 U9271 ( .A(n12991), .ZN(n13201) );
INV_X4 U9272 ( .A(n12991), .ZN(n13200) );
INV_X4 U9273 ( .A(n12991), .ZN(n13205) );
INV_X4 U9274 ( .A(n12991), .ZN(n13207) );
INV_X4 U9275 ( .A(n12991), .ZN(n13203) );
INV_X4 U9276 ( .A(n13430), .ZN(n13181) );
INV_X4 U9277 ( .A(n12994), .ZN(n13212) );
INV_X4 U9278 ( .A(n12994), .ZN(n13211) );
INV_X4 U9279 ( .A(n12994), .ZN(n13210) );
INV_X4 U9280 ( .A(n12994), .ZN(n13209) );
INV_X4 U9281 ( .A(n13182), .ZN(n13185) );
INV_X4 U9282 ( .A(n12994), .ZN(n13213) );
INV_X4 U9283 ( .A(n12991), .ZN(n13208) );
INV_X4 U9284 ( .A(n14701), .ZN(n13235) );
INV_X4 U9285 ( .A(n14702), .ZN(n13238) );
INV_X4 U9286 ( .A(n14703), .ZN(n13241) );
INV_X4 U9287 ( .A(n14709), .ZN(n13262) );
INV_X4 U9288 ( .A(n14710), .ZN(n13247) );
INV_X4 U9289 ( .A(n14711), .ZN(n13250) );
INV_X4 U9290 ( .A(n14720), .ZN(n13256) );
INV_X4 U9291 ( .A(n14710), .ZN(n13246) );
INV_X4 U9292 ( .A(n14711), .ZN(n13249) );
INV_X4 U9293 ( .A(n14720), .ZN(n13255) );
INV_X4 U9294 ( .A(n14701), .ZN(n13234) );
INV_X4 U9295 ( .A(n14702), .ZN(n13237) );
INV_X4 U9296 ( .A(n14703), .ZN(n13240) );
INV_X4 U9297 ( .A(n14709), .ZN(n13261) );
INV_X4 U9298 ( .A(n14701), .ZN(n13236) );
INV_X4 U9299 ( .A(n14702), .ZN(n13239) );
INV_X4 U9300 ( .A(n14703), .ZN(n13242) );
INV_X4 U9301 ( .A(n14709), .ZN(n13263) );
INV_X4 U9302 ( .A(n14710), .ZN(n13248) );
INV_X4 U9303 ( .A(n14711), .ZN(n13251) );
INV_X4 U9304 ( .A(n14720), .ZN(n13257) );
INV_X4 U9305 ( .A(n12992), .ZN(n13199) );
INV_X4 U9306 ( .A(n12992), .ZN(n13198) );
INV_X4 U9307 ( .A(n12992), .ZN(n13195) );
INV_X4 U9308 ( .A(n12992), .ZN(n13196) );
INV_X4 U9309 ( .A(n12996), .ZN(n13172) );
INV_X4 U9310 ( .A(n12992), .ZN(n13197) );
INV_X4 U9311 ( .A(n12992), .ZN(n13193) );
INV_X4 U9312 ( .A(n12992), .ZN(n13194) );
INV_X4 U9313 ( .A(n13121), .ZN(n13222) );
INV_X4 U9314 ( .A(n13121), .ZN(n13223) );
INV_X4 U9315 ( .A(n13430), .ZN(n13178) );
INV_X4 U9316 ( .A(n13119), .ZN(n13231) );
INV_X4 U9317 ( .A(n13119), .ZN(n13232) );
INV_X4 U9318 ( .A(n13119), .ZN(n13233) );
INV_X4 U9319 ( .A(n13120), .ZN(n13333) );
INV_X4 U9320 ( .A(n13120), .ZN(n13334) );
INV_X4 U9321 ( .A(n13118), .ZN(n13354) );
INV_X4 U9322 ( .A(n13118), .ZN(n13353) );
INV_X4 U9323 ( .A(n13120), .ZN(n13335) );
INV_X4 U9324 ( .A(n13118), .ZN(n13355) );
INV_X4 U9325 ( .A(n14698), .ZN(n13362) );
INV_X4 U9326 ( .A(n14706), .ZN(n13374) );
INV_X4 U9327 ( .A(n14713), .ZN(n13383) );
INV_X4 U9328 ( .A(n14692), .ZN(n13356) );
INV_X4 U9329 ( .A(n14696), .ZN(n13359) );
INV_X4 U9330 ( .A(n14692), .ZN(n13357) );
INV_X4 U9331 ( .A(n14696), .ZN(n13360) );
INV_X4 U9332 ( .A(n14698), .ZN(n13363) );
INV_X4 U9333 ( .A(n14706), .ZN(n13375) );
INV_X4 U9334 ( .A(n14713), .ZN(n13384) );
INV_X4 U9335 ( .A(n14725), .ZN(n13259) );
INV_X4 U9336 ( .A(n14725), .ZN(n13258) );
INV_X4 U9337 ( .A(n14713), .ZN(n13385) );
INV_X4 U9338 ( .A(n14692), .ZN(n13358) );
INV_X4 U9339 ( .A(n14696), .ZN(n13361) );
INV_X4 U9340 ( .A(n14698), .ZN(n13364) );
INV_X4 U9341 ( .A(n14706), .ZN(n13376) );
INV_X4 U9342 ( .A(n12998), .ZN(n13149) );
INV_X4 U9343 ( .A(n14725), .ZN(n13260) );
INV_X4 U9344 ( .A(n12996), .ZN(n13175) );
INV_X4 U9345 ( .A(n12996), .ZN(n13176) );
INV_X4 U9346 ( .A(n12996), .ZN(n13173) );
INV_X4 U9347 ( .A(n12996), .ZN(n13174) );
INV_X4 U9348 ( .A(n13121), .ZN(n13215) );
INV_X4 U9349 ( .A(n13121), .ZN(n13221) );
INV_X4 U9350 ( .A(n13121), .ZN(n13220) );
INV_X4 U9351 ( .A(n13121), .ZN(n13219) );
INV_X4 U9352 ( .A(n13121), .ZN(n13218) );
INV_X4 U9353 ( .A(n13121), .ZN(n13217) );
INV_X4 U9354 ( .A(n13121), .ZN(n13216) );
INV_X4 U9355 ( .A(n13121), .ZN(n13214) );
INV_X4 U9356 ( .A(n12998), .ZN(n13148) );
INV_X4 U9357 ( .A(n12997), .ZN(n13169) );
INV_X4 U9358 ( .A(n12997), .ZN(n13170) );
INV_X4 U9359 ( .A(n12997), .ZN(n13167) );
INV_X4 U9360 ( .A(n12997), .ZN(n13168) );
INV_X4 U9361 ( .A(n12997), .ZN(n13166) );
INV_X4 U9362 ( .A(n13121), .ZN(n13224) );
INV_X4 U9363 ( .A(n12996), .ZN(n13177) );
INV_X4 U9364 ( .A(n12997), .ZN(n13171) );
INV_X4 U9365 ( .A(n12998), .ZN(n13150) );
INV_X4 U9366 ( .A(n12990), .ZN(n13321) );
INV_X4 U9367 ( .A(n14601), .ZN(n13182) );
INV_X4 U9368 ( .A(n14000), .ZN(n13156) );
INV_X4 U9369 ( .A(n12993), .ZN(n13192) );
INV_X4 U9370 ( .A(n12993), .ZN(n13188) );
INV_X4 U9371 ( .A(n12993), .ZN(n13189) );
INV_X4 U9372 ( .A(n12993), .ZN(n13191) );
INV_X4 U9373 ( .A(n12993), .ZN(n13190) );
INV_X4 U9374 ( .A(n12993), .ZN(n13187) );
INV_X4 U9375 ( .A(n12993), .ZN(n13186) );
OR2_X2 U9376 ( .A1(n14959), .A2(n13270), .ZN(n13118) );
BUF_X4 U9377 ( .A(n13029), .Z(n13316) );
BUF_X4 U9378 ( .A(n13029), .Z(n13272) );
BUF_X4 U9379 ( .A(n13029), .Z(n13301) );
BUF_X4 U9380 ( .A(n13029), .Z(n13275) );
BUF_X4 U9381 ( .A(n13029), .Z(n13304) );
BUF_X4 U9382 ( .A(n13029), .Z(n13314) );
BUF_X4 U9383 ( .A(n13029), .Z(n13278) );
BUF_X4 U9384 ( .A(n13029), .Z(n13307) );
BUF_X4 U9385 ( .A(n13029), .Z(n13281) );
BUF_X4 U9386 ( .A(n13029), .Z(n13310) );
BUF_X4 U9387 ( .A(n13029), .Z(n13313) );
BUF_X4 U9388 ( .A(n13029), .Z(n13284) );
BUF_X4 U9389 ( .A(n13029), .Z(n13287) );
BUF_X4 U9390 ( .A(n13029), .Z(n13290) );
BUF_X4 U9391 ( .A(n13029), .Z(n13293) );
BUF_X4 U9392 ( .A(n13029), .Z(n13296) );
BUF_X4 U9393 ( .A(n13029), .Z(n13299) );
BUF_X4 U9394 ( .A(n13029), .Z(n13273) );
BUF_X4 U9395 ( .A(n13029), .Z(n13302) );
BUF_X4 U9396 ( .A(n13029), .Z(n13276) );
BUF_X4 U9397 ( .A(n13029), .Z(n13305) );
BUF_X4 U9398 ( .A(n13029), .Z(n13279) );
BUF_X4 U9399 ( .A(n13029), .Z(n13308) );
BUF_X4 U9400 ( .A(n13029), .Z(n13282) );
BUF_X4 U9401 ( .A(n13029), .Z(n13311) );
BUF_X4 U9402 ( .A(n13029), .Z(n13285) );
BUF_X4 U9403 ( .A(n13029), .Z(n13288) );
BUF_X4 U9404 ( .A(n13029), .Z(n13291) );
BUF_X4 U9405 ( .A(n13029), .Z(n13294) );
BUF_X4 U9406 ( .A(n13029), .Z(n13297) );
BUF_X4 U9407 ( .A(n13029), .Z(n13298) );
BUF_X4 U9408 ( .A(n13029), .Z(n13300) );
BUF_X4 U9409 ( .A(n13029), .Z(n13303) );
BUF_X4 U9410 ( .A(n13029), .Z(n13306) );
BUF_X4 U9411 ( .A(n13029), .Z(n13309) );
BUF_X4 U9412 ( .A(n13029), .Z(n13312) );
BUF_X4 U9413 ( .A(n13029), .Z(n13274) );
BUF_X4 U9414 ( .A(n13029), .Z(n13277) );
BUF_X4 U9415 ( .A(n13029), .Z(n13280) );
BUF_X4 U9416 ( .A(n13029), .Z(n13283) );
BUF_X4 U9417 ( .A(n13029), .Z(n13286) );
BUF_X4 U9418 ( .A(n13029), .Z(n13289) );
BUF_X4 U9419 ( .A(n13029), .Z(n13292) );
BUF_X4 U9420 ( .A(n13029), .Z(n13295) );
BUF_X4 U9421 ( .A(n13029), .Z(n13315) );
BUF_X4 U9422 ( .A(n13029), .Z(n13317) );
INV_X4 U9423 ( .A(n14731), .ZN(n14724) );
AND2_X2 U9424 ( .A1(n14700), .A2(n14715), .ZN(n13119) );
OR2_X2 U9425 ( .A1(n14957), .A2(n15425), .ZN(n13120) );
INV_X4 U9426 ( .A(n14690), .ZN(n13270) );
INV_X4 U9427 ( .A(n12990), .ZN(n13328) );
INV_X4 U9428 ( .A(n12990), .ZN(n13323) );
INV_X4 U9429 ( .A(n12990), .ZN(n13322) );
INV_X4 U9430 ( .A(n12990), .ZN(n13325) );
INV_X4 U9431 ( .A(n12990), .ZN(n13324) );
INV_X4 U9432 ( .A(n12990), .ZN(n13326) );
INV_X4 U9433 ( .A(n12990), .ZN(n13327) );
INV_X4 U9434 ( .A(n13124), .ZN(n13343) );
INV_X4 U9435 ( .A(n13124), .ZN(n13342) );
INV_X4 U9436 ( .A(n13124), .ZN(n13344) );
INV_X4 U9437 ( .A(n13126), .ZN(n13225) );
INV_X4 U9438 ( .A(n13123), .ZN(n13228) );
INV_X4 U9439 ( .A(n13127), .ZN(n13243) );
INV_X4 U9440 ( .A(n13125), .ZN(n13252) );
INV_X4 U9441 ( .A(n13126), .ZN(n13226) );
INV_X4 U9442 ( .A(n13123), .ZN(n13229) );
INV_X4 U9443 ( .A(n13127), .ZN(n13244) );
INV_X4 U9444 ( .A(n13125), .ZN(n13253) );
INV_X4 U9445 ( .A(n13125), .ZN(n13254) );
INV_X4 U9446 ( .A(n13126), .ZN(n13227) );
INV_X4 U9447 ( .A(n13123), .ZN(n13230) );
INV_X4 U9448 ( .A(n13127), .ZN(n13245) );
INV_X4 U9449 ( .A(n14690), .ZN(n13271) );
INV_X4 U9450 ( .A(n13017), .ZN(n13264) );
INV_X4 U9451 ( .A(n13017), .ZN(n13265) );
INV_X4 U9452 ( .A(n13017), .ZN(n13266) );
INV_X4 U9453 ( .A(n14718), .ZN(n13386) );
INV_X4 U9454 ( .A(n14000), .ZN(n13155) );
INV_X4 U9455 ( .A(n14000), .ZN(n13154) );
INV_X4 U9456 ( .A(n14721), .ZN(n13389) );
INV_X4 U9457 ( .A(n14728), .ZN(n13267) );
INV_X4 U9458 ( .A(n14718), .ZN(n13387) );
INV_X4 U9459 ( .A(n14721), .ZN(n13390) );
INV_X4 U9460 ( .A(n14001), .ZN(n13318) );
INV_X4 U9461 ( .A(n14001), .ZN(n13319) );
INV_X4 U9462 ( .A(n14728), .ZN(n13268) );
INV_X4 U9463 ( .A(n14718), .ZN(n13388) );
INV_X4 U9464 ( .A(n14721), .ZN(n13391) );
INV_X4 U9465 ( .A(n14001), .ZN(n13320) );
INV_X4 U9466 ( .A(n14728), .ZN(n13269) );
INV_X4 U9467 ( .A(n13352), .ZN(n13349) );
INV_X4 U9468 ( .A(n13352), .ZN(n13350) );
INV_X4 U9469 ( .A(n13352), .ZN(n13347) );
INV_X4 U9470 ( .A(n13352), .ZN(n13348) );
INV_X4 U9471 ( .A(n13352), .ZN(n13346) );
INV_X4 U9472 ( .A(n13352), .ZN(n13345) );
INV_X4 U9473 ( .A(n12990), .ZN(n13329) );
INV_X4 U9474 ( .A(n13352), .ZN(n13351) );
AND2_X2 U9475 ( .A1(n13437), .A2(n13427), .ZN(n13121) );
MUX2_X2 U9476 ( .A(n14368), .B(n13164), .S(n14165), .Z(n14163) );
MUX2_X2 U9477 ( .A(n14368), .B(n13164), .S(n14182), .Z(n14180) );
MUX2_X2 U9478 ( .A(n14368), .B(n13164), .S(n14157), .Z(n14155) );
MUX2_X2 U9479 ( .A(n14174), .B(n13164), .S(n14133), .Z(n14131) );
MUX2_X2 U9480 ( .A(n14368), .B(n13162), .S(n14149), .Z(n14147) );
MUX2_X2 U9481 ( .A(n14174), .B(n13163), .S(n14125), .Z(n14123) );
MUX2_X2 U9482 ( .A(n14174), .B(n13162), .S(n14117), .Z(n14115) );
MUX2_X2 U9483 ( .A(n14174), .B(n13162), .S(n14109), .Z(n14107) );
MUX2_X2 U9484 ( .A(n13096), .B(n13164), .S(n14093), .Z(n14091) );
MUX2_X2 U9485 ( .A(n13096), .B(n13163), .S(n14085), .Z(n14083) );
MUX2_X2 U9486 ( .A(n14174), .B(n13162), .S(n14101), .Z(n14099) );
MUX2_X2 U9487 ( .A(n13096), .B(n13163), .S(n14077), .Z(n14075) );
AND2_X2 U9488 ( .A1(n14242), .A2(n14243), .ZN(n13122) );
MUX2_X2 U9489 ( .A(n14368), .B(n13163), .S(n14173), .Z(n14171) );
MUX2_X2 U9490 ( .A(n14174), .B(n13162), .S(n14141), .Z(n14139) );
INV_X4 U9491 ( .A(n11114), .ZN(n13352) );
AND2_X2 U9492 ( .A1(n14697), .A2(n14700), .ZN(n13123) );
NOR2_X2 U9493 ( .A1(n14730), .A2(n14729), .ZN(n14732) );
AND2_X2 U9494 ( .A1(n14955), .A2(n11840), .ZN(n13124) );
AND2_X2 U9495 ( .A1(n14716), .A2(n14715), .ZN(n13125) );
AND2_X2 U9496 ( .A1(n14695), .A2(n14700), .ZN(n13126) );
AND2_X2 U9497 ( .A1(n14708), .A2(n14715), .ZN(n13127) );
INV_X4 U9498 ( .A(n13134), .ZN(n13396) );
INV_X4 U9499 ( .A(n13134), .ZN(n13395) );
INV_X4 U9500 ( .A(n13133), .ZN(n13151) );
INV_X4 U9501 ( .A(n13133), .ZN(n13153) );
INV_X4 U9502 ( .A(n13133), .ZN(n13152) );
AND2_X2 U9503 ( .A1(n13407), .A2(n14067), .ZN(n13128) );
INV_X4 U9504 ( .A(n13135), .ZN(n13337) );
INV_X4 U9505 ( .A(n13135), .ZN(n13336) );
INV_X4 U9506 ( .A(n13136), .ZN(n13330) );
INV_X4 U9507 ( .A(n13136), .ZN(n13331) );
INV_X4 U9508 ( .A(n13135), .ZN(n13338) );
INV_X4 U9509 ( .A(n13136), .ZN(n13332) );
INV_X4 U9510 ( .A(n13138), .ZN(n13366) );
INV_X4 U9511 ( .A(n13132), .ZN(n13369) );
INV_X4 U9512 ( .A(n13141), .ZN(n13372) );
INV_X4 U9513 ( .A(n13131), .ZN(n13378) );
INV_X4 U9514 ( .A(n13140), .ZN(n13381) );
INV_X4 U9515 ( .A(n13131), .ZN(n13377) );
INV_X4 U9516 ( .A(n13140), .ZN(n13380) );
INV_X4 U9517 ( .A(n13138), .ZN(n13365) );
INV_X4 U9518 ( .A(n13132), .ZN(n13368) );
INV_X4 U9519 ( .A(n13141), .ZN(n13371) );
INV_X4 U9520 ( .A(n13139), .ZN(n13393) );
INV_X4 U9521 ( .A(n13139), .ZN(n13392) );
INV_X4 U9522 ( .A(n13138), .ZN(n13367) );
INV_X4 U9523 ( .A(n13132), .ZN(n13370) );
INV_X4 U9524 ( .A(n13141), .ZN(n13373) );
INV_X4 U9525 ( .A(n13131), .ZN(n13379) );
INV_X4 U9526 ( .A(n13140), .ZN(n13382) );
INV_X4 U9527 ( .A(n13139), .ZN(n13394) );
INV_X4 U9528 ( .A(n13137), .ZN(n13339) );
INV_X4 U9529 ( .A(n13137), .ZN(n13340) );
INV_X4 U9530 ( .A(n13137), .ZN(n13341) );
NOR2_X2 U9531 ( .A1(rst_i), .A2(n13321), .ZN(n11114) );
XNOR2_X2 U9532 ( .A(n461), .B(n14220), .ZN(n14221) );
AND2_X2 U9533 ( .A1(n14067), .A2(n13093), .ZN(n13129) );
NOR2_X2 U9534 ( .A1(n345), .A2(n13998), .ZN(n13805) );
OR2_X2 U9535 ( .A1(n10118), .A2(rst_i), .ZN(n13131) );
OR2_X2 U9536 ( .A1(n10510), .A2(rst_i), .ZN(n13132) );
NOR2_X2 U9537 ( .A1(read_counter[0]), .A2(read_counter[1]), .ZN(n11840) );
NOR2_X2 U9538 ( .A1(n12076), .A2(read_counter[2]), .ZN(n12077) );
NAND3_X2 U9539 ( .A1(n9721), .A2(n9722), .A3(n9723), .ZN(n4431) );
NAND3_X2 U9540 ( .A1(n10905), .A2(n10906), .A3(n10907), .ZN(n4049) );
NAND3_X2 U9541 ( .A1(n9816), .A2(n9817), .A3(n9818), .ZN(n4400) );
NAND3_X2 U9542 ( .A1(n10902), .A2(n10903), .A3(n10904), .ZN(n4050) );
NAND3_X2 U9543 ( .A1(n9813), .A2(n9814), .A3(n9815), .ZN(n4401) );
NAND3_X2 U9544 ( .A1(n10899), .A2(n10900), .A3(n10901), .ZN(n4051) );
NAND3_X2 U9545 ( .A1(n9810), .A2(n9811), .A3(n9812), .ZN(n4402) );
NAND3_X2 U9546 ( .A1(n10896), .A2(n10897), .A3(n10898), .ZN(n4052) );
NAND3_X2 U9547 ( .A1(n9807), .A2(n9808), .A3(n9809), .ZN(n4403) );
NAND3_X2 U9548 ( .A1(n10893), .A2(n10894), .A3(n10895), .ZN(n4053) );
NAND3_X2 U9549 ( .A1(n9804), .A2(n9805), .A3(n9806), .ZN(n4404) );
NAND3_X2 U9550 ( .A1(n10890), .A2(n10891), .A3(n10892), .ZN(n4054) );
NAND3_X2 U9551 ( .A1(n9801), .A2(n9802), .A3(n9803), .ZN(n4405) );
NAND3_X2 U9552 ( .A1(n10887), .A2(n10888), .A3(n10889), .ZN(n4055) );
NAND3_X2 U9553 ( .A1(n9798), .A2(n9799), .A3(n9800), .ZN(n4406) );
NAND3_X2 U9554 ( .A1(n10884), .A2(n10885), .A3(n10886), .ZN(n4056) );
NAND3_X2 U9555 ( .A1(n9795), .A2(n9796), .A3(n9797), .ZN(n4407) );
NAND3_X2 U9556 ( .A1(n10881), .A2(n10882), .A3(n10883), .ZN(n4057) );
NAND3_X2 U9557 ( .A1(n9792), .A2(n9793), .A3(n9794), .ZN(n4408) );
NAND3_X2 U9558 ( .A1(n10878), .A2(n10879), .A3(n10880), .ZN(n4058) );
NAND3_X2 U9559 ( .A1(n9789), .A2(n9790), .A3(n9791), .ZN(n4409) );
NAND3_X2 U9560 ( .A1(n10875), .A2(n10876), .A3(n10877), .ZN(n4059) );
NAND3_X2 U9561 ( .A1(n9786), .A2(n9787), .A3(n9788), .ZN(n4410) );
NAND3_X2 U9562 ( .A1(n10872), .A2(n10873), .A3(n10874), .ZN(n4060) );
NAND3_X2 U9563 ( .A1(n9783), .A2(n9784), .A3(n9785), .ZN(n4411) );
NAND3_X2 U9564 ( .A1(n10869), .A2(n10870), .A3(n10871), .ZN(n4061) );
NAND3_X2 U9565 ( .A1(n9780), .A2(n9781), .A3(n9782), .ZN(n4412) );
NAND3_X2 U9566 ( .A1(n10866), .A2(n10867), .A3(n10868), .ZN(n4062) );
NAND3_X2 U9567 ( .A1(n9777), .A2(n9778), .A3(n9779), .ZN(n4413) );
NAND3_X2 U9568 ( .A1(n10863), .A2(n10864), .A3(n10865), .ZN(n4063) );
NAND3_X2 U9569 ( .A1(n9774), .A2(n9775), .A3(n9776), .ZN(n4414) );
NAND3_X2 U9570 ( .A1(n10860), .A2(n10861), .A3(n10862), .ZN(n4064) );
NAND3_X2 U9571 ( .A1(n9771), .A2(n9772), .A3(n9773), .ZN(n4415) );
NAND3_X2 U9572 ( .A1(n10857), .A2(n10858), .A3(n10859), .ZN(n4065) );
NAND3_X2 U9573 ( .A1(n9768), .A2(n9769), .A3(n9770), .ZN(n4416) );
NAND3_X2 U9574 ( .A1(n10854), .A2(n10855), .A3(n10856), .ZN(n4066) );
NAND3_X2 U9575 ( .A1(n9765), .A2(n9766), .A3(n9767), .ZN(n4417) );
NAND3_X2 U9576 ( .A1(n10851), .A2(n10852), .A3(n10853), .ZN(n4067) );
NAND3_X2 U9577 ( .A1(n9762), .A2(n9763), .A3(n9764), .ZN(n4418) );
NAND3_X2 U9578 ( .A1(n10848), .A2(n10849), .A3(n10850), .ZN(n4068) );
NAND3_X2 U9579 ( .A1(n9759), .A2(n9760), .A3(n9761), .ZN(n4419) );
NAND3_X2 U9580 ( .A1(n10845), .A2(n10846), .A3(n10847), .ZN(n4069) );
NAND3_X2 U9581 ( .A1(n9756), .A2(n9757), .A3(n9758), .ZN(n4420) );
NAND3_X2 U9582 ( .A1(n10842), .A2(n10843), .A3(n10844), .ZN(n4070) );
NAND3_X2 U9583 ( .A1(n9753), .A2(n9754), .A3(n9755), .ZN(n4421) );
NAND3_X2 U9584 ( .A1(n10839), .A2(n10840), .A3(n10841), .ZN(n4071) );
NAND3_X2 U9585 ( .A1(n9750), .A2(n9751), .A3(n9752), .ZN(n4422) );
NAND3_X2 U9586 ( .A1(n10836), .A2(n10837), .A3(n10838), .ZN(n4072) );
NAND3_X2 U9587 ( .A1(n9747), .A2(n9748), .A3(n9749), .ZN(n4423) );
NAND3_X2 U9588 ( .A1(n10833), .A2(n10834), .A3(n10835), .ZN(n4073) );
NAND3_X2 U9589 ( .A1(n9744), .A2(n9745), .A3(n9746), .ZN(n4424) );
NAND3_X2 U9590 ( .A1(n10830), .A2(n10831), .A3(n10832), .ZN(n4074) );
NAND3_X2 U9591 ( .A1(n9741), .A2(n9742), .A3(n9743), .ZN(n4425) );
NAND3_X2 U9592 ( .A1(n10827), .A2(n10828), .A3(n10829), .ZN(n4075) );
NAND3_X2 U9593 ( .A1(n9738), .A2(n9739), .A3(n9740), .ZN(n4426) );
NAND3_X2 U9594 ( .A1(n10824), .A2(n10825), .A3(n10826), .ZN(n4076) );
NAND3_X2 U9595 ( .A1(n9735), .A2(n9736), .A3(n9737), .ZN(n4427) );
NAND3_X2 U9596 ( .A1(n10821), .A2(n10822), .A3(n10823), .ZN(n4077) );
NAND3_X2 U9597 ( .A1(n9732), .A2(n9733), .A3(n9734), .ZN(n4428) );
NAND3_X2 U9598 ( .A1(n10818), .A2(n10819), .A3(n10820), .ZN(n4078) );
NAND3_X2 U9599 ( .A1(n9729), .A2(n9730), .A3(n9731), .ZN(n4429) );
NAND3_X2 U9600 ( .A1(n10815), .A2(n10816), .A3(n10817), .ZN(n4079) );
NAND3_X2 U9601 ( .A1(n9726), .A2(n9727), .A3(n9728), .ZN(n4430) );
NAND3_X2 U9602 ( .A1(n10810), .A2(n10811), .A3(n10812), .ZN(n4080) );
NOR2_X2 U9603 ( .A1(n13395), .A2(n12854), .ZN(n11865) );
NOR2_X2 U9604 ( .A1(n13395), .A2(n12862), .ZN(n11893) );
NOR2_X2 U9605 ( .A1(n13395), .A2(n12852), .ZN(n11853) );
NOR2_X2 U9606 ( .A1(n13395), .A2(n12856), .ZN(n11872) );
NOR2_X2 U9607 ( .A1(n13395), .A2(n12858), .ZN(n11879) );
NOR2_X2 U9608 ( .A1(n13395), .A2(n12860), .ZN(n11886) );
NOR2_X2 U9609 ( .A1(n13396), .A2(n12864), .ZN(n11900) );
NOR2_X2 U9610 ( .A1(n13395), .A2(n12866), .ZN(n11907) );
NOR2_X2 U9611 ( .A1(n13395), .A2(n12868), .ZN(n11914) );
NOR2_X2 U9612 ( .A1(n13395), .A2(n12870), .ZN(n11921) );
NOR2_X2 U9613 ( .A1(n13395), .A2(n12872), .ZN(n11928) );
NOR2_X2 U9614 ( .A1(n13395), .A2(n12874), .ZN(n11935) );
NOR2_X2 U9615 ( .A1(n13395), .A2(n12876), .ZN(n11942) );
NOR2_X2 U9616 ( .A1(n13395), .A2(n12878), .ZN(n11949) );
NOR2_X2 U9617 ( .A1(n13395), .A2(n12880), .ZN(n11956) );
NOR2_X2 U9618 ( .A1(n13396), .A2(n12882), .ZN(n11963) );
NOR2_X2 U9619 ( .A1(n13396), .A2(n12884), .ZN(n11970) );
NOR2_X2 U9620 ( .A1(n13396), .A2(n12886), .ZN(n11977) );
NOR2_X2 U9621 ( .A1(n13396), .A2(n12888), .ZN(n11984) );
NOR2_X2 U9622 ( .A1(n13396), .A2(n12890), .ZN(n11991) );
NOR2_X2 U9623 ( .A1(n13396), .A2(n12892), .ZN(n11998) );
NOR2_X2 U9624 ( .A1(n13396), .A2(n12894), .ZN(n12005) );
NOR2_X2 U9625 ( .A1(n13396), .A2(n12906), .ZN(n12047) );
NOR2_X2 U9626 ( .A1(n13396), .A2(n12908), .ZN(n12054) );
NOR2_X2 U9627 ( .A1(n13396), .A2(n12910), .ZN(n12061) );
NOR2_X2 U9628 ( .A1(n13396), .A2(n12912), .ZN(n12068) );
NOR2_X2 U9629 ( .A1(n13395), .A2(n12914), .ZN(n12075) );
NOR2_X2 U9630 ( .A1(n15426), .A2(rst_i), .ZN(n9301) );
NAND3_X2 U9631 ( .A1(n10974), .A2(n10975), .A3(n10976), .ZN(n4027) );
NAND3_X2 U9632 ( .A1(n10971), .A2(n10972), .A3(n10973), .ZN(n4028) );
NAND3_X2 U9633 ( .A1(n10968), .A2(n10969), .A3(n10970), .ZN(n4029) );
NAND3_X2 U9634 ( .A1(n10965), .A2(n10966), .A3(n10967), .ZN(n4030) );
NAND3_X2 U9635 ( .A1(n10962), .A2(n10963), .A3(n10964), .ZN(n4031) );
NAND3_X2 U9636 ( .A1(n10959), .A2(n10960), .A3(n10961), .ZN(n4032) );
NAND3_X2 U9637 ( .A1(n10956), .A2(n10957), .A3(n10958), .ZN(n4033) );
NAND3_X2 U9638 ( .A1(n10953), .A2(n10954), .A3(n10955), .ZN(n4034) );
NAND3_X2 U9639 ( .A1(n10950), .A2(n10951), .A3(n10952), .ZN(n4035) );
NAND3_X2 U9640 ( .A1(n10947), .A2(n10948), .A3(n10949), .ZN(n4036) );
NAND3_X2 U9641 ( .A1(n10944), .A2(n10945), .A3(n10946), .ZN(n4037) );
NAND3_X2 U9642 ( .A1(n10941), .A2(n10942), .A3(n10943), .ZN(n4038) );
NAND3_X2 U9643 ( .A1(n10938), .A2(n10939), .A3(n10940), .ZN(n4039) );
NAND3_X2 U9644 ( .A1(n10935), .A2(n10936), .A3(n10937), .ZN(n4040) );
NAND3_X2 U9645 ( .A1(n10932), .A2(n10933), .A3(n10934), .ZN(n4041) );
NAND3_X2 U9646 ( .A1(n10929), .A2(n10930), .A3(n10931), .ZN(n4042) );
NAND3_X2 U9647 ( .A1(n10926), .A2(n10927), .A3(n10928), .ZN(n4043) );
NAND3_X2 U9648 ( .A1(n10923), .A2(n10924), .A3(n10925), .ZN(n4044) );
NAND3_X2 U9649 ( .A1(n10920), .A2(n10921), .A3(n10922), .ZN(n4045) );
NAND3_X2 U9650 ( .A1(n10917), .A2(n10918), .A3(n10919), .ZN(n4046) );
NAND3_X2 U9651 ( .A1(n10914), .A2(n10915), .A3(n10916), .ZN(n4047) );
NAND3_X2 U9652 ( .A1(n10909), .A2(n10910), .A3(n10911), .ZN(n4048) );
AND3_X2 U9653 ( .A1(n14933), .A2(n341), .A3(n13437), .ZN(n13133) );
AND2_X2 U9654 ( .A1(cmd_o[0]), .A2(n14953), .ZN(n13134) );
NOR3_X2 U9655 ( .A1(n12010), .A2(n12011), .A3(n12012), .ZN(n12009) );
NOR2_X2 U9656 ( .A1(n13396), .A2(n12896), .ZN(n12012) );
NOR3_X2 U9657 ( .A1(n12017), .A2(n12018), .A3(n12019), .ZN(n12016) );
NOR2_X2 U9658 ( .A1(n13396), .A2(n12898), .ZN(n12019) );
NOR3_X2 U9659 ( .A1(n12024), .A2(n12025), .A3(n12026), .ZN(n12023) );
NOR2_X2 U9660 ( .A1(n13396), .A2(n12900), .ZN(n12026) );
NOR3_X2 U9661 ( .A1(n12031), .A2(n12032), .A3(n12033), .ZN(n12030) );
NOR2_X2 U9662 ( .A1(n13396), .A2(n12902), .ZN(n12033) );
NOR3_X2 U9663 ( .A1(n12038), .A2(n12039), .A3(n12040), .ZN(n12037) );
NOR2_X2 U9664 ( .A1(n13396), .A2(n12904), .ZN(n12040) );
NAND3_X2 U9665 ( .A1(n347), .A2(n14953), .A3(n8326), .ZN(n12076) );
NAND3_X2 U9666 ( .A1(read_counter[1]), .A2(n14952), .A3(n12077), .ZN(n13135));
OR3_X2 U9667 ( .A1(n14952), .A2(read_counter[1]), .A3(n14957), .ZN(n13136));
AND3_X2 U9668 ( .A1(read_counter[1]), .A2(read_counter[0]), .A3(n12077),.ZN(n13137) );
OR2_X2 U9669 ( .A1(n10609), .A2(rst_i), .ZN(n13138) );
OR2_X2 U9670 ( .A1(n10212), .A2(rst_i), .ZN(n13139) );
OR2_X2 U9671 ( .A1(n10019), .A2(rst_i), .ZN(n13140) );
OR2_X2 U9672 ( .A1(n10411), .A2(rst_i), .ZN(n13141) );
NAND3_X2 U9673 ( .A1(n14956), .A2(n11837), .A3(n11840), .ZN(n11839) );
INV_X4 U9674 ( .A(rst_i), .ZN(n14953) );
NAND3_X2 U9675 ( .A1(cmd_o[2]), .A2(n14953), .A3(n15426), .ZN(n9300) );
NAND3_X2 U9676 ( .A1(n11843), .A2(n13395), .A3(n11844), .ZN(n3694) );
NAND3_X2 U9677 ( .A1(n10209), .A2(n10210), .A3(n10211), .ZN(n4273) );
NAND3_X2 U9678 ( .A1(n10206), .A2(n10207), .A3(n10208), .ZN(n4274) );
NAND3_X2 U9679 ( .A1(n10203), .A2(n10204), .A3(n10205), .ZN(n4275) );
NAND3_X2 U9680 ( .A1(n10200), .A2(n10201), .A3(n10202), .ZN(n4276) );
NAND3_X2 U9681 ( .A1(n10197), .A2(n10198), .A3(n10199), .ZN(n4277) );
NAND3_X2 U9682 ( .A1(n10194), .A2(n10195), .A3(n10196), .ZN(n4278) );
NAND3_X2 U9683 ( .A1(n10191), .A2(n10192), .A3(n10193), .ZN(n4279) );
NAND3_X2 U9684 ( .A1(n10188), .A2(n10189), .A3(n10190), .ZN(n4280) );
NAND3_X2 U9685 ( .A1(n10185), .A2(n10186), .A3(n10187), .ZN(n4281) );
NAND3_X2 U9686 ( .A1(n10182), .A2(n10183), .A3(n10184), .ZN(n4282) );
NAND3_X2 U9687 ( .A1(n10179), .A2(n10180), .A3(n10181), .ZN(n4283) );
NAND3_X2 U9688 ( .A1(n10176), .A2(n10177), .A3(n10178), .ZN(n4284) );
NAND3_X2 U9689 ( .A1(n10173), .A2(n10174), .A3(n10175), .ZN(n4285) );
NAND3_X2 U9690 ( .A1(n10170), .A2(n10171), .A3(n10172), .ZN(n4286) );
NAND3_X2 U9691 ( .A1(n10167), .A2(n10168), .A3(n10169), .ZN(n4287) );
NAND3_X2 U9692 ( .A1(n10164), .A2(n10165), .A3(n10166), .ZN(n4288) );
NAND3_X2 U9693 ( .A1(n10161), .A2(n10162), .A3(n10163), .ZN(n4289) );
NAND3_X2 U9694 ( .A1(n10158), .A2(n10159), .A3(n10160), .ZN(n4290) );
NAND3_X2 U9695 ( .A1(n10155), .A2(n10156), .A3(n10157), .ZN(n4291) );
NAND3_X2 U9696 ( .A1(n10152), .A2(n10153), .A3(n10154), .ZN(n4292) );
NAND3_X2 U9697 ( .A1(n10149), .A2(n10150), .A3(n10151), .ZN(n4293) );
NAND3_X2 U9698 ( .A1(n10146), .A2(n10147), .A3(n10148), .ZN(n4294) );
NAND3_X2 U9699 ( .A1(n10143), .A2(n10144), .A3(n10145), .ZN(n4295) );
NAND3_X2 U9700 ( .A1(n10140), .A2(n10141), .A3(n10142), .ZN(n4296) );
NAND3_X2 U9701 ( .A1(n10137), .A2(n10138), .A3(n10139), .ZN(n4297) );
NAND3_X2 U9702 ( .A1(n10134), .A2(n10135), .A3(n10136), .ZN(n4298) );
NAND3_X2 U9703 ( .A1(n10131), .A2(n10132), .A3(n10133), .ZN(n4299) );
NAND3_X2 U9704 ( .A1(n10128), .A2(n10129), .A3(n10130), .ZN(n4300) );
NAND3_X2 U9705 ( .A1(n10125), .A2(n10126), .A3(n10127), .ZN(n4301) );
NAND3_X2 U9706 ( .A1(n10122), .A2(n10123), .A3(n10124), .ZN(n4302) );
NAND3_X2 U9707 ( .A1(n10119), .A2(n10120), .A3(n10121), .ZN(n4303) );
NAND3_X2 U9708 ( .A1(n9315), .A2(n9316), .A3(n9317), .ZN(n4528) );
NAND3_X2 U9709 ( .A1(n10020), .A2(n10021), .A3(n10022), .ZN(n4335) );
NAND3_X2 U9710 ( .A1(n9921), .A2(n9922), .A3(n9923), .ZN(n4367) );
NAND3_X2 U9711 ( .A1(n9820), .A2(n9821), .A3(n9822), .ZN(n4399) );
NAND3_X2 U9712 ( .A1(n9621), .A2(n9622), .A3(n9623), .ZN(n4463) );
NAND3_X2 U9713 ( .A1(n11004), .A2(n11005), .A3(n11006), .ZN(n4017) );
NAND3_X2 U9714 ( .A1(n10806), .A2(n10807), .A3(n10808), .ZN(n4081) );
NAND3_X2 U9715 ( .A1(n10705), .A2(n10706), .A3(n10707), .ZN(n4113) );
NAND3_X2 U9716 ( .A1(n10606), .A2(n10607), .A3(n10608), .ZN(n4145) );
NAND3_X2 U9717 ( .A1(n10507), .A2(n10508), .A3(n10509), .ZN(n4177) );
NAND3_X2 U9718 ( .A1(n10408), .A2(n10409), .A3(n10410), .ZN(n4209) );
NAND3_X2 U9719 ( .A1(n10308), .A2(n10309), .A3(n10310), .ZN(n4241) );
NAND3_X2 U9720 ( .A1(n10115), .A2(n10116), .A3(n10117), .ZN(n4304) );
NAND3_X2 U9721 ( .A1(n10016), .A2(n10017), .A3(n10018), .ZN(n4336) );
NAND3_X2 U9722 ( .A1(n9915), .A2(n9916), .A3(n9917), .ZN(n4368) );
NAND3_X2 U9723 ( .A1(n9716), .A2(n9717), .A3(n9718), .ZN(n4432) );
NAND3_X2 U9724 ( .A1(n9614), .A2(n9615), .A3(n9616), .ZN(n4464) );
NAND3_X2 U9725 ( .A1(n11001), .A2(n11002), .A3(n11003), .ZN(n4018) );
NAND3_X2 U9726 ( .A1(n10803), .A2(n10804), .A3(n10805), .ZN(n4082) );
NAND3_X2 U9727 ( .A1(n10702), .A2(n10703), .A3(n10704), .ZN(n4114) );
NAND3_X2 U9728 ( .A1(n10603), .A2(n10604), .A3(n10605), .ZN(n4146) );
NAND3_X2 U9729 ( .A1(n10504), .A2(n10505), .A3(n10506), .ZN(n4178) );
NAND3_X2 U9730 ( .A1(n10405), .A2(n10406), .A3(n10407), .ZN(n4210) );
NAND3_X2 U9731 ( .A1(n10305), .A2(n10306), .A3(n10307), .ZN(n4242) );
NAND3_X2 U9732 ( .A1(n10112), .A2(n10113), .A3(n10114), .ZN(n4305) );
NAND3_X2 U9733 ( .A1(n10013), .A2(n10014), .A3(n10015), .ZN(n4337) );
NAND3_X2 U9734 ( .A1(n9912), .A2(n9913), .A3(n9914), .ZN(n4369) );
NAND3_X2 U9735 ( .A1(n9713), .A2(n9714), .A3(n9715), .ZN(n4433) );
NAND3_X2 U9736 ( .A1(n9611), .A2(n9612), .A3(n9613), .ZN(n4465) );
NAND3_X2 U9737 ( .A1(n10998), .A2(n10999), .A3(n11000), .ZN(n4019) );
NAND3_X2 U9738 ( .A1(n10800), .A2(n10801), .A3(n10802), .ZN(n4083) );
NAND3_X2 U9739 ( .A1(n10699), .A2(n10700), .A3(n10701), .ZN(n4115) );
NAND3_X2 U9740 ( .A1(n10600), .A2(n10601), .A3(n10602), .ZN(n4147) );
NAND3_X2 U9741 ( .A1(n10501), .A2(n10502), .A3(n10503), .ZN(n4179) );
NAND3_X2 U9742 ( .A1(n10402), .A2(n10403), .A3(n10404), .ZN(n4211) );
NAND3_X2 U9743 ( .A1(n10302), .A2(n10303), .A3(n10304), .ZN(n4243) );
NAND3_X2 U9744 ( .A1(n10109), .A2(n10110), .A3(n10111), .ZN(n4306) );
NAND3_X2 U9745 ( .A1(n10010), .A2(n10011), .A3(n10012), .ZN(n4338) );
NAND3_X2 U9746 ( .A1(n9909), .A2(n9910), .A3(n9911), .ZN(n4370) );
NAND3_X2 U9747 ( .A1(n9710), .A2(n9711), .A3(n9712), .ZN(n4434) );
NAND3_X2 U9748 ( .A1(n9608), .A2(n9609), .A3(n9610), .ZN(n4466) );
NAND3_X2 U9749 ( .A1(n10995), .A2(n10996), .A3(n10997), .ZN(n4020) );
NAND3_X2 U9750 ( .A1(n10797), .A2(n10798), .A3(n10799), .ZN(n4084) );
NAND3_X2 U9751 ( .A1(n10696), .A2(n10697), .A3(n10698), .ZN(n4116) );
NAND3_X2 U9752 ( .A1(n10597), .A2(n10598), .A3(n10599), .ZN(n4148) );
NAND3_X2 U9753 ( .A1(n10498), .A2(n10499), .A3(n10500), .ZN(n4180) );
NAND3_X2 U9754 ( .A1(n10399), .A2(n10400), .A3(n10401), .ZN(n4212) );
NAND3_X2 U9755 ( .A1(n10299), .A2(n10300), .A3(n10301), .ZN(n4244) );
NAND3_X2 U9756 ( .A1(n10106), .A2(n10107), .A3(n10108), .ZN(n4307) );
NAND3_X2 U9757 ( .A1(n10007), .A2(n10008), .A3(n10009), .ZN(n4339) );
NAND3_X2 U9758 ( .A1(n9906), .A2(n9907), .A3(n9908), .ZN(n4371) );
NAND3_X2 U9759 ( .A1(n9707), .A2(n9708), .A3(n9709), .ZN(n4435) );
NAND3_X2 U9760 ( .A1(n9605), .A2(n9606), .A3(n9607), .ZN(n4467) );
NAND3_X2 U9761 ( .A1(n10992), .A2(n10993), .A3(n10994), .ZN(n4021) );
NAND3_X2 U9762 ( .A1(n10794), .A2(n10795), .A3(n10796), .ZN(n4085) );
NAND3_X2 U9763 ( .A1(n10693), .A2(n10694), .A3(n10695), .ZN(n4117) );
NAND3_X2 U9764 ( .A1(n10594), .A2(n10595), .A3(n10596), .ZN(n4149) );
NAND3_X2 U9765 ( .A1(n10495), .A2(n10496), .A3(n10497), .ZN(n4181) );
NAND3_X2 U9766 ( .A1(n10396), .A2(n10397), .A3(n10398), .ZN(n4213) );
NAND3_X2 U9767 ( .A1(n10296), .A2(n10297), .A3(n10298), .ZN(n4245) );
NAND3_X2 U9768 ( .A1(n10103), .A2(n10104), .A3(n10105), .ZN(n4308) );
NAND3_X2 U9769 ( .A1(n10004), .A2(n10005), .A3(n10006), .ZN(n4340) );
NAND3_X2 U9770 ( .A1(n9903), .A2(n9904), .A3(n9905), .ZN(n4372) );
NAND3_X2 U9771 ( .A1(n9704), .A2(n9705), .A3(n9706), .ZN(n4436) );
NAND3_X2 U9772 ( .A1(n9602), .A2(n9603), .A3(n9604), .ZN(n4468) );
NAND3_X2 U9773 ( .A1(n10989), .A2(n10990), .A3(n10991), .ZN(n4022) );
NAND3_X2 U9774 ( .A1(n10791), .A2(n10792), .A3(n10793), .ZN(n4086) );
NAND3_X2 U9775 ( .A1(n10690), .A2(n10691), .A3(n10692), .ZN(n4118) );
NAND3_X2 U9776 ( .A1(n10591), .A2(n10592), .A3(n10593), .ZN(n4150) );
NAND3_X2 U9777 ( .A1(n10492), .A2(n10493), .A3(n10494), .ZN(n4182) );
NAND3_X2 U9778 ( .A1(n10393), .A2(n10394), .A3(n10395), .ZN(n4214) );
NAND3_X2 U9779 ( .A1(n10293), .A2(n10294), .A3(n10295), .ZN(n4246) );
NAND3_X2 U9780 ( .A1(n10100), .A2(n10101), .A3(n10102), .ZN(n4309) );
NAND3_X2 U9781 ( .A1(n10001), .A2(n10002), .A3(n10003), .ZN(n4341) );
NAND3_X2 U9782 ( .A1(n9900), .A2(n9901), .A3(n9902), .ZN(n4373) );
NAND3_X2 U9783 ( .A1(n9701), .A2(n9702), .A3(n9703), .ZN(n4437) );
NAND3_X2 U9784 ( .A1(n9599), .A2(n9600), .A3(n9601), .ZN(n4469) );
NAND3_X2 U9785 ( .A1(n10986), .A2(n10987), .A3(n10988), .ZN(n4023) );
NAND3_X2 U9786 ( .A1(n10788), .A2(n10789), .A3(n10790), .ZN(n4087) );
NAND3_X2 U9787 ( .A1(n10687), .A2(n10688), .A3(n10689), .ZN(n4119) );
NAND3_X2 U9788 ( .A1(n10588), .A2(n10589), .A3(n10590), .ZN(n4151) );
NAND3_X2 U9789 ( .A1(n10489), .A2(n10490), .A3(n10491), .ZN(n4183) );
NAND3_X2 U9790 ( .A1(n10390), .A2(n10391), .A3(n10392), .ZN(n4215) );
NAND3_X2 U9791 ( .A1(n10290), .A2(n10291), .A3(n10292), .ZN(n4247) );
NAND3_X2 U9792 ( .A1(n10097), .A2(n10098), .A3(n10099), .ZN(n4310) );
NAND3_X2 U9793 ( .A1(n9998), .A2(n9999), .A3(n10000), .ZN(n4342) );
NAND3_X2 U9794 ( .A1(n9897), .A2(n9898), .A3(n9899), .ZN(n4374) );
NAND3_X2 U9795 ( .A1(n9698), .A2(n9699), .A3(n9700), .ZN(n4438) );
NAND3_X2 U9796 ( .A1(n9596), .A2(n9597), .A3(n9598), .ZN(n4470) );
NAND3_X2 U9797 ( .A1(n10983), .A2(n10984), .A3(n10985), .ZN(n4024) );
NAND3_X2 U9798 ( .A1(n10785), .A2(n10786), .A3(n10787), .ZN(n4088) );
NAND3_X2 U9799 ( .A1(n10684), .A2(n10685), .A3(n10686), .ZN(n4120) );
NAND3_X2 U9800 ( .A1(n10585), .A2(n10586), .A3(n10587), .ZN(n4152) );
NAND3_X2 U9801 ( .A1(n10486), .A2(n10487), .A3(n10488), .ZN(n4184) );
NAND3_X2 U9802 ( .A1(n10387), .A2(n10388), .A3(n10389), .ZN(n4216) );
NAND3_X2 U9803 ( .A1(n10287), .A2(n10288), .A3(n10289), .ZN(n4248) );
NAND3_X2 U9804 ( .A1(n10094), .A2(n10095), .A3(n10096), .ZN(n4311) );
NAND3_X2 U9805 ( .A1(n9995), .A2(n9996), .A3(n9997), .ZN(n4343) );
NAND3_X2 U9806 ( .A1(n9894), .A2(n9895), .A3(n9896), .ZN(n4375) );
NAND3_X2 U9807 ( .A1(n9695), .A2(n9696), .A3(n9697), .ZN(n4439) );
NAND3_X2 U9808 ( .A1(n9593), .A2(n9594), .A3(n9595), .ZN(n4471) );
NAND3_X2 U9809 ( .A1(n10980), .A2(n10981), .A3(n10982), .ZN(n4025) );
NAND3_X2 U9810 ( .A1(n10782), .A2(n10783), .A3(n10784), .ZN(n4089) );
NAND3_X2 U9811 ( .A1(n10681), .A2(n10682), .A3(n10683), .ZN(n4121) );
NAND3_X2 U9812 ( .A1(n10582), .A2(n10583), .A3(n10584), .ZN(n4153) );
NAND3_X2 U9813 ( .A1(n10483), .A2(n10484), .A3(n10485), .ZN(n4185) );
NAND3_X2 U9814 ( .A1(n10384), .A2(n10385), .A3(n10386), .ZN(n4217) );
NAND3_X2 U9815 ( .A1(n10284), .A2(n10285), .A3(n10286), .ZN(n4249) );
NAND3_X2 U9816 ( .A1(n10091), .A2(n10092), .A3(n10093), .ZN(n4312) );
NAND3_X2 U9817 ( .A1(n9992), .A2(n9993), .A3(n9994), .ZN(n4344) );
NAND3_X2 U9818 ( .A1(n9891), .A2(n9892), .A3(n9893), .ZN(n4376) );
NAND3_X2 U9819 ( .A1(n9692), .A2(n9693), .A3(n9694), .ZN(n4440) );
NAND3_X2 U9820 ( .A1(n9590), .A2(n9591), .A3(n9592), .ZN(n4472) );
NAND3_X2 U9821 ( .A1(n10977), .A2(n10978), .A3(n10979), .ZN(n4026) );
NAND3_X2 U9822 ( .A1(n10779), .A2(n10780), .A3(n10781), .ZN(n4090) );
NAND3_X2 U9823 ( .A1(n10678), .A2(n10679), .A3(n10680), .ZN(n4122) );
NAND3_X2 U9824 ( .A1(n10579), .A2(n10580), .A3(n10581), .ZN(n4154) );
NAND3_X2 U9825 ( .A1(n10480), .A2(n10481), .A3(n10482), .ZN(n4186) );
NAND3_X2 U9826 ( .A1(n10381), .A2(n10382), .A3(n10383), .ZN(n4218) );
NAND3_X2 U9827 ( .A1(n10281), .A2(n10282), .A3(n10283), .ZN(n4250) );
NAND3_X2 U9828 ( .A1(n10088), .A2(n10089), .A3(n10090), .ZN(n4313) );
NAND3_X2 U9829 ( .A1(n9989), .A2(n9990), .A3(n9991), .ZN(n4345) );
NAND3_X2 U9830 ( .A1(n9888), .A2(n9889), .A3(n9890), .ZN(n4377) );
NAND3_X2 U9831 ( .A1(n9689), .A2(n9690), .A3(n9691), .ZN(n4441) );
NAND3_X2 U9832 ( .A1(n9587), .A2(n9588), .A3(n9589), .ZN(n4473) );
NAND3_X2 U9833 ( .A1(n10776), .A2(n10777), .A3(n10778), .ZN(n4091) );
NAND3_X2 U9834 ( .A1(n10675), .A2(n10676), .A3(n10677), .ZN(n4123) );
NAND3_X2 U9835 ( .A1(n10576), .A2(n10577), .A3(n10578), .ZN(n4155) );
NAND3_X2 U9836 ( .A1(n10477), .A2(n10478), .A3(n10479), .ZN(n4187) );
NAND3_X2 U9837 ( .A1(n10378), .A2(n10379), .A3(n10380), .ZN(n4219) );
NAND3_X2 U9838 ( .A1(n10278), .A2(n10279), .A3(n10280), .ZN(n4251) );
NAND3_X2 U9839 ( .A1(n10085), .A2(n10086), .A3(n10087), .ZN(n4314) );
NAND3_X2 U9840 ( .A1(n9986), .A2(n9987), .A3(n9988), .ZN(n4346) );
NAND3_X2 U9841 ( .A1(n9885), .A2(n9886), .A3(n9887), .ZN(n4378) );
NAND3_X2 U9842 ( .A1(n9686), .A2(n9687), .A3(n9688), .ZN(n4442) );
NAND3_X2 U9843 ( .A1(n9584), .A2(n9585), .A3(n9586), .ZN(n4474) );
NAND3_X2 U9844 ( .A1(n10773), .A2(n10774), .A3(n10775), .ZN(n4092) );
NAND3_X2 U9845 ( .A1(n10672), .A2(n10673), .A3(n10674), .ZN(n4124) );
NAND3_X2 U9846 ( .A1(n10573), .A2(n10574), .A3(n10575), .ZN(n4156) );
NAND3_X2 U9847 ( .A1(n10474), .A2(n10475), .A3(n10476), .ZN(n4188) );
NAND3_X2 U9848 ( .A1(n10375), .A2(n10376), .A3(n10377), .ZN(n4220) );
NAND3_X2 U9849 ( .A1(n10275), .A2(n10276), .A3(n10277), .ZN(n4252) );
NAND3_X2 U9850 ( .A1(n10082), .A2(n10083), .A3(n10084), .ZN(n4315) );
NAND3_X2 U9851 ( .A1(n9983), .A2(n9984), .A3(n9985), .ZN(n4347) );
NAND3_X2 U9852 ( .A1(n9882), .A2(n9883), .A3(n9884), .ZN(n4379) );
NAND3_X2 U9853 ( .A1(n9683), .A2(n9684), .A3(n9685), .ZN(n4443) );
NAND3_X2 U9854 ( .A1(n9581), .A2(n9582), .A3(n9583), .ZN(n4475) );
NAND3_X2 U9855 ( .A1(n10770), .A2(n10771), .A3(n10772), .ZN(n4093) );
NAND3_X2 U9856 ( .A1(n10669), .A2(n10670), .A3(n10671), .ZN(n4125) );
NAND3_X2 U9857 ( .A1(n10570), .A2(n10571), .A3(n10572), .ZN(n4157) );
NAND3_X2 U9858 ( .A1(n10471), .A2(n10472), .A3(n10473), .ZN(n4189) );
NAND3_X2 U9859 ( .A1(n10372), .A2(n10373), .A3(n10374), .ZN(n4221) );
NAND3_X2 U9860 ( .A1(n10272), .A2(n10273), .A3(n10274), .ZN(n4253) );
NAND3_X2 U9861 ( .A1(n10079), .A2(n10080), .A3(n10081), .ZN(n4316) );
NAND3_X2 U9862 ( .A1(n9980), .A2(n9981), .A3(n9982), .ZN(n4348) );
NAND3_X2 U9863 ( .A1(n9879), .A2(n9880), .A3(n9881), .ZN(n4380) );
NAND3_X2 U9864 ( .A1(n9680), .A2(n9681), .A3(n9682), .ZN(n4444) );
NAND3_X2 U9865 ( .A1(n9578), .A2(n9579), .A3(n9580), .ZN(n4476) );
NAND3_X2 U9866 ( .A1(n10767), .A2(n10768), .A3(n10769), .ZN(n4094) );
NAND3_X2 U9867 ( .A1(n10666), .A2(n10667), .A3(n10668), .ZN(n4126) );
NAND3_X2 U9868 ( .A1(n10567), .A2(n10568), .A3(n10569), .ZN(n4158) );
NAND3_X2 U9869 ( .A1(n10468), .A2(n10469), .A3(n10470), .ZN(n4190) );
NAND3_X2 U9870 ( .A1(n10369), .A2(n10370), .A3(n10371), .ZN(n4222) );
NAND3_X2 U9871 ( .A1(n10269), .A2(n10270), .A3(n10271), .ZN(n4254) );
NAND3_X2 U9872 ( .A1(n10076), .A2(n10077), .A3(n10078), .ZN(n4317) );
NAND3_X2 U9873 ( .A1(n9977), .A2(n9978), .A3(n9979), .ZN(n4349) );
NAND3_X2 U9874 ( .A1(n9876), .A2(n9877), .A3(n9878), .ZN(n4381) );
NAND3_X2 U9875 ( .A1(n9677), .A2(n9678), .A3(n9679), .ZN(n4445) );
NAND3_X2 U9876 ( .A1(n9575), .A2(n9576), .A3(n9577), .ZN(n4477) );
NAND3_X2 U9877 ( .A1(n10764), .A2(n10765), .A3(n10766), .ZN(n4095) );
NAND3_X2 U9878 ( .A1(n10663), .A2(n10664), .A3(n10665), .ZN(n4127) );
NAND3_X2 U9879 ( .A1(n10564), .A2(n10565), .A3(n10566), .ZN(n4159) );
NAND3_X2 U9880 ( .A1(n10465), .A2(n10466), .A3(n10467), .ZN(n4191) );
NAND3_X2 U9881 ( .A1(n10366), .A2(n10367), .A3(n10368), .ZN(n4223) );
NAND3_X2 U9882 ( .A1(n10266), .A2(n10267), .A3(n10268), .ZN(n4255) );
NAND3_X2 U9883 ( .A1(n10073), .A2(n10074), .A3(n10075), .ZN(n4318) );
NAND3_X2 U9884 ( .A1(n9974), .A2(n9975), .A3(n9976), .ZN(n4350) );
NAND3_X2 U9885 ( .A1(n9873), .A2(n9874), .A3(n9875), .ZN(n4382) );
NAND3_X2 U9886 ( .A1(n9674), .A2(n9675), .A3(n9676), .ZN(n4446) );
NAND3_X2 U9887 ( .A1(n10761), .A2(n10762), .A3(n10763), .ZN(n4096) );
NAND3_X2 U9888 ( .A1(n10660), .A2(n10661), .A3(n10662), .ZN(n4128) );
NAND3_X2 U9889 ( .A1(n10561), .A2(n10562), .A3(n10563), .ZN(n4160) );
NAND3_X2 U9890 ( .A1(n10462), .A2(n10463), .A3(n10464), .ZN(n4192) );
NAND3_X2 U9891 ( .A1(n10363), .A2(n10364), .A3(n10365), .ZN(n4224) );
NAND3_X2 U9892 ( .A1(n10263), .A2(n10264), .A3(n10265), .ZN(n4256) );
NAND3_X2 U9893 ( .A1(n10070), .A2(n10071), .A3(n10072), .ZN(n4319) );
NAND3_X2 U9894 ( .A1(n9971), .A2(n9972), .A3(n9973), .ZN(n4351) );
NAND3_X2 U9895 ( .A1(n9870), .A2(n9871), .A3(n9872), .ZN(n4383) );
NAND3_X2 U9896 ( .A1(n9671), .A2(n9672), .A3(n9673), .ZN(n4447) );
NAND3_X2 U9897 ( .A1(n10758), .A2(n10759), .A3(n10760), .ZN(n4097) );
NAND3_X2 U9898 ( .A1(n10657), .A2(n10658), .A3(n10659), .ZN(n4129) );
NAND3_X2 U9899 ( .A1(n10558), .A2(n10559), .A3(n10560), .ZN(n4161) );
NAND3_X2 U9900 ( .A1(n10459), .A2(n10460), .A3(n10461), .ZN(n4193) );
NAND3_X2 U9901 ( .A1(n10360), .A2(n10361), .A3(n10362), .ZN(n4225) );
NAND3_X2 U9902 ( .A1(n10260), .A2(n10261), .A3(n10262), .ZN(n4257) );
NAND3_X2 U9903 ( .A1(n10067), .A2(n10068), .A3(n10069), .ZN(n4320) );
NAND3_X2 U9904 ( .A1(n9968), .A2(n9969), .A3(n9970), .ZN(n4352) );
NAND3_X2 U9905 ( .A1(n9867), .A2(n9868), .A3(n9869), .ZN(n4384) );
NAND3_X2 U9906 ( .A1(n9668), .A2(n9669), .A3(n9670), .ZN(n4448) );
NAND3_X2 U9907 ( .A1(n10755), .A2(n10756), .A3(n10757), .ZN(n4098) );
NAND3_X2 U9908 ( .A1(n10654), .A2(n10655), .A3(n10656), .ZN(n4130) );
NAND3_X2 U9909 ( .A1(n10555), .A2(n10556), .A3(n10557), .ZN(n4162) );
NAND3_X2 U9910 ( .A1(n10456), .A2(n10457), .A3(n10458), .ZN(n4194) );
NAND3_X2 U9911 ( .A1(n10357), .A2(n10358), .A3(n10359), .ZN(n4226) );
NAND3_X2 U9912 ( .A1(n10257), .A2(n10258), .A3(n10259), .ZN(n4258) );
NAND3_X2 U9913 ( .A1(n10064), .A2(n10065), .A3(n10066), .ZN(n4321) );
NAND3_X2 U9914 ( .A1(n9965), .A2(n9966), .A3(n9967), .ZN(n4353) );
NAND3_X2 U9915 ( .A1(n9864), .A2(n9865), .A3(n9866), .ZN(n4385) );
NAND3_X2 U9916 ( .A1(n9665), .A2(n9666), .A3(n9667), .ZN(n4449) );
NAND3_X2 U9917 ( .A1(n10752), .A2(n10753), .A3(n10754), .ZN(n4099) );
NAND3_X2 U9918 ( .A1(n10651), .A2(n10652), .A3(n10653), .ZN(n4131) );
NAND3_X2 U9919 ( .A1(n10552), .A2(n10553), .A3(n10554), .ZN(n4163) );
NAND3_X2 U9920 ( .A1(n10453), .A2(n10454), .A3(n10455), .ZN(n4195) );
NAND3_X2 U9921 ( .A1(n10354), .A2(n10355), .A3(n10356), .ZN(n4227) );
NAND3_X2 U9922 ( .A1(n10254), .A2(n10255), .A3(n10256), .ZN(n4259) );
NAND3_X2 U9923 ( .A1(n10061), .A2(n10062), .A3(n10063), .ZN(n4322) );
NAND3_X2 U9924 ( .A1(n9962), .A2(n9963), .A3(n9964), .ZN(n4354) );
NAND3_X2 U9925 ( .A1(n9861), .A2(n9862), .A3(n9863), .ZN(n4386) );
NAND3_X2 U9926 ( .A1(n9662), .A2(n9663), .A3(n9664), .ZN(n4450) );
NAND3_X2 U9927 ( .A1(n10749), .A2(n10750), .A3(n10751), .ZN(n4100) );
NAND3_X2 U9928 ( .A1(n10648), .A2(n10649), .A3(n10650), .ZN(n4132) );
NAND3_X2 U9929 ( .A1(n10549), .A2(n10550), .A3(n10551), .ZN(n4164) );
NAND3_X2 U9930 ( .A1(n10450), .A2(n10451), .A3(n10452), .ZN(n4196) );
NAND3_X2 U9931 ( .A1(n10351), .A2(n10352), .A3(n10353), .ZN(n4228) );
NAND3_X2 U9932 ( .A1(n10251), .A2(n10252), .A3(n10253), .ZN(n4260) );
NAND3_X2 U9933 ( .A1(n10058), .A2(n10059), .A3(n10060), .ZN(n4323) );
NAND3_X2 U9934 ( .A1(n9959), .A2(n9960), .A3(n9961), .ZN(n4355) );
NAND3_X2 U9935 ( .A1(n9858), .A2(n9859), .A3(n9860), .ZN(n4387) );
NAND3_X2 U9936 ( .A1(n9659), .A2(n9660), .A3(n9661), .ZN(n4451) );
NAND3_X2 U9937 ( .A1(n10746), .A2(n10747), .A3(n10748), .ZN(n4101) );
NAND3_X2 U9938 ( .A1(n10645), .A2(n10646), .A3(n10647), .ZN(n4133) );
NAND3_X2 U9939 ( .A1(n10546), .A2(n10547), .A3(n10548), .ZN(n4165) );
NAND3_X2 U9940 ( .A1(n10447), .A2(n10448), .A3(n10449), .ZN(n4197) );
NAND3_X2 U9941 ( .A1(n10348), .A2(n10349), .A3(n10350), .ZN(n4229) );
NAND3_X2 U9942 ( .A1(n10248), .A2(n10249), .A3(n10250), .ZN(n4261) );
NAND3_X2 U9943 ( .A1(n10055), .A2(n10056), .A3(n10057), .ZN(n4324) );
NAND3_X2 U9944 ( .A1(n9956), .A2(n9957), .A3(n9958), .ZN(n4356) );
NAND3_X2 U9945 ( .A1(n9855), .A2(n9856), .A3(n9857), .ZN(n4388) );
NAND3_X2 U9946 ( .A1(n9656), .A2(n9657), .A3(n9658), .ZN(n4452) );
NAND3_X2 U9947 ( .A1(n10743), .A2(n10744), .A3(n10745), .ZN(n4102) );
NAND3_X2 U9948 ( .A1(n10642), .A2(n10643), .A3(n10644), .ZN(n4134) );
NAND3_X2 U9949 ( .A1(n10543), .A2(n10544), .A3(n10545), .ZN(n4166) );
NAND3_X2 U9950 ( .A1(n10444), .A2(n10445), .A3(n10446), .ZN(n4198) );
NAND3_X2 U9951 ( .A1(n10345), .A2(n10346), .A3(n10347), .ZN(n4230) );
NAND3_X2 U9952 ( .A1(n10245), .A2(n10246), .A3(n10247), .ZN(n4262) );
NAND3_X2 U9953 ( .A1(n10052), .A2(n10053), .A3(n10054), .ZN(n4325) );
NAND3_X2 U9954 ( .A1(n9953), .A2(n9954), .A3(n9955), .ZN(n4357) );
NAND3_X2 U9955 ( .A1(n9852), .A2(n9853), .A3(n9854), .ZN(n4389) );
NAND3_X2 U9956 ( .A1(n9653), .A2(n9654), .A3(n9655), .ZN(n4453) );
NAND3_X2 U9957 ( .A1(n10740), .A2(n10741), .A3(n10742), .ZN(n4103) );
NAND3_X2 U9958 ( .A1(n10639), .A2(n10640), .A3(n10641), .ZN(n4135) );
NAND3_X2 U9959 ( .A1(n10540), .A2(n10541), .A3(n10542), .ZN(n4167) );
NAND3_X2 U9960 ( .A1(n10441), .A2(n10442), .A3(n10443), .ZN(n4199) );
NAND3_X2 U9961 ( .A1(n10342), .A2(n10343), .A3(n10344), .ZN(n4231) );
NAND3_X2 U9962 ( .A1(n10242), .A2(n10243), .A3(n10244), .ZN(n4263) );
NAND3_X2 U9963 ( .A1(n10049), .A2(n10050), .A3(n10051), .ZN(n4326) );
NAND3_X2 U9964 ( .A1(n9950), .A2(n9951), .A3(n9952), .ZN(n4358) );
NAND3_X2 U9965 ( .A1(n9849), .A2(n9850), .A3(n9851), .ZN(n4390) );
NAND3_X2 U9966 ( .A1(n9650), .A2(n9651), .A3(n9652), .ZN(n4454) );
NAND3_X2 U9967 ( .A1(n10737), .A2(n10738), .A3(n10739), .ZN(n4104) );
NAND3_X2 U9968 ( .A1(n10636), .A2(n10637), .A3(n10638), .ZN(n4136) );
NAND3_X2 U9969 ( .A1(n10537), .A2(n10538), .A3(n10539), .ZN(n4168) );
NAND3_X2 U9970 ( .A1(n10438), .A2(n10439), .A3(n10440), .ZN(n4200) );
NAND3_X2 U9971 ( .A1(n10339), .A2(n10340), .A3(n10341), .ZN(n4232) );
NAND3_X2 U9972 ( .A1(n10239), .A2(n10240), .A3(n10241), .ZN(n4264) );
NAND3_X2 U9973 ( .A1(n10046), .A2(n10047), .A3(n10048), .ZN(n4327) );
NAND3_X2 U9974 ( .A1(n9947), .A2(n9948), .A3(n9949), .ZN(n4359) );
NAND3_X2 U9975 ( .A1(n9846), .A2(n9847), .A3(n9848), .ZN(n4391) );
NAND3_X2 U9976 ( .A1(n9647), .A2(n9648), .A3(n9649), .ZN(n4455) );
NAND3_X2 U9977 ( .A1(n10734), .A2(n10735), .A3(n10736), .ZN(n4105) );
NAND3_X2 U9978 ( .A1(n10633), .A2(n10634), .A3(n10635), .ZN(n4137) );
NAND3_X2 U9979 ( .A1(n10534), .A2(n10535), .A3(n10536), .ZN(n4169) );
NAND3_X2 U9980 ( .A1(n10435), .A2(n10436), .A3(n10437), .ZN(n4201) );
NAND3_X2 U9981 ( .A1(n10336), .A2(n10337), .A3(n10338), .ZN(n4233) );
NAND3_X2 U9982 ( .A1(n10236), .A2(n10237), .A3(n10238), .ZN(n4265) );
NAND3_X2 U9983 ( .A1(n10043), .A2(n10044), .A3(n10045), .ZN(n4328) );
NAND3_X2 U9984 ( .A1(n9944), .A2(n9945), .A3(n9946), .ZN(n4360) );
NAND3_X2 U9985 ( .A1(n9843), .A2(n9844), .A3(n9845), .ZN(n4392) );
NAND3_X2 U9986 ( .A1(n9644), .A2(n9645), .A3(n9646), .ZN(n4456) );
NAND3_X2 U9987 ( .A1(n10731), .A2(n10732), .A3(n10733), .ZN(n4106) );
NAND3_X2 U9988 ( .A1(n10630), .A2(n10631), .A3(n10632), .ZN(n4138) );
NAND3_X2 U9989 ( .A1(n10531), .A2(n10532), .A3(n10533), .ZN(n4170) );
NAND3_X2 U9990 ( .A1(n10432), .A2(n10433), .A3(n10434), .ZN(n4202) );
NAND3_X2 U9991 ( .A1(n10333), .A2(n10334), .A3(n10335), .ZN(n4234) );
NAND3_X2 U9992 ( .A1(n10233), .A2(n10234), .A3(n10235), .ZN(n4266) );
NAND3_X2 U9993 ( .A1(n10040), .A2(n10041), .A3(n10042), .ZN(n4329) );
NAND3_X2 U9994 ( .A1(n9941), .A2(n9942), .A3(n9943), .ZN(n4361) );
NAND3_X2 U9995 ( .A1(n9840), .A2(n9841), .A3(n9842), .ZN(n4393) );
NAND3_X2 U9996 ( .A1(n9641), .A2(n9642), .A3(n9643), .ZN(n4457) );
NAND3_X2 U9997 ( .A1(n10728), .A2(n10729), .A3(n10730), .ZN(n4107) );
NAND3_X2 U9998 ( .A1(n10627), .A2(n10628), .A3(n10629), .ZN(n4139) );
NAND3_X2 U9999 ( .A1(n10528), .A2(n10529), .A3(n10530), .ZN(n4171) );
NAND3_X2 U10000 ( .A1(n10429), .A2(n10430), .A3(n10431), .ZN(n4203) );
NAND3_X2 U10001 ( .A1(n10330), .A2(n10331), .A3(n10332), .ZN(n4235) );
NAND3_X2 U10002 ( .A1(n10230), .A2(n10231), .A3(n10232), .ZN(n4267) );
NAND3_X2 U10003 ( .A1(n10037), .A2(n10038), .A3(n10039), .ZN(n4330) );
NAND3_X2 U10004 ( .A1(n9938), .A2(n9939), .A3(n9940), .ZN(n4362) );
NAND3_X2 U10005 ( .A1(n9837), .A2(n9838), .A3(n9839), .ZN(n4394) );
NAND3_X2 U10006 ( .A1(n9638), .A2(n9639), .A3(n9640), .ZN(n4458) );
NAND3_X2 U10007 ( .A1(n10725), .A2(n10726), .A3(n10727), .ZN(n4108) );
NAND3_X2 U10008 ( .A1(n10624), .A2(n10625), .A3(n10626), .ZN(n4140) );
NAND3_X2 U10009 ( .A1(n10525), .A2(n10526), .A3(n10527), .ZN(n4172) );
NAND3_X2 U10010 ( .A1(n10426), .A2(n10427), .A3(n10428), .ZN(n4204) );
NAND3_X2 U10011 ( .A1(n10327), .A2(n10328), .A3(n10329), .ZN(n4236) );
NAND3_X2 U10012 ( .A1(n10227), .A2(n10228), .A3(n10229), .ZN(n4268) );
NAND3_X2 U10013 ( .A1(n10034), .A2(n10035), .A3(n10036), .ZN(n4331) );
NAND3_X2 U10014 ( .A1(n9935), .A2(n9936), .A3(n9937), .ZN(n4363) );
NAND3_X2 U10015 ( .A1(n9834), .A2(n9835), .A3(n9836), .ZN(n4395) );
NAND3_X2 U10016 ( .A1(n9635), .A2(n9636), .A3(n9637), .ZN(n4459) );
NAND3_X2 U10017 ( .A1(n10722), .A2(n10723), .A3(n10724), .ZN(n4109) );
NAND3_X2 U10018 ( .A1(n10621), .A2(n10622), .A3(n10623), .ZN(n4141) );
NAND3_X2 U10019 ( .A1(n10522), .A2(n10523), .A3(n10524), .ZN(n4173) );
NAND3_X2 U10020 ( .A1(n10423), .A2(n10424), .A3(n10425), .ZN(n4205) );
NAND3_X2 U10021 ( .A1(n10324), .A2(n10325), .A3(n10326), .ZN(n4237) );
NAND3_X2 U10022 ( .A1(n10224), .A2(n10225), .A3(n10226), .ZN(n4269) );
NAND3_X2 U10023 ( .A1(n10031), .A2(n10032), .A3(n10033), .ZN(n4332) );
NAND3_X2 U10024 ( .A1(n9932), .A2(n9933), .A3(n9934), .ZN(n4364) );
NAND3_X2 U10025 ( .A1(n9831), .A2(n9832), .A3(n9833), .ZN(n4396) );
NAND3_X2 U10026 ( .A1(n9632), .A2(n9633), .A3(n9634), .ZN(n4460) );
NAND3_X2 U10027 ( .A1(n10719), .A2(n10720), .A3(n10721), .ZN(n4110) );
NAND3_X2 U10028 ( .A1(n10618), .A2(n10619), .A3(n10620), .ZN(n4142) );
NAND3_X2 U10029 ( .A1(n10519), .A2(n10520), .A3(n10521), .ZN(n4174) );
NAND3_X2 U10030 ( .A1(n10420), .A2(n10421), .A3(n10422), .ZN(n4206) );
NAND3_X2 U10031 ( .A1(n10321), .A2(n10322), .A3(n10323), .ZN(n4238) );
NAND3_X2 U10032 ( .A1(n10221), .A2(n10222), .A3(n10223), .ZN(n4270) );
NAND3_X2 U10033 ( .A1(n10028), .A2(n10029), .A3(n10030), .ZN(n4333) );
NAND3_X2 U10034 ( .A1(n9929), .A2(n9930), .A3(n9931), .ZN(n4365) );
NAND3_X2 U10035 ( .A1(n9828), .A2(n9829), .A3(n9830), .ZN(n4397) );
NAND3_X2 U10036 ( .A1(n9629), .A2(n9630), .A3(n9631), .ZN(n4461) );
NAND3_X2 U10037 ( .A1(n10716), .A2(n10717), .A3(n10718), .ZN(n4111) );
NAND3_X2 U10038 ( .A1(n10615), .A2(n10616), .A3(n10617), .ZN(n4143) );
NAND3_X2 U10039 ( .A1(n10516), .A2(n10517), .A3(n10518), .ZN(n4175) );
NAND3_X2 U10040 ( .A1(n10417), .A2(n10418), .A3(n10419), .ZN(n4207) );
NAND3_X2 U10041 ( .A1(n10318), .A2(n10319), .A3(n10320), .ZN(n4239) );
NAND3_X2 U10042 ( .A1(n10218), .A2(n10219), .A3(n10220), .ZN(n4271) );
NAND3_X2 U10043 ( .A1(n10025), .A2(n10026), .A3(n10027), .ZN(n4334) );
NAND3_X2 U10044 ( .A1(n9926), .A2(n9927), .A3(n9928), .ZN(n4366) );
NAND3_X2 U10045 ( .A1(n9825), .A2(n9826), .A3(n9827), .ZN(n4398) );
NAND3_X2 U10046 ( .A1(n9626), .A2(n9627), .A3(n9628), .ZN(n4462) );
NAND3_X2 U10047 ( .A1(n10711), .A2(n10712), .A3(n10713), .ZN(n4112) );
NAND3_X2 U10048 ( .A1(n10610), .A2(n10611), .A3(n10612), .ZN(n4144) );
NAND3_X2 U10049 ( .A1(n10511), .A2(n10512), .A3(n10513), .ZN(n4176) );
NAND3_X2 U10050 ( .A1(n10412), .A2(n10413), .A3(n10414), .ZN(n4208) );
NAND3_X2 U10051 ( .A1(n10313), .A2(n10314), .A3(n10315), .ZN(n4240) );
NAND3_X2 U10052 ( .A1(n10213), .A2(n10214), .A3(n10215), .ZN(n4272) );
NAND2_X4 U10053 ( .A1(n14267), .A2(n14279), .ZN(n14371) );
NAND2_X4 U10054 ( .A1(n14367), .A2(n14366), .ZN(n14929) );
NOR3_X4 U10055 ( .A1(n14254), .A2(n465), .A3(n14255), .ZN(n14262) );
XOR2_X1 U10056 ( .A(n13419), .B(n13077), .Z(n13420) );
NAND2_X1 U10057 ( .A1(n13071), .A2(n13076), .ZN(n13975) );
NAND3_X1 U10058 ( .A1(n13071), .A2(n14953), .A3(n14266), .ZN(n13982) );
NAND2_X1 U10059 ( .A1(n13197), .A2(n13081), .ZN(n14521) );
NAND2_X1 U10060 ( .A1(n13081), .A2(n13224), .ZN(n13761) );
NAND2_X1 U10061 ( .A1(n13203), .A2(n13081), .ZN(n13763) );
INV_X1 U10062 ( .A(n13081), .ZN(n14771) );
NAND2_X1 U10063 ( .A1(n13081), .A2(n14770), .ZN(n14311) );
NAND2_X1 U10064 ( .A1(round[0]), .A2(round[1]), .ZN(n13411) );
NAND3_X1 U10065 ( .A1(round[1]), .A2(n13398), .A3(n14067), .ZN(n14729) );
NAND4_X4 U10066 ( .A1(n14338), .A2(n14341), .A3(n14339), .A4(n14340), .ZN(SHA1_ft_BCD[3]) );
NAND3_X1 U10067 ( .A1(next_C[4]), .A2(SHA1_result[70]), .A3(n14334), .ZN(n14305) );
NAND2_X4 U10068 ( .A1(n13075), .A2(n13102), .ZN(n14334) );
NAND2_X1 U10069 ( .A1(n12983), .A2(n13208), .ZN(n13459) );
NAND2_X1 U10070 ( .A1(n13128), .A2(n13145), .ZN(n13409) );
NAND2_X1 U10071 ( .A1(n13087), .A2(n13145), .ZN(n14730) );
NAND2_X1 U10072 ( .A1(n13145), .A2(n12980), .ZN(n14707) );
NOR2_X1 U10073 ( .A1(n14359), .A2(n13143), .ZN(n14363) );
NAND3_X1 U10074 ( .A1(n14270), .A2(n14269), .A3(n14321), .ZN(n14271) );
NAND2_X1 U10075 ( .A1(next_A[26]), .A2(n13208), .ZN(n13506) );
NOR2_X1 U10076 ( .A1(n13146), .A2(n13027), .ZN(n13418) );
NAND2_X1 U10077 ( .A1(n13027), .A2(n13146), .ZN(n13419) );
NAND3_X1 U10078 ( .A1(round[5]), .A2(n13146), .A3(n14726), .ZN(n13968) );
NAND2_X1 U10079 ( .A1(n13146), .A2(n13069), .ZN(n13434) );
NAND2_X1 U10080 ( .A1(n13094), .A2(n13207), .ZN(n13567) );
NAND2_X1 U10081 ( .A1(next_A[22]), .A2(n13207), .ZN(n13553) );
NAND2_X1 U10082 ( .A1(n13106), .A2(n13207), .ZN(n13579) );
NAND2_X4 U10083 ( .A1(n14265), .A2(n14264), .ZN(SHA1_ft_BCD[10]) );
NAND2_X4 U10084 ( .A1(n13122), .A2(n14241), .ZN(SHA1_ft_BCD[12]) );
NAND3_X1 U10085 ( .A1(n463), .A2(n14368), .A3(n14239), .ZN(n14242) );
NAND2_X4 U10086 ( .A1(n14240), .A2(n14817), .ZN(n14241) );
NAND2_X1 U10087 ( .A1(n12989), .A2(n12980), .ZN(n14694) );
NAND2_X1 U10088 ( .A1(n13087), .A2(n12989), .ZN(n14714) );
INV_X16 U10089 ( .A(n13144), .ZN(n14688) );
INV_X16 U10090 ( .A(n14344), .ZN(n14368) );
INV_X4 U10091 ( .A(n11846), .ZN(n14955) );
INV_X4 U10092 ( .A(n14694), .ZN(n14691) );
INV_X4 U10093 ( .A(n13402), .ZN(n13424) );
NAND2_X2 U10094 ( .A1(n13424), .A2(n14688), .ZN(n13403) );
INV_X4 U10095 ( .A(n13403), .ZN(n13398) );
NAND2_X2 U10096 ( .A1(n12999), .A2(n13398), .ZN(n13998) );
INV_X4 U10097 ( .A(n13998), .ZN(n13397) );
NAND2_X2 U10098 ( .A1(n13397), .A2(n14953), .ZN(n14959) );
INV_X4 U10099 ( .A(n14959), .ZN(n14933) );
NAND2_X2 U10100 ( .A1(cmd_o[1]), .A2(n14933), .ZN(n13405) );
INV_X4 U10101 ( .A(n13411), .ZN(n13413) );
NAND2_X2 U10102 ( .A1(n13398), .A2(n13413), .ZN(n14699) );
INV_X4 U10103 ( .A(n14730), .ZN(n14726) );
NAND2_X2 U10104 ( .A1(n13025), .A2(n14726), .ZN(n14719) );
INV_X4 U10105 ( .A(n14714), .ZN(n14712) );
NAND2_X2 U10106 ( .A1(n14712), .A2(n13025), .ZN(n10212) );
INV_X4 U10107 ( .A(n10212), .ZN(n13400) );
INV_X4 U10108 ( .A(n14707), .ZN(n14705) );
NAND2_X2 U10109 ( .A1(n14705), .A2(n13025), .ZN(n10609) );
INV_X4 U10110 ( .A(n10609), .ZN(n13399) );
INV_X4 U10111 ( .A(n14693), .ZN(n14722) );
NOR3_X2 U10112 ( .A1(n13400), .A2(n13399), .A3(n14722), .ZN(n13401) );
NAND2_X2 U10113 ( .A1(n13069), .A2(n13402), .ZN(n14733) );
NAND2_X2 U10114 ( .A1(n14733), .A2(n13403), .ZN(n14687) );
NAND2_X2 U10115 ( .A1(n13026), .A2(n14687), .ZN(n13404) );
NAND2_X2 U10116 ( .A1(n13404), .A2(n14953), .ZN(n13436) );
NAND2_X2 U10117 ( .A1(n13405), .A2(n13436), .ZN(n13407) );
INV_X4 U10118 ( .A(n13407), .ZN(n13421) );
NOR2_X2 U10119 ( .A1(n13421), .A2(n14067), .ZN(n13406) );
MUX2_X2 U10120 ( .A(n13406), .B(n13128), .S(round[1]), .Z(N1715) );
MUX2_X2 U10121 ( .A(n13413), .B(n13093), .S(n13145), .Z(n13408) );
NAND2_X2 U10122 ( .A1(n13408), .A2(n13407), .ZN(n13410) );
NAND2_X2 U10123 ( .A1(n13410), .A2(n13409), .ZN(N1716) );
NOR2_X2 U10124 ( .A1(n13087), .A2(n13412), .ZN(n13414) );
NOR3_X2 U10125 ( .A1(n13414), .A2(n13421), .A3(n13027), .ZN(N1717) );
NOR2_X2 U10126 ( .A1(n13069), .A2(n13415), .ZN(n13416) );
NOR2_X2 U10127 ( .A1(n13421), .A2(n13416), .ZN(N1720) );
INV_X4 U10128 ( .A(n13419), .ZN(n13417) );
NOR3_X2 U10129 ( .A1(n13418), .A2(n13421), .A3(n13417), .ZN(N1718) );
NOR2_X2 U10130 ( .A1(n13421), .A2(n13420), .ZN(N1719) );
NAND2_X2 U10131 ( .A1(n12999), .A2(n13424), .ZN(n13422) );
NAND2_X2 U10132 ( .A1(n13422), .A2(n14688), .ZN(n13428) );
NAND2_X2 U10133 ( .A1(n345), .A2(n14688), .ZN(n13423) );
NAND2_X2 U10134 ( .A1(n13424), .A2(n13423), .ZN(n13425) );
NAND3_X2 U10135 ( .A1(n13428), .A2(n14953), .A3(n13425), .ZN(n14000) );
NAND2_X2 U10136 ( .A1(n13156), .A2(n13426), .ZN(n13437) );
NAND2_X2 U10137 ( .A1(n14933), .A2(cmd_o[2]), .ZN(n13427) );
NAND2_X2 U10138 ( .A1(next_A[0]), .A2(n13206), .ZN(n13433) );
NAND3_X2 U10139 ( .A1(n13429), .A2(n13428), .A3(n12995), .ZN(n13430) );
NAND2_X2 U10140 ( .A1(N852), .A2(n13180), .ZN(n13432) );
NAND2_X2 U10141 ( .A1(n13214), .A2(SHA1_result_128), .ZN(n13431) );
NAND4_X2 U10142 ( .A1(n13433), .A2(n13432), .A3(n13431), .A4(n13185), .ZN(n4016) );
INV_X4 U10143 ( .A(n13434), .ZN(n13435) );
NAND2_X2 U10144 ( .A1(N884), .A2(n13166), .ZN(n13441) );
NAND2_X2 U10145 ( .A1(next_C[30]), .A2(n13150), .ZN(n13440) );
INV_X4 U10146 ( .A(n13436), .ZN(n13438) );
NAND2_X2 U10147 ( .A1(n13172), .A2(SHA1_result_128), .ZN(n13439) );
NAND4_X2 U10148 ( .A1(n13441), .A2(n13151), .A3(n13440), .A4(n13439), .ZN(n3952) );
NAND2_X2 U10149 ( .A1(n13200), .A2(next_C[30]), .ZN(n13444) );
NAND2_X2 U10150 ( .A1(N946), .A2(n13213), .ZN(n13443) );
NAND2_X2 U10151 ( .A1(n13222), .A2(SHA1_result[94]), .ZN(n13442) );
NAND3_X2 U10152 ( .A1(n13444), .A2(n13443), .A3(n13442), .ZN(n3890) );
NAND2_X2 U10153 ( .A1(n13200), .A2(SHA1_result[94]), .ZN(n13447) );
NAND2_X2 U10154 ( .A1(N978), .A2(n13213), .ZN(n13446) );
NAND2_X2 U10155 ( .A1(n13224), .A2(SHA1_result[62]), .ZN(n13445) );
NAND3_X2 U10156 ( .A1(n13447), .A2(n13446), .A3(n13445), .ZN(n3858) );
NAND2_X2 U10157 ( .A1(N915), .A2(n13166), .ZN(n13450) );
NAND2_X2 U10158 ( .A1(next_C[29]), .A2(n13150), .ZN(n13449) );
NAND2_X2 U10159 ( .A1(n13172), .A2(n14464), .ZN(n13448) );
NAND4_X2 U10160 ( .A1(n13450), .A2(n13153), .A3(n13449), .A4(n13448), .ZN(n3921) );
NAND2_X2 U10161 ( .A1(n13200), .A2(next_C[29]), .ZN(n13453) );
NAND2_X2 U10162 ( .A1(N945), .A2(n13213), .ZN(n13452) );
NAND2_X2 U10163 ( .A1(n13224), .A2(SHA1_result[93]), .ZN(n13451) );
NAND3_X2 U10164 ( .A1(n13453), .A2(n13452), .A3(n13451), .ZN(n3891) );
NAND2_X2 U10165 ( .A1(n13200), .A2(SHA1_result[93]), .ZN(n13456) );
NAND2_X2 U10166 ( .A1(N977), .A2(n13213), .ZN(n13455) );
NAND2_X2 U10167 ( .A1(n13223), .A2(SHA1_result[61]), .ZN(n13454) );
NAND3_X2 U10168 ( .A1(n13456), .A2(n13455), .A3(n13454), .ZN(n3859) );
NAND2_X2 U10169 ( .A1(n13223), .A2(n14382), .ZN(n13458) );
NAND2_X2 U10170 ( .A1(N882), .A2(n13178), .ZN(n13457) );
NAND4_X2 U10171 ( .A1(n13457), .A2(n13184), .A3(n13458), .A4(n13459), .ZN(n3986) );
NAND2_X2 U10172 ( .A1(n13172), .A2(n14382), .ZN(n13462) );
NAND2_X2 U10173 ( .A1(N914), .A2(n13166), .ZN(n13461) );
NAND2_X2 U10174 ( .A1(next_C[28]), .A2(n13149), .ZN(n13460) );
NAND4_X2 U10175 ( .A1(n13462), .A2(n13461), .A3(n13460), .A4(n13151), .ZN(n3922) );
NAND2_X2 U10176 ( .A1(N944), .A2(n13178), .ZN(n13465) );
NAND2_X2 U10177 ( .A1(n13223), .A2(SHA1_result[92]), .ZN(n13464) );
NAND2_X2 U10178 ( .A1(n13200), .A2(next_C[28]), .ZN(n13463) );
NAND4_X2 U10179 ( .A1(n13465), .A2(n13185), .A3(n13464), .A4(n13463), .ZN(n3892) );
NAND2_X2 U10180 ( .A1(N976), .A2(n13178), .ZN(n13468) );
NAND2_X2 U10181 ( .A1(n13223), .A2(SHA1_result[60]), .ZN(n13467) );
NAND2_X2 U10182 ( .A1(n13200), .A2(SHA1_result[92]), .ZN(n13466) );
NAND4_X2 U10183 ( .A1(n13468), .A2(n13185), .A3(n13467), .A4(n13466), .ZN(n3860) );
NAND2_X2 U10184 ( .A1(N881), .A2(n13178), .ZN(n13470) );
NAND2_X2 U10185 ( .A1(n13223), .A2(n14385), .ZN(n13469) );
NAND4_X2 U10186 ( .A1(n13470), .A2(n13471), .A3(n13185), .A4(n13469), .ZN(n3987) );
NAND2_X2 U10187 ( .A1(N913), .A2(n13166), .ZN(n13474) );
NAND2_X2 U10188 ( .A1(next_C[27]), .A2(n13149), .ZN(n13473) );
NAND2_X2 U10189 ( .A1(n13172), .A2(n14385), .ZN(n13472) );
NAND4_X2 U10190 ( .A1(n13474), .A2(n13153), .A3(n13473), .A4(n13472), .ZN(n3923) );
NAND2_X2 U10191 ( .A1(N943), .A2(n13178), .ZN(n13477) );
NAND2_X2 U10192 ( .A1(n13223), .A2(SHA1_result[91]), .ZN(n13476) );
NAND2_X2 U10193 ( .A1(n13200), .A2(next_C[27]), .ZN(n13475) );
NAND4_X2 U10194 ( .A1(n13477), .A2(n13185), .A3(n13476), .A4(n13475), .ZN(n3893) );
NAND2_X2 U10195 ( .A1(n13200), .A2(SHA1_result[91]), .ZN(n13480) );
NAND2_X2 U10196 ( .A1(N975), .A2(n13213), .ZN(n13479) );
NAND2_X2 U10197 ( .A1(n13223), .A2(SHA1_result[59]), .ZN(n13478) );
NAND3_X2 U10198 ( .A1(n13480), .A2(n13479), .A3(n13478), .ZN(n3861) );
NAND2_X2 U10199 ( .A1(n13223), .A2(n14388), .ZN(n13481) );
NAND2_X2 U10200 ( .A1(N912), .A2(n13166), .ZN(n13486) );
NAND2_X2 U10201 ( .A1(next_C[26]), .A2(n13224), .ZN(n13485) );
NAND2_X2 U10202 ( .A1(n13172), .A2(n14388), .ZN(n13484) );
NAND3_X2 U10203 ( .A1(n13486), .A2(n13485), .A3(n13484), .ZN(n3924) );
NAND2_X2 U10204 ( .A1(n13200), .A2(next_C[26]), .ZN(n13489) );
NAND2_X2 U10205 ( .A1(N942), .A2(n13213), .ZN(n13488) );
NAND2_X2 U10206 ( .A1(n13223), .A2(SHA1_result[90]), .ZN(n13487) );
NAND3_X2 U10207 ( .A1(n13489), .A2(n13488), .A3(n13487), .ZN(n3894) );
NAND2_X2 U10208 ( .A1(n13201), .A2(SHA1_result[90]), .ZN(n13492) );
NAND2_X2 U10209 ( .A1(N974), .A2(n13213), .ZN(n13491) );
NAND2_X2 U10210 ( .A1(n13222), .A2(SHA1_result[58]), .ZN(n13490) );
NAND3_X2 U10211 ( .A1(n13492), .A2(n13491), .A3(n13490), .ZN(n3862) );
NAND2_X2 U10212 ( .A1(N911), .A2(n13166), .ZN(n13498) );
NAND2_X2 U10213 ( .A1(next_C[25]), .A2(n13149), .ZN(n13497) );
NAND2_X2 U10214 ( .A1(n13172), .A2(n14391), .ZN(n13496) );
NAND4_X2 U10215 ( .A1(n13498), .A2(n13153), .A3(n13497), .A4(n13496), .ZN(n3925) );
NAND2_X2 U10216 ( .A1(n13201), .A2(next_C[25]), .ZN(n13501) );
NAND2_X2 U10217 ( .A1(N941), .A2(n13212), .ZN(n13500) );
NAND2_X2 U10218 ( .A1(n13222), .A2(SHA1_result[89]), .ZN(n13499) );
NAND3_X2 U10219 ( .A1(n13501), .A2(n13500), .A3(n13499), .ZN(n3895) );
NAND2_X2 U10220 ( .A1(n13201), .A2(SHA1_result[89]), .ZN(n13504) );
NAND2_X2 U10221 ( .A1(N973), .A2(n13212), .ZN(n13503) );
NAND2_X2 U10222 ( .A1(n13223), .A2(SHA1_result[57]), .ZN(n13502) );
NAND3_X2 U10223 ( .A1(n13504), .A2(n13503), .A3(n13502), .ZN(n3863) );
NAND2_X2 U10224 ( .A1(n13222), .A2(n14394), .ZN(n13507) );
NAND2_X2 U10225 ( .A1(N910), .A2(n13166), .ZN(n13510) );
NAND2_X2 U10226 ( .A1(next_C[24]), .A2(n13149), .ZN(n13509) );
NAND2_X2 U10227 ( .A1(n13172), .A2(n14394), .ZN(n13508) );
NAND4_X2 U10228 ( .A1(n13510), .A2(n13153), .A3(n13509), .A4(n13508), .ZN(n3926) );
NAND2_X2 U10229 ( .A1(n13201), .A2(next_C[24]), .ZN(n13513) );
NAND2_X2 U10230 ( .A1(N940), .A2(n13212), .ZN(n13512) );
NAND2_X2 U10231 ( .A1(n13223), .A2(SHA1_result[88]), .ZN(n13511) );
NAND3_X2 U10232 ( .A1(n13513), .A2(n13512), .A3(n13511), .ZN(n3896) );
NAND2_X2 U10233 ( .A1(n13201), .A2(SHA1_result[88]), .ZN(n13516) );
NAND2_X2 U10234 ( .A1(N972), .A2(n13212), .ZN(n13515) );
NAND2_X2 U10235 ( .A1(n13222), .A2(SHA1_result[56]), .ZN(n13514) );
NAND3_X2 U10236 ( .A1(n13516), .A2(n13515), .A3(n13514), .ZN(n3864) );
NAND2_X2 U10237 ( .A1(N877), .A2(n13178), .ZN(n13519) );
NAND2_X2 U10238 ( .A1(n13222), .A2(n14397), .ZN(n13518) );
NAND4_X2 U10239 ( .A1(n13519), .A2(n13185), .A3(n13518), .A4(n13517), .ZN(n3991) );
NAND2_X2 U10240 ( .A1(N909), .A2(n13166), .ZN(n13522) );
NAND2_X2 U10241 ( .A1(next_C[23]), .A2(n13149), .ZN(n13521) );
NAND2_X2 U10242 ( .A1(n13172), .A2(n14397), .ZN(n13520) );
NAND4_X2 U10243 ( .A1(n13522), .A2(n13153), .A3(n13521), .A4(n13520), .ZN(n3927) );
NAND2_X2 U10244 ( .A1(N939), .A2(n13178), .ZN(n13525) );
NAND2_X2 U10245 ( .A1(n13222), .A2(SHA1_result[87]), .ZN(n13524) );
NAND2_X2 U10246 ( .A1(n13201), .A2(next_C[23]), .ZN(n13523) );
NAND4_X2 U10247 ( .A1(n13525), .A2(n13185), .A3(n13524), .A4(n13523), .ZN(n3897) );
NAND2_X2 U10248 ( .A1(n13201), .A2(SHA1_result[87]), .ZN(n13528) );
NAND2_X2 U10249 ( .A1(N971), .A2(n13212), .ZN(n13527) );
NAND2_X2 U10250 ( .A1(n13222), .A2(SHA1_result[55]), .ZN(n13526) );
NAND3_X2 U10251 ( .A1(n13528), .A2(n13527), .A3(n13526), .ZN(n3865) );
NAND2_X2 U10252 ( .A1(n13221), .A2(n14400), .ZN(n13530) );
NAND2_X2 U10253 ( .A1(N876), .A2(n13179), .ZN(n13529) );
NAND2_X2 U10254 ( .A1(N908), .A2(n13166), .ZN(n13534) );
NAND2_X2 U10255 ( .A1(next_C[22]), .A2(n13149), .ZN(n13533) );
NAND2_X2 U10256 ( .A1(n13172), .A2(n14400), .ZN(n13532) );
NAND4_X2 U10257 ( .A1(n13534), .A2(n13153), .A3(n13533), .A4(n13532), .ZN(n3928) );
NAND2_X2 U10258 ( .A1(n13201), .A2(next_C[22]), .ZN(n13537) );
NAND2_X2 U10259 ( .A1(N938), .A2(n13212), .ZN(n13536) );
NAND2_X2 U10260 ( .A1(n13221), .A2(SHA1_result[86]), .ZN(n13535) );
NAND3_X2 U10261 ( .A1(n13537), .A2(n13536), .A3(n13535), .ZN(n3898) );
NAND2_X2 U10262 ( .A1(n13202), .A2(SHA1_result[86]), .ZN(n13540) );
NAND2_X2 U10263 ( .A1(N970), .A2(n13212), .ZN(n13539) );
NAND2_X2 U10264 ( .A1(n13222), .A2(n14681), .ZN(n13538) );
NAND3_X2 U10265 ( .A1(n13540), .A2(n13539), .A3(n13538), .ZN(n3866) );
NAND2_X2 U10266 ( .A1(n13221), .A2(SHA1_result_151), .ZN(n13541) );
NAND2_X2 U10267 ( .A1(N907), .A2(n13166), .ZN(n13546) );
NAND2_X2 U10268 ( .A1(next_C[21]), .A2(n13149), .ZN(n13545) );
NAND2_X2 U10269 ( .A1(n13172), .A2(SHA1_result_151), .ZN(n13544) );
NAND4_X2 U10270 ( .A1(n13546), .A2(n13153), .A3(n13545), .A4(n13544), .ZN(n3929) );
NAND2_X2 U10271 ( .A1(N937), .A2(n13179), .ZN(n13549) );
NAND2_X2 U10272 ( .A1(n13219), .A2(SHA1_result[85]), .ZN(n13548) );
NAND2_X2 U10273 ( .A1(n13202), .A2(next_C[21]), .ZN(n13547) );
NAND4_X2 U10274 ( .A1(n13549), .A2(n13185), .A3(n13548), .A4(n13547), .ZN(n3899) );
NAND2_X2 U10275 ( .A1(N969), .A2(n13179), .ZN(n13552) );
INV_X4 U10276 ( .A(n422), .ZN(n14682) );
NAND2_X2 U10277 ( .A1(n13222), .A2(n14682), .ZN(n13551) );
NAND2_X2 U10278 ( .A1(n13202), .A2(SHA1_result[85]), .ZN(n13550) );
NAND4_X2 U10279 ( .A1(n13552), .A2(n13184), .A3(n13551), .A4(n13550), .ZN(n3867) );
NAND2_X2 U10280 ( .A1(N874), .A2(n13179), .ZN(n13555) );
NAND2_X2 U10281 ( .A1(n13221), .A2(n14405), .ZN(n13554) );
NAND4_X2 U10282 ( .A1(n13555), .A2(n13184), .A3(n13554), .A4(n13553), .ZN(n3994) );
NAND2_X2 U10283 ( .A1(N906), .A2(n13166), .ZN(n13558) );
NAND2_X2 U10284 ( .A1(next_C[20]), .A2(n13149), .ZN(n13557) );
NAND2_X2 U10285 ( .A1(n13172), .A2(n14405), .ZN(n13556) );
NAND4_X2 U10286 ( .A1(n13558), .A2(n13153), .A3(n13557), .A4(n13556), .ZN(n3930) );
NAND2_X2 U10287 ( .A1(N936), .A2(n13179), .ZN(n13561) );
NAND2_X2 U10288 ( .A1(n13221), .A2(SHA1_result[84]), .ZN(n13560) );
NAND2_X2 U10289 ( .A1(n13201), .A2(next_C[20]), .ZN(n13559) );
NAND4_X2 U10290 ( .A1(n13561), .A2(n13184), .A3(n13560), .A4(n13559), .ZN(n3900) );
NAND2_X2 U10291 ( .A1(N968), .A2(n13179), .ZN(n13564) );
INV_X4 U10292 ( .A(n423), .ZN(n14868) );
NAND2_X2 U10293 ( .A1(n13221), .A2(n14868), .ZN(n13563) );
NAND2_X2 U10294 ( .A1(n13202), .A2(SHA1_result[84]), .ZN(n13562) );
NAND4_X2 U10295 ( .A1(n13564), .A2(n13184), .A3(n13563), .A4(n13562), .ZN(n3868) );
NAND2_X2 U10296 ( .A1(n13221), .A2(n14408), .ZN(n13566) );
NAND2_X2 U10297 ( .A1(N873), .A2(n13212), .ZN(n13565) );
NAND3_X2 U10298 ( .A1(n13565), .A2(n13566), .A3(n13567), .ZN(n3995) );
NAND2_X2 U10299 ( .A1(N905), .A2(n13167), .ZN(n13570) );
NAND2_X2 U10300 ( .A1(next_C[19]), .A2(n13224), .ZN(n13569) );
NAND2_X2 U10301 ( .A1(n13173), .A2(n14408), .ZN(n13568) );
NAND3_X2 U10302 ( .A1(n13570), .A2(n13569), .A3(n13568), .ZN(n3931) );
NAND2_X2 U10303 ( .A1(N935), .A2(n13179), .ZN(n13573) );
NAND2_X2 U10304 ( .A1(n13221), .A2(SHA1_result[83]), .ZN(n13572) );
NAND2_X2 U10305 ( .A1(n13202), .A2(next_C[19]), .ZN(n13571) );
NAND4_X2 U10306 ( .A1(n13573), .A2(n13184), .A3(n13572), .A4(n13571), .ZN(n3901) );
NAND2_X2 U10307 ( .A1(n13202), .A2(SHA1_result[83]), .ZN(n13576) );
NAND2_X2 U10308 ( .A1(N967), .A2(n13212), .ZN(n13575) );
NAND2_X2 U10309 ( .A1(n13221), .A2(SHA1_result[51]), .ZN(n13574) );
NAND3_X2 U10310 ( .A1(n13576), .A2(n13575), .A3(n13574), .ZN(n3869) );
NAND2_X2 U10311 ( .A1(N872), .A2(n13211), .ZN(n13578) );
NAND2_X2 U10312 ( .A1(n13221), .A2(SHA1_result_148), .ZN(n13577) );
NAND3_X2 U10313 ( .A1(n13578), .A2(n13579), .A3(n13577), .ZN(n3996) );
NAND2_X2 U10314 ( .A1(N904), .A2(n13167), .ZN(n13582) );
NAND2_X2 U10315 ( .A1(next_C[18]), .A2(n13224), .ZN(n13581) );
NAND2_X2 U10316 ( .A1(n13173), .A2(SHA1_result_148), .ZN(n13580) );
NAND3_X2 U10317 ( .A1(n13582), .A2(n13581), .A3(n13580), .ZN(n3932) );
NAND2_X2 U10318 ( .A1(n13202), .A2(next_C[18]), .ZN(n13585) );
NAND2_X2 U10319 ( .A1(N934), .A2(n13211), .ZN(n13584) );
NAND2_X2 U10320 ( .A1(n13221), .A2(SHA1_result[82]), .ZN(n13583) );
NAND3_X2 U10321 ( .A1(n13585), .A2(n13584), .A3(n13583), .ZN(n3902) );
NAND2_X2 U10322 ( .A1(n13203), .A2(SHA1_result[82]), .ZN(n13588) );
NAND2_X2 U10323 ( .A1(N966), .A2(n13211), .ZN(n13587) );
NAND2_X2 U10324 ( .A1(n13220), .A2(SHA1_result[50]), .ZN(n13586) );
NAND3_X2 U10325 ( .A1(n13588), .A2(n13587), .A3(n13586), .ZN(n3870) );
NAND2_X2 U10326 ( .A1(N871), .A2(n13211), .ZN(n13590) );
NAND2_X2 U10327 ( .A1(n13220), .A2(n14413), .ZN(n13589) );
NAND2_X2 U10328 ( .A1(N903), .A2(n13167), .ZN(n13594) );
NAND2_X2 U10329 ( .A1(next_C[17]), .A2(n13149), .ZN(n13593) );
NAND2_X2 U10330 ( .A1(n13173), .A2(n14413), .ZN(n13592) );
NAND4_X2 U10331 ( .A1(n13594), .A2(n13153), .A3(n13593), .A4(n13592), .ZN(n3933) );
NAND2_X2 U10332 ( .A1(N933), .A2(n13179), .ZN(n13597) );
NAND2_X2 U10333 ( .A1(n13220), .A2(SHA1_result[81]), .ZN(n13596) );
NAND2_X2 U10334 ( .A1(n13203), .A2(next_C[17]), .ZN(n13595) );
NAND4_X2 U10335 ( .A1(n13597), .A2(n13184), .A3(n13596), .A4(n13595), .ZN(n3903) );
NAND2_X2 U10336 ( .A1(N965), .A2(n13179), .ZN(n13600) );
NAND2_X2 U10337 ( .A1(n13220), .A2(SHA1_result[49]), .ZN(n13599) );
NAND2_X2 U10338 ( .A1(n13200), .A2(SHA1_result[81]), .ZN(n13598) );
NAND4_X2 U10339 ( .A1(n13600), .A2(n13184), .A3(n13599), .A4(n13598), .ZN(n3871) );
NAND2_X2 U10340 ( .A1(N870), .A2(n13179), .ZN(n13603) );
NAND2_X2 U10341 ( .A1(n13220), .A2(n14416), .ZN(n13602) );
NAND4_X2 U10342 ( .A1(n13603), .A2(n13184), .A3(n13602), .A4(n13601), .ZN(n3998) );
NAND2_X2 U10343 ( .A1(N902), .A2(n13167), .ZN(n13606) );
NAND2_X2 U10344 ( .A1(next_C[16]), .A2(n13149), .ZN(n13605) );
NAND2_X2 U10345 ( .A1(n13173), .A2(n14416), .ZN(n13604) );
NAND4_X2 U10346 ( .A1(n13606), .A2(n13153), .A3(n13605), .A4(n13604), .ZN(n3934) );
NAND2_X2 U10347 ( .A1(n13202), .A2(next_C[16]), .ZN(n13609) );
NAND2_X2 U10348 ( .A1(N932), .A2(n13211), .ZN(n13608) );
NAND2_X2 U10349 ( .A1(n13220), .A2(SHA1_result[80]), .ZN(n13607) );
NAND3_X2 U10350 ( .A1(n13609), .A2(n13608), .A3(n13607), .ZN(n3904) );
NAND2_X2 U10351 ( .A1(n13203), .A2(SHA1_result[80]), .ZN(n13612) );
NAND2_X2 U10352 ( .A1(N964), .A2(n13211), .ZN(n13611) );
NAND2_X2 U10353 ( .A1(n13220), .A2(SHA1_result[48]), .ZN(n13610) );
NAND3_X2 U10354 ( .A1(n13612), .A2(n13611), .A3(n13610), .ZN(n3872) );
NAND2_X2 U10355 ( .A1(n13220), .A2(n14419), .ZN(n13613) );
NAND2_X2 U10356 ( .A1(N901), .A2(n13167), .ZN(n13618) );
NAND2_X2 U10357 ( .A1(next_C[15]), .A2(n13224), .ZN(n13617) );
NAND2_X2 U10358 ( .A1(n13173), .A2(n14419), .ZN(n13616) );
NAND3_X2 U10359 ( .A1(n13618), .A2(n13617), .A3(n13616), .ZN(n3935) );
NAND2_X2 U10360 ( .A1(N931), .A2(n13179), .ZN(n13621) );
NAND2_X2 U10361 ( .A1(n13220), .A2(SHA1_result[79]), .ZN(n13620) );
NAND2_X2 U10362 ( .A1(n13203), .A2(next_C[15]), .ZN(n13619) );
NAND4_X2 U10363 ( .A1(n13621), .A2(n13184), .A3(n13620), .A4(n13619), .ZN(n3905) );
NAND2_X2 U10364 ( .A1(n13203), .A2(SHA1_result[79]), .ZN(n13624) );
NAND2_X2 U10365 ( .A1(N963), .A2(n13211), .ZN(n13623) );
NAND2_X2 U10366 ( .A1(n13220), .A2(SHA1_result[47]), .ZN(n13622) );
NAND3_X2 U10367 ( .A1(n13624), .A2(n13623), .A3(n13622), .ZN(n3873) );
NAND2_X2 U10368 ( .A1(N868), .A2(n13179), .ZN(n13627) );
NAND2_X2 U10369 ( .A1(n13219), .A2(n14422), .ZN(n13626) );
NAND2_X2 U10370 ( .A1(n13108), .A2(n13207), .ZN(n13625) );
NAND4_X2 U10371 ( .A1(n13627), .A2(n13184), .A3(n13626), .A4(n13625), .ZN(n4000) );
NAND2_X2 U10372 ( .A1(N900), .A2(n13167), .ZN(n13630) );
NAND2_X2 U10373 ( .A1(next_C[14]), .A2(n13149), .ZN(n13629) );
NAND2_X2 U10374 ( .A1(n13173), .A2(n14422), .ZN(n13628) );
NAND4_X2 U10375 ( .A1(n13630), .A2(n13153), .A3(n13629), .A4(n13628), .ZN(n3936) );
NAND2_X2 U10376 ( .A1(N930), .A2(n13180), .ZN(n13633) );
NAND2_X2 U10377 ( .A1(n13220), .A2(SHA1_result[78]), .ZN(n13632) );
NAND2_X2 U10378 ( .A1(n13203), .A2(next_C[14]), .ZN(n13631) );
NAND4_X2 U10379 ( .A1(n13633), .A2(n13184), .A3(n13632), .A4(n13631), .ZN(n3906) );
NAND2_X2 U10380 ( .A1(N962), .A2(n13180), .ZN(n13636) );
NAND2_X2 U10381 ( .A1(n13219), .A2(n14830), .ZN(n13635) );
NAND2_X2 U10382 ( .A1(n13204), .A2(SHA1_result[78]), .ZN(n13634) );
NAND4_X2 U10383 ( .A1(n13636), .A2(n13184), .A3(n13635), .A4(n13634), .ZN(n3874) );
NAND2_X2 U10384 ( .A1(N867), .A2(n13211), .ZN(n13638) );
NAND2_X2 U10385 ( .A1(n13219), .A2(n14425), .ZN(n13637) );
NAND3_X2 U10386 ( .A1(n13639), .A2(n13638), .A3(n13637), .ZN(n4001) );
NAND2_X2 U10387 ( .A1(N899), .A2(n13167), .ZN(n13642) );
NAND2_X2 U10388 ( .A1(next_C[13]), .A2(n13149), .ZN(n13641) );
NAND2_X2 U10389 ( .A1(n13173), .A2(n14425), .ZN(n13640) );
NAND4_X2 U10390 ( .A1(n13642), .A2(n13153), .A3(n13641), .A4(n13640), .ZN(n3937) );
NAND2_X2 U10391 ( .A1(n13204), .A2(next_C[13]), .ZN(n13645) );
NAND2_X2 U10392 ( .A1(N929), .A2(n13211), .ZN(n13644) );
NAND2_X2 U10393 ( .A1(n13219), .A2(SHA1_result[77]), .ZN(n13643) );
NAND3_X2 U10394 ( .A1(n13645), .A2(n13644), .A3(n13643), .ZN(n3907) );
NAND2_X2 U10395 ( .A1(n13204), .A2(SHA1_result[77]), .ZN(n13648) );
NAND2_X2 U10396 ( .A1(N961), .A2(n13211), .ZN(n13647) );
NAND2_X2 U10397 ( .A1(n13219), .A2(SHA1_result[45]), .ZN(n13646) );
NAND3_X2 U10398 ( .A1(n13648), .A2(n13647), .A3(n13646), .ZN(n3875) );
NAND2_X2 U10399 ( .A1(N866), .A2(n13210), .ZN(n13650) );
NAND2_X2 U10400 ( .A1(n13219), .A2(n14428), .ZN(n13649) );
NAND3_X2 U10401 ( .A1(n13651), .A2(n13650), .A3(n13649), .ZN(n4002) );
NAND2_X2 U10402 ( .A1(N898), .A2(n13167), .ZN(n13654) );
NAND2_X2 U10403 ( .A1(next_C[12]), .A2(n13224), .ZN(n13653) );
NAND2_X2 U10404 ( .A1(n13173), .A2(n14428), .ZN(n13652) );
NAND3_X2 U10405 ( .A1(n13654), .A2(n13653), .A3(n13652), .ZN(n3938) );
NAND2_X2 U10406 ( .A1(N928), .A2(n13180), .ZN(n13657) );
NAND2_X2 U10407 ( .A1(n13219), .A2(SHA1_result[76]), .ZN(n13656) );
NAND2_X2 U10408 ( .A1(n13203), .A2(next_C[12]), .ZN(n13655) );
NAND4_X2 U10409 ( .A1(n13657), .A2(n13183), .A3(n13656), .A4(n13655), .ZN(n3908) );
NAND2_X2 U10410 ( .A1(N960), .A2(n13180), .ZN(n13660) );
NAND2_X2 U10411 ( .A1(n13219), .A2(n14817), .ZN(n13659) );
NAND2_X2 U10412 ( .A1(n13204), .A2(SHA1_result[76]), .ZN(n13658) );
NAND4_X2 U10413 ( .A1(n13660), .A2(n13183), .A3(n13659), .A4(n13658), .ZN(n3876) );
NAND2_X2 U10414 ( .A1(N865), .A2(n13180), .ZN(n13663) );
NAND2_X2 U10415 ( .A1(n13219), .A2(n14431), .ZN(n13662) );
NAND4_X2 U10416 ( .A1(n13663), .A2(n13183), .A3(n13662), .A4(n13661), .ZN(n4003) );
NAND2_X2 U10417 ( .A1(N897), .A2(n13167), .ZN(n13666) );
NAND2_X2 U10418 ( .A1(next_C[11]), .A2(n13148), .ZN(n13665) );
NAND2_X2 U10419 ( .A1(n13173), .A2(n14431), .ZN(n13664) );
NAND4_X2 U10420 ( .A1(n13666), .A2(n13152), .A3(n13665), .A4(n13664), .ZN(n3939) );
NAND2_X2 U10421 ( .A1(N927), .A2(n13180), .ZN(n13669) );
NAND2_X2 U10422 ( .A1(n13218), .A2(SHA1_result[75]), .ZN(n13668) );
NAND2_X2 U10423 ( .A1(n13204), .A2(next_C[11]), .ZN(n13667) );
NAND4_X2 U10424 ( .A1(n13669), .A2(n13183), .A3(n13668), .A4(n13667), .ZN(n3909) );
NAND2_X2 U10425 ( .A1(n13204), .A2(SHA1_result[75]), .ZN(n13672) );
NAND2_X2 U10426 ( .A1(N959), .A2(n13210), .ZN(n13671) );
NAND2_X2 U10427 ( .A1(n13218), .A2(n14810), .ZN(n13670) );
NAND3_X2 U10428 ( .A1(n13672), .A2(n13671), .A3(n13670), .ZN(n3877) );
NAND2_X2 U10429 ( .A1(N864), .A2(n13210), .ZN(n13674) );
NAND2_X2 U10430 ( .A1(n13218), .A2(n14434), .ZN(n13673) );
NAND3_X2 U10431 ( .A1(n13675), .A2(n13674), .A3(n13673), .ZN(n4004) );
NAND2_X2 U10432 ( .A1(N896), .A2(n13167), .ZN(n13678) );
NAND2_X2 U10433 ( .A1(next_C[10]), .A2(n13224), .ZN(n13677) );
NAND2_X2 U10434 ( .A1(n13173), .A2(n14434), .ZN(n13676) );
NAND3_X2 U10435 ( .A1(n13678), .A2(n13677), .A3(n13676), .ZN(n3940) );
NAND2_X2 U10436 ( .A1(N926), .A2(n13180), .ZN(n13681) );
NAND2_X2 U10437 ( .A1(n13218), .A2(SHA1_result[74]), .ZN(n13680) );
NAND2_X2 U10438 ( .A1(n13204), .A2(next_C[10]), .ZN(n13679) );
NAND4_X2 U10439 ( .A1(n13681), .A2(n13183), .A3(n13680), .A4(n13679), .ZN(n3910) );
NAND2_X2 U10440 ( .A1(N958), .A2(n13180), .ZN(n13684) );
NAND2_X2 U10441 ( .A1(n13218), .A2(SHA1_result[42]), .ZN(n13683) );
NAND2_X2 U10442 ( .A1(n13205), .A2(SHA1_result[74]), .ZN(n13682) );
NAND4_X2 U10443 ( .A1(n13684), .A2(n13183), .A3(n13683), .A4(n13682), .ZN(n3878) );
NAND2_X2 U10444 ( .A1(next_A[11]), .A2(n13206), .ZN(n13687) );
NAND2_X2 U10445 ( .A1(N863), .A2(n13210), .ZN(n13686) );
NAND2_X2 U10446 ( .A1(n13218), .A2(n14437), .ZN(n13685) );
NAND3_X2 U10447 ( .A1(n13687), .A2(n13686), .A3(n13685), .ZN(n4005) );
NAND2_X2 U10448 ( .A1(N895), .A2(n13167), .ZN(n13690) );
NAND2_X2 U10449 ( .A1(next_C[9]), .A2(n13148), .ZN(n13689) );
NAND2_X2 U10450 ( .A1(n13173), .A2(n14437), .ZN(n13688) );
NAND4_X2 U10451 ( .A1(n13690), .A2(n13152), .A3(n13689), .A4(n13688), .ZN(n3941) );
NAND2_X2 U10452 ( .A1(n13205), .A2(next_C[9]), .ZN(n13693) );
NAND2_X2 U10453 ( .A1(N925), .A2(n13210), .ZN(n13692) );
NAND2_X2 U10454 ( .A1(n13218), .A2(SHA1_result[73]), .ZN(n13691) );
NAND3_X2 U10455 ( .A1(n13693), .A2(n13692), .A3(n13691), .ZN(n3911) );
NAND2_X2 U10456 ( .A1(n13205), .A2(SHA1_result[73]), .ZN(n13696) );
NAND2_X2 U10457 ( .A1(N957), .A2(n13210), .ZN(n13695) );
NAND2_X2 U10458 ( .A1(n13218), .A2(n14797), .ZN(n13694) );
NAND3_X2 U10459 ( .A1(n13696), .A2(n13695), .A3(n13694), .ZN(n3879) );
NAND2_X2 U10460 ( .A1(N862), .A2(n13210), .ZN(n13698) );
NAND2_X2 U10461 ( .A1(n13218), .A2(n14440), .ZN(n13697) );
NAND3_X2 U10462 ( .A1(n13699), .A2(n13698), .A3(n13697), .ZN(n4006) );
NAND2_X2 U10463 ( .A1(N894), .A2(n13168), .ZN(n13702) );
NAND2_X2 U10464 ( .A1(next_C[8]), .A2(n13224), .ZN(n13701) );
NAND2_X2 U10465 ( .A1(n13174), .A2(n14440), .ZN(n13700) );
NAND3_X2 U10466 ( .A1(n13702), .A2(n13701), .A3(n13700), .ZN(n3942) );
NAND2_X2 U10467 ( .A1(n13204), .A2(next_C[8]), .ZN(n13705) );
NAND2_X2 U10468 ( .A1(N924), .A2(n13210), .ZN(n13704) );
NAND2_X2 U10469 ( .A1(n13218), .A2(SHA1_result[72]), .ZN(n13703) );
NAND3_X2 U10470 ( .A1(n13705), .A2(n13704), .A3(n13703), .ZN(n3912) );
NAND2_X2 U10471 ( .A1(n13205), .A2(SHA1_result[72]), .ZN(n13708) );
NAND2_X2 U10472 ( .A1(N956), .A2(n13210), .ZN(n13707) );
NAND2_X2 U10473 ( .A1(n13218), .A2(SHA1_result[40]), .ZN(n13706) );
NAND3_X2 U10474 ( .A1(n13708), .A2(n13707), .A3(n13706), .ZN(n3880) );
NAND2_X2 U10475 ( .A1(N861), .A2(n13180), .ZN(n13711) );
NAND2_X2 U10476 ( .A1(n13217), .A2(n14443), .ZN(n13710) );
NAND4_X2 U10477 ( .A1(n13711), .A2(n13183), .A3(n13710), .A4(n13709), .ZN(n4007) );
NAND2_X2 U10478 ( .A1(N893), .A2(n13168), .ZN(n13714) );
NAND2_X2 U10479 ( .A1(next_C[7]), .A2(n13148), .ZN(n13713) );
NAND2_X2 U10480 ( .A1(n13174), .A2(n14443), .ZN(n13712) );
NAND4_X2 U10481 ( .A1(n13714), .A2(n13152), .A3(n13713), .A4(n13712), .ZN(n3943) );
NAND2_X2 U10482 ( .A1(N923), .A2(n13180), .ZN(n13717) );
NAND2_X2 U10483 ( .A1(n13217), .A2(SHA1_result[71]), .ZN(n13716) );
NAND2_X2 U10484 ( .A1(n13205), .A2(next_C[7]), .ZN(n13715) );
NAND4_X2 U10485 ( .A1(n13717), .A2(n13183), .A3(n13716), .A4(n13715), .ZN(n3913) );
NAND2_X2 U10486 ( .A1(n13205), .A2(SHA1_result[71]), .ZN(n13720) );
NAND2_X2 U10487 ( .A1(N955), .A2(n13210), .ZN(n13719) );
NAND2_X2 U10488 ( .A1(n13217), .A2(SHA1_result[39]), .ZN(n13718) );
NAND3_X2 U10489 ( .A1(n13720), .A2(n13719), .A3(n13718), .ZN(n3881) );
NAND2_X2 U10490 ( .A1(N860), .A2(n13180), .ZN(n13723) );
NAND2_X2 U10491 ( .A1(n13217), .A2(SHA1_result_136), .ZN(n13722) );
NAND2_X2 U10492 ( .A1(next_A[8]), .A2(n13206), .ZN(n13721) );
NAND4_X2 U10493 ( .A1(n13723), .A2(n13183), .A3(n13722), .A4(n13721), .ZN(n4008) );
NAND2_X2 U10494 ( .A1(N892), .A2(n13168), .ZN(n13726) );
NAND2_X2 U10495 ( .A1(next_C[6]), .A2(n13148), .ZN(n13725) );
NAND2_X2 U10496 ( .A1(n13174), .A2(SHA1_result_136), .ZN(n13724) );
NAND4_X2 U10497 ( .A1(n13726), .A2(n13152), .A3(n13725), .A4(n13724), .ZN(n3944) );
NAND2_X2 U10498 ( .A1(N922), .A2(n13181), .ZN(n13729) );
NAND2_X2 U10499 ( .A1(n13217), .A2(SHA1_result[70]), .ZN(n13728) );
NAND2_X2 U10500 ( .A1(n13203), .A2(next_C[6]), .ZN(n13727) );
NAND4_X2 U10501 ( .A1(n13729), .A2(n13183), .A3(n13728), .A4(n13727), .ZN(n3914) );
NAND2_X2 U10502 ( .A1(N954), .A2(n13181), .ZN(n13732) );
INV_X4 U10503 ( .A(n437), .ZN(n14778) );
NAND2_X2 U10504 ( .A1(n13217), .A2(n14778), .ZN(n13731) );
NAND2_X2 U10505 ( .A1(n13205), .A2(SHA1_result[70]), .ZN(n13730) );
NAND4_X2 U10506 ( .A1(n13732), .A2(n13183), .A3(n13731), .A4(n13730), .ZN(n3882) );
NAND2_X2 U10507 ( .A1(N859), .A2(n13210), .ZN(n13734) );
NAND2_X2 U10508 ( .A1(n13217), .A2(SHA1_result_135), .ZN(n13733) );
NAND3_X2 U10509 ( .A1(n13735), .A2(n13734), .A3(n13733), .ZN(n4009) );
NAND2_X2 U10510 ( .A1(N891), .A2(n13168), .ZN(n13738) );
NAND2_X2 U10511 ( .A1(next_C[5]), .A2(n13148), .ZN(n13737) );
NAND2_X2 U10512 ( .A1(n13174), .A2(SHA1_result_135), .ZN(n13736) );
NAND4_X2 U10513 ( .A1(n13738), .A2(n13152), .A3(n13737), .A4(n13736), .ZN(n3945) );
NAND2_X2 U10514 ( .A1(N921), .A2(n13181), .ZN(n13741) );
NAND2_X2 U10515 ( .A1(n13217), .A2(SHA1_result[69]), .ZN(n13740) );
NAND2_X2 U10516 ( .A1(n13204), .A2(next_C[5]), .ZN(n13739) );
NAND4_X2 U10517 ( .A1(n13741), .A2(n13183), .A3(n13740), .A4(n13739), .ZN(n3915) );
NAND2_X2 U10518 ( .A1(N953), .A2(n13181), .ZN(n13744) );
INV_X4 U10519 ( .A(n438), .ZN(n14770) );
NAND2_X2 U10520 ( .A1(n13217), .A2(n14770), .ZN(n13743) );
NAND2_X2 U10521 ( .A1(n13205), .A2(SHA1_result[69]), .ZN(n13742) );
NAND4_X2 U10522 ( .A1(n13744), .A2(n13185), .A3(n13743), .A4(n13742), .ZN(n3883) );
NAND2_X2 U10523 ( .A1(next_A[6]), .A2(n13206), .ZN(n13747) );
NAND2_X2 U10524 ( .A1(N858), .A2(n13209), .ZN(n13746) );
NAND2_X2 U10525 ( .A1(n13217), .A2(SHA1_result_134), .ZN(n13745) );
NAND3_X2 U10526 ( .A1(n13747), .A2(n13746), .A3(n13745), .ZN(n4010) );
NAND2_X2 U10527 ( .A1(N890), .A2(n13168), .ZN(n13750) );
NAND2_X2 U10528 ( .A1(next_C[4]), .A2(n13224), .ZN(n13749) );
NAND2_X2 U10529 ( .A1(n13174), .A2(SHA1_result_134), .ZN(n13748) );
NAND3_X2 U10530 ( .A1(n13750), .A2(n13749), .A3(n13748), .ZN(n3946) );
NAND2_X2 U10531 ( .A1(N920), .A2(n13181), .ZN(n13753) );
NAND2_X2 U10532 ( .A1(n13217), .A2(SHA1_result[68]), .ZN(n13752) );
NAND2_X2 U10533 ( .A1(n13204), .A2(next_C[4]), .ZN(n13751) );
NAND4_X2 U10534 ( .A1(n13753), .A2(n13185), .A3(n13752), .A4(n13751), .ZN(n3916) );
NAND2_X2 U10535 ( .A1(N952), .A2(n13181), .ZN(n13756) );
NAND2_X2 U10536 ( .A1(n13216), .A2(SHA1_result[36]), .ZN(n13755) );
NAND2_X2 U10537 ( .A1(n13204), .A2(SHA1_result[68]), .ZN(n13754) );
NAND4_X2 U10538 ( .A1(n13756), .A2(n13185), .A3(n13755), .A4(n13754), .ZN(n3884) );
NAND2_X2 U10539 ( .A1(next_A[5]), .A2(n13206), .ZN(n13759) );
NAND2_X2 U10540 ( .A1(N857), .A2(n13209), .ZN(n13758) );
NAND2_X2 U10541 ( .A1(n13216), .A2(SHA1_result_133), .ZN(n13757) );
NAND3_X2 U10542 ( .A1(n13759), .A2(n13758), .A3(n13757), .ZN(n4011) );
NAND2_X2 U10543 ( .A1(N889), .A2(n13168), .ZN(n13762) );
NAND2_X2 U10544 ( .A1(n13174), .A2(SHA1_result_133), .ZN(n13760) );
NAND3_X2 U10545 ( .A1(n13762), .A2(n13761), .A3(n13760), .ZN(n3947) );
NAND2_X2 U10546 ( .A1(N919), .A2(n13181), .ZN(n13765) );
NAND2_X2 U10547 ( .A1(n13216), .A2(SHA1_result[67]), .ZN(n13764) );
NAND4_X2 U10548 ( .A1(n13765), .A2(n14601), .A3(n13764), .A4(n13763), .ZN(n3917) );
NAND2_X2 U10549 ( .A1(n13203), .A2(SHA1_result[67]), .ZN(n13768) );
NAND2_X2 U10550 ( .A1(N951), .A2(n13209), .ZN(n13767) );
NAND2_X2 U10551 ( .A1(n13216), .A2(SHA1_result[35]), .ZN(n13766) );
NAND3_X2 U10552 ( .A1(n13768), .A2(n13767), .A3(n13766), .ZN(n3885) );
NAND2_X2 U10553 ( .A1(next_A[4]), .A2(n13206), .ZN(n13771) );
NAND2_X2 U10554 ( .A1(N856), .A2(n13209), .ZN(n13770) );
NAND2_X2 U10555 ( .A1(n13216), .A2(SHA1_result_132), .ZN(n13769) );
NAND3_X2 U10556 ( .A1(n13771), .A2(n13770), .A3(n13769), .ZN(n4012) );
NAND2_X2 U10557 ( .A1(N888), .A2(n13168), .ZN(n13774) );
NAND2_X2 U10558 ( .A1(next_C[2]), .A2(n13224), .ZN(n13773) );
NAND2_X2 U10559 ( .A1(n13174), .A2(SHA1_result_132), .ZN(n13772) );
NAND3_X2 U10560 ( .A1(n13774), .A2(n13773), .A3(n13772), .ZN(n3948) );
NAND2_X2 U10561 ( .A1(N918), .A2(n13181), .ZN(n13777) );
NAND2_X2 U10562 ( .A1(n13216), .A2(SHA1_result[66]), .ZN(n13776) );
NAND2_X2 U10563 ( .A1(n13203), .A2(next_C[2]), .ZN(n13775) );
NAND4_X2 U10564 ( .A1(n13777), .A2(n14601), .A3(n13776), .A4(n13775), .ZN(n3918) );
NAND2_X2 U10565 ( .A1(N950), .A2(n13181), .ZN(n13780) );
NAND2_X2 U10566 ( .A1(n13216), .A2(SHA1_result[34]), .ZN(n13779) );
NAND2_X2 U10567 ( .A1(n13202), .A2(SHA1_result[66]), .ZN(n13778) );
NAND4_X2 U10568 ( .A1(n13780), .A2(n13185), .A3(n13779), .A4(n13778), .ZN(n3886) );
NAND2_X2 U10569 ( .A1(next_A[3]), .A2(n13205), .ZN(n13783) );
NAND2_X2 U10570 ( .A1(N855), .A2(n13209), .ZN(n13782) );
NAND2_X2 U10571 ( .A1(n13216), .A2(SHA1_result_131), .ZN(n13781) );
NAND3_X2 U10572 ( .A1(n13783), .A2(n13782), .A3(n13781), .ZN(n4013) );
NAND2_X2 U10573 ( .A1(N887), .A2(n13168), .ZN(n13786) );
NAND2_X2 U10574 ( .A1(next_C[1]), .A2(n13148), .ZN(n13785) );
NAND2_X2 U10575 ( .A1(n13174), .A2(SHA1_result_131), .ZN(n13784) );
NAND4_X2 U10576 ( .A1(n13786), .A2(n13152), .A3(n13785), .A4(n13784), .ZN(n3949) );
NAND2_X2 U10577 ( .A1(N917), .A2(n13181), .ZN(n13789) );
NAND2_X2 U10578 ( .A1(n13216), .A2(SHA1_result[65]), .ZN(n13788) );
NAND2_X2 U10579 ( .A1(n13202), .A2(next_C[1]), .ZN(n13787) );
NAND4_X2 U10580 ( .A1(n13789), .A2(n14601), .A3(n13788), .A4(n13787), .ZN(n3919) );
NAND2_X2 U10581 ( .A1(N949), .A2(n13181), .ZN(n13792) );
NAND2_X2 U10582 ( .A1(n13216), .A2(n14742), .ZN(n13791) );
NAND2_X2 U10583 ( .A1(n13202), .A2(SHA1_result[65]), .ZN(n13790) );
NAND4_X2 U10584 ( .A1(n13792), .A2(n13185), .A3(n13791), .A4(n13790), .ZN(n3887) );
NAND2_X2 U10585 ( .A1(next_A[2]), .A2(n13206), .ZN(n13795) );
NAND2_X2 U10586 ( .A1(N854), .A2(n13209), .ZN(n13794) );
NAND2_X2 U10587 ( .A1(n13216), .A2(SHA1_result_130), .ZN(n13793) );
NAND3_X2 U10588 ( .A1(n13795), .A2(n13794), .A3(n13793), .ZN(n4014) );
NAND2_X2 U10589 ( .A1(N886), .A2(n13168), .ZN(n13798) );
NAND2_X2 U10590 ( .A1(next_C[0]), .A2(n13224), .ZN(n13797) );
NAND2_X2 U10591 ( .A1(n13174), .A2(SHA1_result_130), .ZN(n13796) );
NAND3_X2 U10592 ( .A1(n13798), .A2(n13797), .A3(n13796), .ZN(n3950) );
NAND2_X2 U10593 ( .A1(n13201), .A2(next_C[0]), .ZN(n13801) );
NAND2_X2 U10594 ( .A1(N916), .A2(n13209), .ZN(n13800) );
NAND2_X2 U10595 ( .A1(n13215), .A2(SHA1_result[64]), .ZN(n13799) );
NAND3_X2 U10596 ( .A1(n13801), .A2(n13800), .A3(n13799), .ZN(n3920) );
NAND2_X2 U10597 ( .A1(n13201), .A2(SHA1_result[64]), .ZN(n13804) );
NAND2_X2 U10598 ( .A1(N948), .A2(n13209), .ZN(n13803) );
NAND2_X2 U10599 ( .A1(n13215), .A2(SHA1_result[32]), .ZN(n13802) );
NAND3_X2 U10600 ( .A1(n13804), .A2(n13803), .A3(n13802), .ZN(n3888) );
NAND2_X2 U10601 ( .A1(H4[31]), .A2(n13329), .ZN(n13807) );
NAND2_X2 U10602 ( .A1(n13351), .A2(SHA1_result[31]), .ZN(n13806) );
NAND3_X2 U10603 ( .A1(n13807), .A2(n13186), .A3(n13806), .ZN(n3761) );
NAND2_X2 U10604 ( .A1(N1010), .A2(n13168), .ZN(n13810) );
NAND2_X2 U10605 ( .A1(n13148), .A2(SHA1_result[30]), .ZN(n13809) );
NAND2_X2 U10606 ( .A1(n13174), .A2(SHA1_result[62]), .ZN(n13808) );
NAND4_X2 U10607 ( .A1(n13810), .A2(n13152), .A3(n13809), .A4(n13808), .ZN(n3794) );
NAND2_X2 U10608 ( .A1(H4[30]), .A2(n13329), .ZN(n13812) );
NAND2_X2 U10609 ( .A1(n13351), .A2(SHA1_result[30]), .ZN(n13811) );
NAND3_X2 U10610 ( .A1(n13812), .A2(n13187), .A3(n13811), .ZN(n3762) );
NAND2_X2 U10611 ( .A1(N1009), .A2(n13168), .ZN(n13815) );
NAND2_X2 U10612 ( .A1(n13215), .A2(SHA1_result[29]), .ZN(n13814) );
NAND2_X2 U10613 ( .A1(n13174), .A2(SHA1_result[61]), .ZN(n13813) );
NAND3_X2 U10614 ( .A1(n13815), .A2(n13814), .A3(n13813), .ZN(n3795) );
NAND2_X2 U10615 ( .A1(n13193), .A2(SHA1_result[29]), .ZN(n13817) );
NAND2_X2 U10616 ( .A1(H4[29]), .A2(n13329), .ZN(n13816) );
NAND2_X2 U10617 ( .A1(n13817), .A2(n13816), .ZN(n3763) );
NAND2_X2 U10618 ( .A1(N1008), .A2(n13169), .ZN(n13820) );
NAND2_X2 U10619 ( .A1(n13215), .A2(SHA1_result[28]), .ZN(n13819) );
NAND2_X2 U10620 ( .A1(n13175), .A2(SHA1_result[60]), .ZN(n13818) );
NAND3_X2 U10621 ( .A1(n13820), .A2(n13819), .A3(n13818), .ZN(n3796) );
NAND2_X2 U10622 ( .A1(n13193), .A2(SHA1_result[28]), .ZN(n13822) );
NAND2_X2 U10623 ( .A1(H4[28]), .A2(n13329), .ZN(n13821) );
NAND2_X2 U10624 ( .A1(n13822), .A2(n13821), .ZN(n3764) );
NAND2_X2 U10625 ( .A1(N1007), .A2(n13169), .ZN(n13825) );
NAND2_X2 U10626 ( .A1(n13215), .A2(SHA1_result[27]), .ZN(n13824) );
NAND2_X2 U10627 ( .A1(n13175), .A2(SHA1_result[59]), .ZN(n13823) );
NAND3_X2 U10628 ( .A1(n13825), .A2(n13824), .A3(n13823), .ZN(n3797) );
NAND2_X2 U10629 ( .A1(n13193), .A2(SHA1_result[27]), .ZN(n13827) );
NAND2_X2 U10630 ( .A1(H4[27]), .A2(n13329), .ZN(n13826) );
NAND2_X2 U10631 ( .A1(n13827), .A2(n13826), .ZN(n3765) );
NAND2_X2 U10632 ( .A1(N1006), .A2(n13169), .ZN(n13830) );
NAND2_X2 U10633 ( .A1(n13215), .A2(SHA1_result[26]), .ZN(n13829) );
NAND2_X2 U10634 ( .A1(n13175), .A2(SHA1_result[58]), .ZN(n13828) );
NAND3_X2 U10635 ( .A1(n13830), .A2(n13829), .A3(n13828), .ZN(n3798) );
NAND2_X2 U10636 ( .A1(n13193), .A2(SHA1_result[26]), .ZN(n13832) );
NAND2_X2 U10637 ( .A1(H4[26]), .A2(n13329), .ZN(n13831) );
NAND2_X2 U10638 ( .A1(n13832), .A2(n13831), .ZN(n3766) );
NAND2_X2 U10639 ( .A1(N1005), .A2(n13169), .ZN(n13835) );
NAND2_X2 U10640 ( .A1(n13148), .A2(SHA1_result[25]), .ZN(n13834) );
NAND2_X2 U10641 ( .A1(n13175), .A2(SHA1_result[57]), .ZN(n13833) );
NAND4_X2 U10642 ( .A1(n13835), .A2(n13152), .A3(n13834), .A4(n13833), .ZN(n3799) );
NAND2_X2 U10643 ( .A1(H4[25]), .A2(n13329), .ZN(n13837) );
NAND2_X2 U10644 ( .A1(n13351), .A2(SHA1_result[25]), .ZN(n13836) );
NAND3_X2 U10645 ( .A1(n13837), .A2(n13186), .A3(n13836), .ZN(n3767) );
NAND2_X2 U10646 ( .A1(N1004), .A2(n13169), .ZN(n13840) );
NAND2_X2 U10647 ( .A1(n13148), .A2(SHA1_result[24]), .ZN(n13839) );
NAND2_X2 U10648 ( .A1(n13175), .A2(SHA1_result[56]), .ZN(n13838) );
NAND4_X2 U10649 ( .A1(n13840), .A2(n13152), .A3(n13839), .A4(n13838), .ZN(n3800) );
NAND2_X2 U10650 ( .A1(H4[24]), .A2(n13329), .ZN(n13842) );
NAND2_X2 U10651 ( .A1(n13351), .A2(SHA1_result[24]), .ZN(n13841) );
NAND3_X2 U10652 ( .A1(n13842), .A2(n13192), .A3(n13841), .ZN(n3768) );
NAND2_X2 U10653 ( .A1(N1003), .A2(n13169), .ZN(n13845) );
NAND2_X2 U10654 ( .A1(n13148), .A2(SHA1_result[23]), .ZN(n13844) );
NAND2_X2 U10655 ( .A1(n13175), .A2(SHA1_result[55]), .ZN(n13843) );
NAND4_X2 U10656 ( .A1(n13845), .A2(n13152), .A3(n13844), .A4(n13843), .ZN(n3801) );
NAND2_X2 U10657 ( .A1(H4[23]), .A2(n13329), .ZN(n13847) );
NAND2_X2 U10658 ( .A1(n13351), .A2(SHA1_result[23]), .ZN(n13846) );
NAND3_X2 U10659 ( .A1(n13847), .A2(n13192), .A3(n13846), .ZN(n3769) );
NAND2_X2 U10660 ( .A1(N1002), .A2(n13169), .ZN(n13850) );
NAND2_X2 U10661 ( .A1(n13148), .A2(SHA1_result[22]), .ZN(n13849) );
NAND2_X2 U10662 ( .A1(n13175), .A2(n14681), .ZN(n13848) );
NAND4_X2 U10663 ( .A1(n13850), .A2(n13152), .A3(n13849), .A4(n13848), .ZN(n3802) );
NAND2_X2 U10664 ( .A1(H4[22]), .A2(n13329), .ZN(n13852) );
NAND2_X2 U10665 ( .A1(n13350), .A2(SHA1_result[22]), .ZN(n13851) );
NAND3_X2 U10666 ( .A1(n13852), .A2(n13192), .A3(n13851), .ZN(n3770) );
NAND2_X2 U10667 ( .A1(N1001), .A2(n13169), .ZN(n13855) );
NAND2_X2 U10668 ( .A1(n13215), .A2(SHA1_result[21]), .ZN(n13854) );
NAND2_X2 U10669 ( .A1(n13175), .A2(n14682), .ZN(n13853) );
NAND3_X2 U10670 ( .A1(n13855), .A2(n13854), .A3(n13853), .ZN(n3803) );
NAND2_X2 U10671 ( .A1(n13193), .A2(SHA1_result[21]), .ZN(n13857) );
NAND2_X2 U10672 ( .A1(H4[21]), .A2(n13328), .ZN(n13856) );
NAND2_X2 U10673 ( .A1(n13857), .A2(n13856), .ZN(n3771) );
NAND2_X2 U10674 ( .A1(N1000), .A2(n13169), .ZN(n13860) );
NAND2_X2 U10675 ( .A1(n13150), .A2(SHA1_result[20]), .ZN(n13859) );
NAND2_X2 U10676 ( .A1(n13175), .A2(n14868), .ZN(n13858) );
NAND4_X2 U10677 ( .A1(n13860), .A2(n13151), .A3(n13859), .A4(n13858), .ZN(n3804) );
NAND2_X2 U10678 ( .A1(H4[20]), .A2(n13328), .ZN(n13862) );
NAND2_X2 U10679 ( .A1(n13345), .A2(SHA1_result[20]), .ZN(n13861) );
NAND3_X2 U10680 ( .A1(n13862), .A2(n13192), .A3(n13861), .ZN(n3772) );
NAND2_X2 U10681 ( .A1(N999), .A2(n13169), .ZN(n13865) );
NAND2_X2 U10682 ( .A1(n13219), .A2(SHA1_result[19]), .ZN(n13864) );
NAND2_X2 U10683 ( .A1(n13175), .A2(SHA1_result[51]), .ZN(n13863) );
NAND3_X2 U10684 ( .A1(n13865), .A2(n13864), .A3(n13863), .ZN(n3805) );
NAND2_X2 U10685 ( .A1(n13193), .A2(SHA1_result[19]), .ZN(n13867) );
NAND2_X2 U10686 ( .A1(H4[19]), .A2(n13328), .ZN(n13866) );
NAND2_X2 U10687 ( .A1(n13867), .A2(n13866), .ZN(n3773) );
NAND2_X2 U10688 ( .A1(N998), .A2(n13169), .ZN(n13870) );
NAND2_X2 U10689 ( .A1(n13215), .A2(SHA1_result[18]), .ZN(n13869) );
NAND2_X2 U10690 ( .A1(n13175), .A2(SHA1_result[50]), .ZN(n13868) );
NAND3_X2 U10691 ( .A1(n13870), .A2(n13869), .A3(n13868), .ZN(n3806) );
NAND2_X2 U10692 ( .A1(n13193), .A2(SHA1_result[18]), .ZN(n13872) );
NAND2_X2 U10693 ( .A1(H4[18]), .A2(n13328), .ZN(n13871) );
NAND2_X2 U10694 ( .A1(n13872), .A2(n13871), .ZN(n3774) );
NAND2_X2 U10695 ( .A1(N997), .A2(n13170), .ZN(n13875) );
NAND2_X2 U10696 ( .A1(n13150), .A2(SHA1_result[17]), .ZN(n13874) );
NAND2_X2 U10697 ( .A1(n13176), .A2(SHA1_result[49]), .ZN(n13873) );
NAND4_X2 U10698 ( .A1(n13875), .A2(n13151), .A3(n13874), .A4(n13873), .ZN(n3807) );
NAND2_X2 U10699 ( .A1(H4[17]), .A2(n13328), .ZN(n13877) );
NAND2_X2 U10700 ( .A1(n13351), .A2(SHA1_result[17]), .ZN(n13876) );
NAND3_X2 U10701 ( .A1(n13877), .A2(n13192), .A3(n13876), .ZN(n3775) );
NAND2_X2 U10702 ( .A1(N996), .A2(n13170), .ZN(n13880) );
NAND2_X2 U10703 ( .A1(n13215), .A2(SHA1_result[16]), .ZN(n13879) );
NAND2_X2 U10704 ( .A1(n13176), .A2(SHA1_result[48]), .ZN(n13878) );
NAND3_X2 U10705 ( .A1(n13880), .A2(n13879), .A3(n13878), .ZN(n3808) );
NAND2_X2 U10706 ( .A1(n13193), .A2(SHA1_result[16]), .ZN(n13882) );
NAND2_X2 U10707 ( .A1(H4[16]), .A2(n13328), .ZN(n13881) );
NAND2_X2 U10708 ( .A1(n13882), .A2(n13881), .ZN(n3776) );
NAND2_X2 U10709 ( .A1(N995), .A2(n13170), .ZN(n13885) );
NAND2_X2 U10710 ( .A1(n13150), .A2(SHA1_result[15]), .ZN(n13884) );
NAND2_X2 U10711 ( .A1(n13176), .A2(SHA1_result[47]), .ZN(n13883) );
NAND4_X2 U10712 ( .A1(n13885), .A2(n13151), .A3(n13884), .A4(n13883), .ZN(n3809) );
NAND2_X2 U10713 ( .A1(H4[15]), .A2(n13328), .ZN(n13887) );
NAND2_X2 U10714 ( .A1(n13351), .A2(SHA1_result[15]), .ZN(n13886) );
NAND3_X2 U10715 ( .A1(n13887), .A2(n13192), .A3(n13886), .ZN(n3777) );
NAND2_X2 U10716 ( .A1(N994), .A2(n13170), .ZN(n13890) );
NAND2_X2 U10717 ( .A1(n13150), .A2(SHA1_result[14]), .ZN(n13889) );
NAND2_X2 U10718 ( .A1(n13176), .A2(n14830), .ZN(n13888) );
NAND4_X2 U10719 ( .A1(n13890), .A2(n13151), .A3(n13889), .A4(n13888), .ZN(n3810) );
NAND2_X2 U10720 ( .A1(H4[14]), .A2(n13328), .ZN(n13892) );
NAND2_X2 U10721 ( .A1(n13345), .A2(SHA1_result[14]), .ZN(n13891) );
NAND3_X2 U10722 ( .A1(n13892), .A2(n13192), .A3(n13891), .ZN(n3778) );
NAND2_X2 U10723 ( .A1(N993), .A2(n13170), .ZN(n13895) );
NAND2_X2 U10724 ( .A1(n13150), .A2(SHA1_result[13]), .ZN(n13894) );
NAND2_X2 U10725 ( .A1(n13176), .A2(SHA1_result[45]), .ZN(n13893) );
NAND4_X2 U10726 ( .A1(n13895), .A2(n13151), .A3(n13894), .A4(n13893), .ZN(n3811) );
NAND2_X2 U10727 ( .A1(H4[13]), .A2(n13328), .ZN(n13897) );
NAND2_X2 U10728 ( .A1(n13345), .A2(SHA1_result[13]), .ZN(n13896) );
NAND3_X2 U10729 ( .A1(n13897), .A2(n13192), .A3(n13896), .ZN(n3779) );
NAND2_X2 U10730 ( .A1(N992), .A2(n13170), .ZN(n13900) );
NAND2_X2 U10731 ( .A1(n13215), .A2(SHA1_result[12]), .ZN(n13899) );
NAND2_X2 U10732 ( .A1(n13176), .A2(n14817), .ZN(n13898) );
NAND3_X2 U10733 ( .A1(n13900), .A2(n13899), .A3(n13898), .ZN(n3812) );
NAND2_X2 U10734 ( .A1(n13193), .A2(SHA1_result[12]), .ZN(n13902) );
NAND2_X2 U10735 ( .A1(H4[12]), .A2(n13328), .ZN(n13901) );
NAND2_X2 U10736 ( .A1(n13902), .A2(n13901), .ZN(n3780) );
NAND2_X2 U10737 ( .A1(N991), .A2(n13170), .ZN(n13905) );
NAND2_X2 U10738 ( .A1(n13214), .A2(SHA1_result[11]), .ZN(n13904) );
NAND2_X2 U10739 ( .A1(n13176), .A2(n14810), .ZN(n13903) );
NAND3_X2 U10740 ( .A1(n13905), .A2(n13904), .A3(n13903), .ZN(n3813) );
NAND2_X2 U10741 ( .A1(n13193), .A2(SHA1_result[11]), .ZN(n13907) );
NAND2_X2 U10742 ( .A1(H4[11]), .A2(n13328), .ZN(n13906) );
NAND2_X2 U10743 ( .A1(n13907), .A2(n13906), .ZN(n3781) );
NAND2_X2 U10744 ( .A1(N990), .A2(n13170), .ZN(n13910) );
NAND2_X2 U10745 ( .A1(n13214), .A2(SHA1_result[10]), .ZN(n13909) );
NAND2_X2 U10746 ( .A1(n13176), .A2(SHA1_result[42]), .ZN(n13908) );
NAND3_X2 U10747 ( .A1(n13910), .A2(n13909), .A3(n13908), .ZN(n3814) );
NAND2_X2 U10748 ( .A1(n13193), .A2(SHA1_result[10]), .ZN(n13912) );
NAND2_X2 U10749 ( .A1(H4[10]), .A2(n13328), .ZN(n13911) );
NAND2_X2 U10750 ( .A1(n13912), .A2(n13911), .ZN(n3782) );
NAND2_X2 U10751 ( .A1(N989), .A2(n13170), .ZN(n13915) );
NAND2_X2 U10752 ( .A1(n13214), .A2(SHA1_result[9]), .ZN(n13914) );
NAND2_X2 U10753 ( .A1(n13176), .A2(n14797), .ZN(n13913) );
NAND3_X2 U10754 ( .A1(n13915), .A2(n13914), .A3(n13913), .ZN(n3815) );
NAND2_X2 U10755 ( .A1(n13194), .A2(SHA1_result[9]), .ZN(n13917) );
NAND2_X2 U10756 ( .A1(H4[9]), .A2(n13328), .ZN(n13916) );
NAND2_X2 U10757 ( .A1(n13917), .A2(n13916), .ZN(n3783) );
NAND2_X2 U10758 ( .A1(N988), .A2(n13170), .ZN(n13920) );
NAND2_X2 U10759 ( .A1(n13150), .A2(SHA1_result[8]), .ZN(n13919) );
NAND2_X2 U10760 ( .A1(n13176), .A2(SHA1_result[40]), .ZN(n13918) );
NAND4_X2 U10761 ( .A1(n13920), .A2(n13151), .A3(n13919), .A4(n13918), .ZN(n3816) );
NAND2_X2 U10762 ( .A1(H4[8]), .A2(n13328), .ZN(n13922) );
NAND2_X2 U10763 ( .A1(n13345), .A2(SHA1_result[8]), .ZN(n13921) );
NAND3_X2 U10764 ( .A1(n13922), .A2(n13192), .A3(n13921), .ZN(n3784) );
NAND2_X2 U10765 ( .A1(N987), .A2(n13170), .ZN(n13925) );
NAND2_X2 U10766 ( .A1(n13150), .A2(SHA1_result[7]), .ZN(n13924) );
NAND2_X2 U10767 ( .A1(n13176), .A2(SHA1_result[39]), .ZN(n13923) );
NAND4_X2 U10768 ( .A1(n13925), .A2(n13151), .A3(n13924), .A4(n13923), .ZN(n3817) );
NAND2_X2 U10769 ( .A1(H4[7]), .A2(n13328), .ZN(n13927) );
NAND2_X2 U10770 ( .A1(n13345), .A2(SHA1_result[7]), .ZN(n13926) );
NAND3_X2 U10771 ( .A1(n13927), .A2(n13192), .A3(n13926), .ZN(n3785) );
NAND2_X2 U10772 ( .A1(N986), .A2(n13171), .ZN(n13930) );
NAND2_X2 U10773 ( .A1(n13150), .A2(SHA1_result[6]), .ZN(n13929) );
NAND2_X2 U10774 ( .A1(n13177), .A2(n14778), .ZN(n13928) );
NAND4_X2 U10775 ( .A1(n13930), .A2(n13151), .A3(n13929), .A4(n13928), .ZN(n3818) );
NAND2_X2 U10776 ( .A1(H4[6]), .A2(n13328), .ZN(n13932) );
NAND2_X2 U10777 ( .A1(n13345), .A2(SHA1_result[6]), .ZN(n13931) );
NAND3_X2 U10778 ( .A1(n13932), .A2(n13192), .A3(n13931), .ZN(n3786) );
NAND2_X2 U10779 ( .A1(N985), .A2(n13171), .ZN(n13935) );
NAND2_X2 U10780 ( .A1(n13150), .A2(SHA1_result[5]), .ZN(n13934) );
NAND2_X2 U10781 ( .A1(n13177), .A2(n14770), .ZN(n13933) );
NAND4_X2 U10782 ( .A1(n13935), .A2(n13151), .A3(n13934), .A4(n13933), .ZN(n3819) );
NAND2_X2 U10783 ( .A1(H4[5]), .A2(n13328), .ZN(n13937) );
NAND2_X2 U10784 ( .A1(n13345), .A2(SHA1_result[5]), .ZN(n13936) );
NAND3_X2 U10785 ( .A1(n13937), .A2(n13192), .A3(n13936), .ZN(n3787) );
NAND2_X2 U10786 ( .A1(N984), .A2(n13171), .ZN(n13940) );
NAND2_X2 U10787 ( .A1(n13150), .A2(SHA1_result[4]), .ZN(n13939) );
NAND2_X2 U10788 ( .A1(n13177), .A2(SHA1_result[36]), .ZN(n13938) );
NAND4_X2 U10789 ( .A1(n13940), .A2(n13151), .A3(n13939), .A4(n13938), .ZN(n3820) );
NAND2_X2 U10790 ( .A1(H4[4]), .A2(n13328), .ZN(n13942) );
NAND2_X2 U10791 ( .A1(n13345), .A2(SHA1_result[4]), .ZN(n13941) );
NAND3_X2 U10792 ( .A1(n13942), .A2(n13191), .A3(n13941), .ZN(n3788) );
NAND2_X2 U10793 ( .A1(N983), .A2(n13171), .ZN(n13945) );
NAND2_X2 U10794 ( .A1(n13214), .A2(SHA1_result[3]), .ZN(n13944) );
NAND2_X2 U10795 ( .A1(n13177), .A2(SHA1_result[35]), .ZN(n13943) );
NAND3_X2 U10796 ( .A1(n13945), .A2(n13944), .A3(n13943), .ZN(n3821) );
NAND2_X2 U10797 ( .A1(n13194), .A2(SHA1_result[3]), .ZN(n13947) );
NAND2_X2 U10798 ( .A1(H4[3]), .A2(n13328), .ZN(n13946) );
NAND2_X2 U10799 ( .A1(n13947), .A2(n13946), .ZN(n3789) );
NAND2_X2 U10800 ( .A1(N982), .A2(n13171), .ZN(n13950) );
NAND2_X2 U10801 ( .A1(n13214), .A2(SHA1_result[2]), .ZN(n13949) );
NAND2_X2 U10802 ( .A1(n13177), .A2(SHA1_result[34]), .ZN(n13948) );
NAND3_X2 U10803 ( .A1(n13950), .A2(n13949), .A3(n13948), .ZN(n3822) );
NAND2_X2 U10804 ( .A1(n13194), .A2(SHA1_result[2]), .ZN(n13952) );
NAND2_X2 U10805 ( .A1(H4[2]), .A2(n13327), .ZN(n13951) );
NAND2_X2 U10806 ( .A1(n13952), .A2(n13951), .ZN(n3790) );
NAND2_X2 U10807 ( .A1(N981), .A2(n13171), .ZN(n13955) );
NAND2_X2 U10808 ( .A1(n13214), .A2(SHA1_result[1]), .ZN(n13954) );
NAND2_X2 U10809 ( .A1(n13177), .A2(n14742), .ZN(n13953) );
NAND3_X2 U10810 ( .A1(n13955), .A2(n13954), .A3(n13953), .ZN(n3823) );
NAND2_X2 U10811 ( .A1(n13194), .A2(SHA1_result[1]), .ZN(n13957) );
NAND2_X2 U10812 ( .A1(H4[1]), .A2(n13327), .ZN(n13956) );
NAND2_X2 U10813 ( .A1(n13957), .A2(n13956), .ZN(n3791) );
NAND2_X2 U10814 ( .A1(N980), .A2(n13171), .ZN(n13960) );
NAND2_X2 U10815 ( .A1(n13214), .A2(SHA1_result[0]), .ZN(n13959) );
NAND2_X2 U10816 ( .A1(n13177), .A2(SHA1_result[32]), .ZN(n13958) );
NAND3_X2 U10817 ( .A1(n13960), .A2(n13959), .A3(n13958), .ZN(n3824) );
NAND2_X2 U10818 ( .A1(n13194), .A2(SHA1_result[0]), .ZN(n13962) );
NAND2_X2 U10819 ( .A1(H4[0]), .A2(n13327), .ZN(n13961) );
NAND2_X2 U10820 ( .A1(n13962), .A2(n13961), .ZN(n3792) );
NAND2_X2 U10821 ( .A1(N1011), .A2(n13171), .ZN(n13965) );
NAND2_X2 U10822 ( .A1(n13150), .A2(SHA1_result[31]), .ZN(n13964) );
NAND2_X2 U10823 ( .A1(n13177), .A2(SHA1_result[63]), .ZN(n13963) );
NAND4_X2 U10824 ( .A1(n13965), .A2(n13152), .A3(n13964), .A4(n13963), .ZN(n3793) );
NAND3_X2 U10825 ( .A1(n13966), .A2(n13967), .A3(n14688), .ZN(n14273) );
INV_X4 U10826 ( .A(n13970), .ZN(n13969) );
NAND2_X2 U10827 ( .A1(n13970), .A2(n14953), .ZN(n13978) );
NAND2_X2 U10828 ( .A1(n13983), .A2(n13978), .ZN(N2585) );
NAND2_X2 U10829 ( .A1(n13116), .A2(n14061), .ZN(n13971) );
NAND2_X2 U10830 ( .A1(n14688), .A2(n13076), .ZN(n13972) );
INV_X4 U10831 ( .A(n13972), .ZN(n14266) );
NAND3_X2 U10832 ( .A1(n13975), .A2(n14953), .A3(n13974), .ZN(n13980) );
NAND2_X2 U10833 ( .A1(n13982), .A2(n13980), .ZN(N2583) );
INV_X4 U10834 ( .A(N2583), .ZN(n13976) );
NAND2_X2 U10835 ( .A1(n13978), .A2(n13976), .ZN(N2590) );
INV_X4 U10836 ( .A(n13980), .ZN(n14962) );
INV_X4 U10837 ( .A(n13982), .ZN(n8328) );
INV_X4 U10838 ( .A(N2590), .ZN(n13977) );
NAND2_X2 U10839 ( .A1(n13983), .A2(n13977), .ZN(N2589) );
NAND2_X2 U10840 ( .A1(n13983), .A2(n13980), .ZN(n8330) );
INV_X4 U10841 ( .A(n13983), .ZN(n14931) );
NAND2_X2 U10842 ( .A1(n13978), .A2(n13980), .ZN(N2595) );
INV_X4 U10843 ( .A(n13978), .ZN(n14932) );
INV_X4 U10844 ( .A(N2585), .ZN(n13979) );
NAND2_X2 U10845 ( .A1(n13982), .A2(n13979), .ZN(N2587) );
NAND2_X2 U10846 ( .A1(n13980), .A2(n13979), .ZN(n14960) );
INV_X4 U10847 ( .A(n8330), .ZN(n13981) );
NAND2_X2 U10848 ( .A1(n13982), .A2(n13981), .ZN(N2592) );
NAND2_X2 U10849 ( .A1(n13983), .A2(n13982), .ZN(n14961) );
NAND2_X2 U10850 ( .A1(n13156), .A2(Wt[31]), .ZN(n13984) );
NAND3_X2 U10851 ( .A1(n9509), .A2(n9510), .A3(n13984), .ZN(n4496) );
NAND2_X2 U10852 ( .A1(n13156), .A2(Wt[30]), .ZN(n13985) );
NAND3_X2 U10853 ( .A1(n9503), .A2(n9504), .A3(n13985), .ZN(n4497) );
NAND2_X2 U10854 ( .A1(n13156), .A2(Wt[29]), .ZN(n13986) );
NAND3_X2 U10855 ( .A1(n9497), .A2(n9498), .A3(n13986), .ZN(n4498) );
NAND2_X2 U10856 ( .A1(n13156), .A2(Wt[28]), .ZN(n13987) );
NAND3_X2 U10857 ( .A1(n9491), .A2(n9492), .A3(n13987), .ZN(n4499) );
NAND2_X2 U10858 ( .A1(n13156), .A2(Wt[27]), .ZN(n13988) );
NAND3_X2 U10859 ( .A1(n9485), .A2(n9486), .A3(n13988), .ZN(n4500) );
NAND2_X2 U10860 ( .A1(n13156), .A2(Wt[26]), .ZN(n13989) );
NAND3_X2 U10861 ( .A1(n9479), .A2(n9480), .A3(n13989), .ZN(n4501) );
NAND2_X2 U10862 ( .A1(n13156), .A2(Wt[25]), .ZN(n13990) );
NAND3_X2 U10863 ( .A1(n9473), .A2(n9474), .A3(n13990), .ZN(n4502) );
NAND2_X2 U10864 ( .A1(n13156), .A2(Wt[24]), .ZN(n13991) );
NAND3_X2 U10865 ( .A1(n9467), .A2(n9468), .A3(n13991), .ZN(n4503) );
NAND2_X2 U10866 ( .A1(n13156), .A2(Wt[23]), .ZN(n13992) );
NAND3_X2 U10867 ( .A1(n9461), .A2(n9462), .A3(n13992), .ZN(n4504) );
NAND2_X2 U10868 ( .A1(n13156), .A2(Wt[22]), .ZN(n13993) );
NAND3_X2 U10869 ( .A1(n9455), .A2(n9456), .A3(n13993), .ZN(n4505) );
NAND2_X2 U10870 ( .A1(n13155), .A2(Wt[21]), .ZN(n13994) );
NAND3_X2 U10871 ( .A1(n9449), .A2(n9450), .A3(n13994), .ZN(n4506) );
NAND2_X2 U10872 ( .A1(n13155), .A2(Wt[20]), .ZN(n13995) );
NAND3_X2 U10873 ( .A1(n9443), .A2(n9444), .A3(n13995), .ZN(n4507) );
NAND2_X2 U10874 ( .A1(n13155), .A2(Wt[19]), .ZN(n13996) );
NAND3_X2 U10875 ( .A1(n9437), .A2(n9438), .A3(n13996), .ZN(n4508) );
NAND2_X2 U10876 ( .A1(n13155), .A2(Wt[18]), .ZN(n13997) );
NAND3_X2 U10877 ( .A1(n9431), .A2(n9432), .A3(n13997), .ZN(n4509) );
NAND2_X2 U10878 ( .A1(n13026), .A2(n13998), .ZN(n13999) );
NAND3_X2 U10879 ( .A1(n14000), .A2(n14953), .A3(n13999), .ZN(n14001) );
NAND2_X2 U10880 ( .A1(n13155), .A2(Wt[17]), .ZN(n14004) );
INV_X4 U10881 ( .A(n14687), .ZN(n14002) );
NAND2_X2 U10882 ( .A1(n9428), .A2(n13317), .ZN(n14003) );
NAND3_X2 U10883 ( .A1(n14005), .A2(n14004), .A3(n14003), .ZN(n4510) );
NAND2_X2 U10884 ( .A1(n13155), .A2(Wt[16]), .ZN(n14007) );
NAND2_X2 U10885 ( .A1(n9422), .A2(n13317), .ZN(n14006) );
NAND3_X2 U10886 ( .A1(n14008), .A2(n14007), .A3(n14006), .ZN(n4511) );
NAND2_X2 U10887 ( .A1(n13155), .A2(Wt[15]), .ZN(n14010) );
NAND2_X2 U10888 ( .A1(n9416), .A2(n13317), .ZN(n14009) );
NAND3_X2 U10889 ( .A1(n14011), .A2(n14010), .A3(n14009), .ZN(n4512) );
NAND2_X2 U10890 ( .A1(n13155), .A2(Wt[14]), .ZN(n14013) );
NAND2_X2 U10891 ( .A1(n9410), .A2(n13317), .ZN(n14012) );
NAND3_X2 U10892 ( .A1(n14014), .A2(n14013), .A3(n14012), .ZN(n4513) );
NAND2_X2 U10893 ( .A1(n13155), .A2(Wt[13]), .ZN(n14016) );
NAND2_X2 U10894 ( .A1(n9404), .A2(n13317), .ZN(n14015) );
NAND3_X2 U10895 ( .A1(n14017), .A2(n14016), .A3(n14015), .ZN(n4514) );
NAND2_X2 U10896 ( .A1(n13155), .A2(Wt[12]), .ZN(n14019) );
NAND2_X2 U10897 ( .A1(n9398), .A2(n13316), .ZN(n14018) );
NAND3_X2 U10898 ( .A1(n14020), .A2(n14019), .A3(n14018), .ZN(n4515) );
NAND2_X2 U10899 ( .A1(n13155), .A2(Wt[11]), .ZN(n14022) );
NAND2_X2 U10900 ( .A1(n9392), .A2(n13316), .ZN(n14021) );
NAND3_X2 U10901 ( .A1(n14023), .A2(n14022), .A3(n14021), .ZN(n4516) );
NAND2_X2 U10902 ( .A1(n13154), .A2(Wt[10]), .ZN(n14025) );
NAND2_X2 U10903 ( .A1(n9386), .A2(n13316), .ZN(n14024) );
NAND3_X2 U10904 ( .A1(n14026), .A2(n14025), .A3(n14024), .ZN(n4517) );
NAND2_X2 U10905 ( .A1(n13154), .A2(Wt[9]), .ZN(n14028) );
NAND2_X2 U10906 ( .A1(n9380), .A2(n13316), .ZN(n14027) );
NAND3_X2 U10907 ( .A1(n14029), .A2(n14028), .A3(n14027), .ZN(n4518) );
NAND2_X2 U10908 ( .A1(n13154), .A2(Wt[8]), .ZN(n14031) );
NAND2_X2 U10909 ( .A1(n9374), .A2(n13316), .ZN(n14030) );
NAND3_X2 U10910 ( .A1(n14032), .A2(n14031), .A3(n14030), .ZN(n4519) );
NAND2_X2 U10911 ( .A1(n13154), .A2(Wt[7]), .ZN(n14034) );
NAND2_X2 U10912 ( .A1(n9368), .A2(n13316), .ZN(n14033) );
NAND3_X2 U10913 ( .A1(n14035), .A2(n14034), .A3(n14033), .ZN(n4520) );
NAND2_X2 U10914 ( .A1(n13154), .A2(Wt[6]), .ZN(n14037) );
NAND2_X2 U10915 ( .A1(n9362), .A2(n13316), .ZN(n14036) );
NAND3_X2 U10916 ( .A1(n14038), .A2(n14037), .A3(n14036), .ZN(n4521) );
NAND2_X2 U10917 ( .A1(n13154), .A2(Wt[5]), .ZN(n14040) );
NAND2_X2 U10918 ( .A1(n9356), .A2(n13316), .ZN(n14039) );
NAND3_X2 U10919 ( .A1(n14041), .A2(n14040), .A3(n14039), .ZN(n4522) );
NAND2_X2 U10920 ( .A1(n13154), .A2(Wt[4]), .ZN(n14043) );
NAND2_X2 U10921 ( .A1(n9350), .A2(n13316), .ZN(n14042) );
NAND3_X2 U10922 ( .A1(n14044), .A2(n14043), .A3(n14042), .ZN(n4523) );
NAND2_X2 U10923 ( .A1(n13154), .A2(Wt[3]), .ZN(n14046) );
NAND2_X2 U10924 ( .A1(n9344), .A2(n13316), .ZN(n14045) );
NAND3_X2 U10925 ( .A1(n14047), .A2(n14046), .A3(n14045), .ZN(n4524) );
NAND2_X2 U10926 ( .A1(n13154), .A2(Wt[2]), .ZN(n14049) );
NAND2_X2 U10927 ( .A1(n9338), .A2(n13316), .ZN(n14048) );
NAND3_X2 U10928 ( .A1(n14050), .A2(n14049), .A3(n14048), .ZN(n4525) );
NAND2_X2 U10929 ( .A1(n13154), .A2(Wt[1]), .ZN(n14052) );
NAND2_X2 U10930 ( .A1(n9332), .A2(n13316), .ZN(n14051) );
NAND3_X2 U10931 ( .A1(n14053), .A2(n14052), .A3(n14051), .ZN(n4526) );
NAND2_X2 U10932 ( .A1(n13319), .A2(n13063), .ZN(n14056) );
NAND2_X2 U10933 ( .A1(n13154), .A2(Wt[0]), .ZN(n14055) );
NAND2_X2 U10934 ( .A1(n9325), .A2(n13317), .ZN(n14054) );
NAND3_X2 U10935 ( .A1(n14056), .A2(n14055), .A3(n14054), .ZN(n4527) );
NAND2_X2 U10936 ( .A1(next_A[1]), .A2(n13205), .ZN(n14059) );
NAND2_X2 U10937 ( .A1(N853), .A2(n13209), .ZN(n14058) );
NAND2_X2 U10938 ( .A1(n13214), .A2(SHA1_result_129), .ZN(n14057) );
NAND3_X2 U10939 ( .A1(n14059), .A2(n14058), .A3(n14057), .ZN(n4015) );
INV_X4 U10940 ( .A(n14063), .ZN(n14074) );
MUX2_X2 U10941 ( .A(n13158), .B(n13162), .S(next_C[29]), .Z(n14070) );
NAND2_X2 U10942 ( .A1(n14070), .A2(SHA1_result[63]), .ZN(n14081) );
XOR2_X2 U10943 ( .A(n13002), .B(n412), .Z(n14077) );
NOR2_X2 U10944 ( .A1(n14076), .A2(n14075), .ZN(n14079) );
NAND2_X2 U10945 ( .A1(n13096), .A2(n14077), .ZN(n14078) );
MUX2_X2 U10946 ( .A(n14079), .B(n14078), .S(n444), .Z(n14080) );
NAND2_X2 U10947 ( .A1(n14081), .A2(n14080), .ZN(SHA1_ft_BCD[31]) );
MUX2_X2 U10948 ( .A(n13158), .B(n13164), .S(next_C[28]), .Z(n14082) );
NAND2_X2 U10949 ( .A1(n14082), .A2(SHA1_result[62]), .ZN(n14089) );
XOR2_X2 U10950 ( .A(SHA1_result[62]), .B(next_C[28]), .Z(n14085) );
NOR2_X2 U10951 ( .A1(n14084), .A2(n14083), .ZN(n14087) );
NAND2_X2 U10952 ( .A1(n13096), .A2(n14085), .ZN(n14086) );
MUX2_X2 U10953 ( .A(n14087), .B(n14086), .S(n445), .Z(n14088) );
NAND2_X2 U10954 ( .A1(n14089), .A2(n14088), .ZN(SHA1_ft_BCD[30]) );
MUX2_X2 U10955 ( .A(n13159), .B(n13162), .S(next_C[27]), .Z(n14090) );
NAND2_X2 U10956 ( .A1(n14090), .A2(SHA1_result[61]), .ZN(n14097) );
XOR2_X2 U10957 ( .A(SHA1_result[61]), .B(next_C[27]), .Z(n14093) );
NOR2_X2 U10958 ( .A1(n14092), .A2(n14091), .ZN(n14095) );
NAND2_X2 U10959 ( .A1(n13096), .A2(n14093), .ZN(n14094) );
MUX2_X2 U10960 ( .A(n14095), .B(n14094), .S(n446), .Z(n14096) );
NAND2_X2 U10961 ( .A1(n14097), .A2(n14096), .ZN(SHA1_ft_BCD[29]) );
MUX2_X2 U10962 ( .A(n13158), .B(n13163), .S(next_C[26]), .Z(n14098) );
NAND2_X2 U10963 ( .A1(n14098), .A2(SHA1_result[60]), .ZN(n14105) );
XOR2_X2 U10964 ( .A(SHA1_result[60]), .B(next_C[26]), .Z(n14101) );
NOR2_X2 U10965 ( .A1(n14100), .A2(n14099), .ZN(n14103) );
NAND2_X2 U10966 ( .A1(n13096), .A2(n14101), .ZN(n14102) );
MUX2_X2 U10967 ( .A(n14103), .B(n14102), .S(n447), .Z(n14104) );
NAND2_X2 U10968 ( .A1(n14105), .A2(n14104), .ZN(SHA1_ft_BCD[28]) );
MUX2_X2 U10969 ( .A(n13158), .B(n13163), .S(next_C[25]), .Z(n14106) );
NAND2_X2 U10970 ( .A1(n14106), .A2(SHA1_result[59]), .ZN(n14113) );
NOR2_X2 U10971 ( .A1(n13082), .A2(n13008), .ZN(n14108) );
XOR2_X2 U10972 ( .A(SHA1_result[59]), .B(next_C[25]), .Z(n14109) );
NOR2_X2 U10973 ( .A1(n14108), .A2(n14107), .ZN(n14111) );
NAND2_X2 U10974 ( .A1(n13096), .A2(n14109), .ZN(n14110) );
MUX2_X2 U10975 ( .A(n14111), .B(n14110), .S(n448), .Z(n14112) );
NAND2_X2 U10976 ( .A1(n14113), .A2(n14112), .ZN(SHA1_ft_BCD[27]) );
MUX2_X2 U10977 ( .A(n13159), .B(n13164), .S(next_C[24]), .Z(n14114) );
NAND2_X2 U10978 ( .A1(n14114), .A2(SHA1_result[58]), .ZN(n14121) );
NOR2_X2 U10979 ( .A1(n13161), .A2(n13003), .ZN(n14116) );
XOR2_X2 U10980 ( .A(SHA1_result[58]), .B(next_C[24]), .Z(n14117) );
NOR2_X2 U10981 ( .A1(n14116), .A2(n14115), .ZN(n14119) );
NAND2_X2 U10982 ( .A1(n14174), .A2(n14117), .ZN(n14118) );
MUX2_X2 U10983 ( .A(n14119), .B(n14118), .S(n449), .Z(n14120) );
NAND2_X2 U10984 ( .A1(n14121), .A2(n14120), .ZN(SHA1_ft_BCD[26]) );
MUX2_X2 U10985 ( .A(n13158), .B(n13163), .S(next_C[23]), .Z(n14122) );
NAND2_X2 U10986 ( .A1(n14122), .A2(SHA1_result[57]), .ZN(n14129) );
NOR2_X2 U10987 ( .A1(n13161), .A2(n13009), .ZN(n14124) );
XOR2_X2 U10988 ( .A(SHA1_result[57]), .B(next_C[23]), .Z(n14125) );
NOR2_X2 U10989 ( .A1(n14124), .A2(n14123), .ZN(n14127) );
NAND2_X2 U10990 ( .A1(n14174), .A2(n14125), .ZN(n14126) );
MUX2_X2 U10991 ( .A(n14127), .B(n14126), .S(n450), .Z(n14128) );
NAND2_X2 U10992 ( .A1(n14129), .A2(n14128), .ZN(SHA1_ft_BCD[25]) );
MUX2_X2 U10993 ( .A(n13158), .B(n13162), .S(next_C[22]), .Z(n14130) );
NAND2_X2 U10994 ( .A1(n14130), .A2(SHA1_result[56]), .ZN(n14137) );
NOR2_X2 U10995 ( .A1(n13161), .A2(n13010), .ZN(n14132) );
XOR2_X2 U10996 ( .A(SHA1_result[56]), .B(next_C[22]), .Z(n14133) );
NOR2_X2 U10997 ( .A1(n14132), .A2(n14131), .ZN(n14135) );
NAND2_X2 U10998 ( .A1(n14174), .A2(n14133), .ZN(n14134) );
MUX2_X2 U10999 ( .A(n14135), .B(n14134), .S(n451), .Z(n14136) );
NAND2_X2 U11000 ( .A1(n14137), .A2(n14136), .ZN(SHA1_ft_BCD[24]) );
MUX2_X2 U11001 ( .A(n13158), .B(n13163), .S(next_C[21]), .Z(n14138) );
NAND2_X2 U11002 ( .A1(n14138), .A2(SHA1_result[55]), .ZN(n14145) );
NOR2_X2 U11003 ( .A1(n13161), .A2(n14680), .ZN(n14140) );
XOR2_X2 U11004 ( .A(SHA1_result[55]), .B(next_C[21]), .Z(n14141) );
NOR2_X2 U11005 ( .A1(n14140), .A2(n14139), .ZN(n14143) );
NAND2_X2 U11006 ( .A1(n14174), .A2(n14141), .ZN(n14142) );
MUX2_X2 U11007 ( .A(n14143), .B(n14142), .S(n452), .Z(n14144) );
NAND2_X2 U11008 ( .A1(n14145), .A2(n14144), .ZN(SHA1_ft_BCD[23]) );
MUX2_X2 U11009 ( .A(n13159), .B(n13164), .S(next_C[20]), .Z(n14146) );
NAND2_X2 U11010 ( .A1(n14146), .A2(n14681), .ZN(n14153) );
NOR2_X2 U11011 ( .A1(n13161), .A2(n13006), .ZN(n14148) );
XOR2_X2 U11012 ( .A(n14681), .B(next_C[20]), .Z(n14149) );
NOR2_X2 U11013 ( .A1(n14148), .A2(n14147), .ZN(n14151) );
MUX2_X2 U11014 ( .A(n14151), .B(n14150), .S(n453), .Z(n14152) );
NAND2_X2 U11015 ( .A1(n14153), .A2(n14152), .ZN(SHA1_ft_BCD[22]) );
MUX2_X2 U11016 ( .A(n13159), .B(n13162), .S(next_C[19]), .Z(n14154) );
NAND2_X2 U11017 ( .A1(n14154), .A2(n14682), .ZN(n14161) );
NOR2_X2 U11018 ( .A1(n13161), .A2(n13011), .ZN(n14156) );
XOR2_X2 U11019 ( .A(n14682), .B(next_C[19]), .Z(n14157) );
NOR2_X2 U11020 ( .A1(n14156), .A2(n14155), .ZN(n14159) );
MUX2_X2 U11021 ( .A(n14159), .B(n14158), .S(n454), .Z(n14160) );
NAND2_X2 U11022 ( .A1(n14161), .A2(n14160), .ZN(SHA1_ft_BCD[21]) );
MUX2_X2 U11023 ( .A(n13159), .B(n13164), .S(next_C[18]), .Z(n14162) );
NAND2_X2 U11024 ( .A1(n14162), .A2(n14868), .ZN(n14169) );
NOR2_X2 U11025 ( .A1(n13161), .A2(n13012), .ZN(n14164) );
XOR2_X2 U11026 ( .A(n14868), .B(next_C[18]), .Z(n14165) );
NOR2_X2 U11027 ( .A1(n14164), .A2(n14163), .ZN(n14167) );
MUX2_X2 U11028 ( .A(n14167), .B(n14166), .S(n455), .Z(n14168) );
MUX2_X2 U11029 ( .A(n13159), .B(n13162), .S(next_C[17]), .Z(n14170) );
NAND2_X2 U11030 ( .A1(n14170), .A2(SHA1_result[51]), .ZN(n14178) );
NOR2_X2 U11031 ( .A1(n13161), .A2(n14861), .ZN(n14172) );
XOR2_X2 U11032 ( .A(SHA1_result[51]), .B(next_C[17]), .Z(n14173) );
NOR2_X2 U11033 ( .A1(n14172), .A2(n14171), .ZN(n14176) );
MUX2_X2 U11034 ( .A(n14176), .B(n14175), .S(n456), .Z(n14177) );
NAND2_X2 U11035 ( .A1(n14178), .A2(n14177), .ZN(SHA1_ft_BCD[19]) );
MUX2_X2 U11036 ( .A(n13158), .B(n13162), .S(next_C[16]), .Z(n14179) );
NAND2_X2 U11037 ( .A1(n14179), .A2(SHA1_result[50]), .ZN(n14186) );
NOR2_X2 U11038 ( .A1(n13161), .A2(n13004), .ZN(n14181) );
XOR2_X2 U11039 ( .A(SHA1_result[50]), .B(next_C[16]), .Z(n14182) );
NOR2_X2 U11040 ( .A1(n14181), .A2(n14180), .ZN(n14184) );
NAND2_X2 U11041 ( .A1(n14368), .A2(n14182), .ZN(n14183) );
MUX2_X2 U11042 ( .A(n14184), .B(n14183), .S(n457), .Z(n14185) );
XOR2_X2 U11043 ( .A(SHA1_result[49]), .B(next_C[15]), .Z(n14187) );
NAND3_X2 U11044 ( .A1(n14368), .A2(n14187), .A3(n458), .ZN(n14197) );
NAND2_X2 U11045 ( .A1(n14187), .A2(n13117), .ZN(n14190) );
INV_X4 U11046 ( .A(n14187), .ZN(n14188) );
NAND2_X2 U11047 ( .A1(n14188), .A2(n13147), .ZN(n14189) );
NAND2_X2 U11048 ( .A1(n14190), .A2(n14189), .ZN(n14192) );
NAND2_X2 U11049 ( .A1(n14192), .A2(n14191), .ZN(n14193) );
NAND2_X2 U11050 ( .A1(n14193), .A2(SHA1_result[81]), .ZN(n14196) );
MUX2_X2 U11051 ( .A(n13158), .B(n13164), .S(next_C[15]), .Z(n14194) );
NAND2_X2 U11052 ( .A1(n14194), .A2(SHA1_result[49]), .ZN(n14195) );
XOR2_X2 U11053 ( .A(SHA1_result[48]), .B(next_C[14]), .Z(n14201) );
NAND3_X2 U11054 ( .A1(n14368), .A2(n14201), .A3(n459), .ZN(n14207) );
INV_X4 U11055 ( .A(n14201), .ZN(n14199) );
NAND2_X2 U11056 ( .A1(next_C[14]), .A2(n13158), .ZN(n14200) );
NAND3_X2 U11057 ( .A1(n14199), .A2(n13147), .A3(n14200), .ZN(n14203) );
NAND3_X2 U11058 ( .A1(n14201), .A2(n13117), .A3(n14200), .ZN(n14202) );
NAND3_X2 U11059 ( .A1(n14203), .A2(SHA1_result[80]), .A3(n14202), .ZN(n14206) );
MUX2_X2 U11060 ( .A(n13159), .B(n13162), .S(next_C[14]), .Z(n14204) );
NAND2_X2 U11061 ( .A1(n14204), .A2(SHA1_result[48]), .ZN(n14205) );
NAND3_X2 U11062 ( .A1(n14207), .A2(n14206), .A3(n14205), .ZN(SHA1_ft_BCD[16]) );
NAND2_X2 U11063 ( .A1(next_C[13]), .A2(n14334), .ZN(n14209) );
XOR2_X2 U11064 ( .A(SHA1_result[47]), .B(next_C[13]), .Z(n14212) );
INV_X4 U11065 ( .A(n14212), .ZN(n14208) );
NAND3_X2 U11066 ( .A1(n14209), .A2(n14208), .A3(n14356), .ZN(n14211) );
NAND3_X2 U11067 ( .A1(n14212), .A2(n14209), .A3(n13117), .ZN(n14210) );
NAND3_X2 U11068 ( .A1(n14211), .A2(SHA1_result[79]), .A3(n14210), .ZN(n14217) );
NAND3_X2 U11069 ( .A1(n460), .A2(n14368), .A3(n14212), .ZN(n14216) );
MUX2_X2 U11070 ( .A(n13142), .B(n14330), .S(next_C[13]), .Z(n14214) );
NAND2_X2 U11071 ( .A1(n14214), .A2(SHA1_result[47]), .ZN(n14215) );
NAND3_X2 U11072 ( .A1(n14217), .A2(n14216), .A3(n14215), .ZN(SHA1_ft_BCD[15]) );
NAND2_X2 U11073 ( .A1(n13161), .A2(n13005), .ZN(n14219) );
NAND3_X2 U11074 ( .A1(n14219), .A2(n14830), .A3(n14218), .ZN(n14225) );
XOR2_X2 U11075 ( .A(n14830), .B(next_C[12]), .Z(n14220) );
NAND2_X2 U11076 ( .A1(n14368), .A2(n14221), .ZN(n14222) );
MUX2_X2 U11077 ( .A(n13142), .B(n14330), .S(next_C[11]), .Z(n14226) );
NAND2_X2 U11078 ( .A1(n14226), .A2(SHA1_result[45]), .ZN(n14234) );
XOR2_X2 U11079 ( .A(SHA1_result[45]), .B(next_C[11]), .Z(n14227) );
NAND3_X2 U11080 ( .A1(n462), .A2(n14368), .A3(n14227), .ZN(n14233) );
NAND2_X2 U11081 ( .A1(next_C[11]), .A2(n14334), .ZN(n14229) );
NAND3_X2 U11082 ( .A1(n14227), .A2(n14229), .A3(n13165), .ZN(n14231) );
INV_X4 U11083 ( .A(n14227), .ZN(n14228) );
NAND3_X2 U11084 ( .A1(n14229), .A2(n14228), .A3(n13147), .ZN(n14230) );
NAND3_X2 U11085 ( .A1(n14231), .A2(SHA1_result[77]), .A3(n14230), .ZN(n14232) );
NAND2_X2 U11086 ( .A1(next_C[10]), .A2(n13157), .ZN(n14235) );
XOR2_X2 U11087 ( .A(n14817), .B(next_C[10]), .Z(n14239) );
NAND3_X2 U11088 ( .A1(n14235), .A2(n13117), .A3(n14239), .ZN(n14238) );
INV_X4 U11089 ( .A(n14239), .ZN(n14236) );
NAND3_X2 U11090 ( .A1(n14236), .A2(n13147), .A3(n14235), .ZN(n14237) );
NAND3_X2 U11091 ( .A1(n14238), .A2(SHA1_result[76]), .A3(n14237), .ZN(n14243) );
MUX2_X2 U11092 ( .A(n13159), .B(n13162), .S(next_C[10]), .Z(n14240) );
XOR2_X2 U11093 ( .A(n14810), .B(next_C[9]), .Z(n14246) );
NAND3_X2 U11094 ( .A1(n464), .A2(n14368), .A3(n14246), .ZN(n14253) );
NAND2_X2 U11095 ( .A1(n13161), .A2(n13001), .ZN(n14245) );
NAND2_X2 U11096 ( .A1(next_C[9]), .A2(n13117), .ZN(n14244) );
NAND3_X2 U11097 ( .A1(n14245), .A2(n14810), .A3(n14244), .ZN(n14252) );
NAND2_X2 U11098 ( .A1(next_C[9]), .A2(n13157), .ZN(n14248) );
NAND3_X2 U11099 ( .A1(n14248), .A2(n13117), .A3(n14246), .ZN(n14250) );
INV_X4 U11100 ( .A(n14246), .ZN(n14247) );
NAND3_X2 U11101 ( .A1(n14248), .A2(n13074), .A3(n14247), .ZN(n14249) );
NAND3_X2 U11102 ( .A1(n14250), .A2(SHA1_result[75]), .A3(n14249), .ZN(n14251) );
NAND3_X2 U11103 ( .A1(n14253), .A2(n14252), .A3(n14251), .ZN(SHA1_ft_BCD[11]) );
XOR2_X2 U11104 ( .A(SHA1_result[42]), .B(next_C[8]), .Z(n14263) );
NAND2_X2 U11105 ( .A1(n14255), .A2(SHA1_result[74]), .ZN(n14258) );
NOR2_X2 U11106 ( .A1(n14331), .A2(n13098), .ZN(n14257) );
NOR2_X2 U11107 ( .A1(next_C[8]), .A2(n13157), .ZN(n14256) );
NOR2_X2 U11108 ( .A1(n13090), .A2(n14258), .ZN(n14259) );
XOR2_X2 U11109 ( .A(n14797), .B(next_C[7]), .Z(n14270) );
NAND3_X2 U11110 ( .A1(n466), .A2(n14270), .A3(n14368), .ZN(n14277) );
NAND2_X2 U11111 ( .A1(n13075), .A2(n13088), .ZN(n14342) );
INV_X4 U11112 ( .A(n14270), .ZN(n14268) );
NAND3_X2 U11113 ( .A1(n14269), .A2(n14344), .A3(n14268), .ZN(n14272) );
NAND3_X2 U11114 ( .A1(n14271), .A2(SHA1_result[73]), .A3(n14272), .ZN(n14276) );
NAND2_X2 U11115 ( .A1(n14274), .A2(n14797), .ZN(n14275) );
NAND3_X2 U11116 ( .A1(n14275), .A2(n14277), .A3(n14276), .ZN(SHA1_ft_BCD[9]));
XOR2_X2 U11117 ( .A(SHA1_result[40]), .B(next_C[6]), .Z(n14284) );
INV_X4 U11118 ( .A(n14284), .ZN(n14281) );
NAND3_X2 U11119 ( .A1(n14283), .A2(SHA1_result[72]), .A3(n14282), .ZN(n14288) );
NAND3_X2 U11120 ( .A1(n467), .A2(n14349), .A3(n14284), .ZN(n14287) );
MUX2_X2 U11121 ( .A(n13142), .B(n14331), .S(next_C[6]), .Z(n14285) );
NAND2_X2 U11122 ( .A1(n14285), .A2(SHA1_result[40]), .ZN(n14286) );
NAND3_X2 U11123 ( .A1(n14288), .A2(n14286), .A3(n14287), .ZN(SHA1_ft_BCD[8]));
NAND2_X2 U11124 ( .A1(next_C[5]), .A2(n14334), .ZN(n14290) );
XOR2_X2 U11125 ( .A(SHA1_result[39]), .B(next_C[5]), .Z(n14293) );
INV_X4 U11126 ( .A(n14293), .ZN(n14289) );
NAND3_X2 U11127 ( .A1(n14290), .A2(n14289), .A3(n13147), .ZN(n14292) );
NAND3_X2 U11128 ( .A1(n14293), .A2(n14290), .A3(n13117), .ZN(n14291) );
NAND3_X2 U11129 ( .A1(n14292), .A2(SHA1_result[71]), .A3(n14291), .ZN(n14297) );
NAND3_X2 U11130 ( .A1(n468), .A2(n14368), .A3(n14293), .ZN(n14296) );
NAND2_X2 U11131 ( .A1(n14294), .A2(SHA1_result[39]), .ZN(n14295) );
XOR2_X2 U11132 ( .A(n14778), .B(next_C[4]), .Z(n14298) );
NAND3_X2 U11133 ( .A1(n14298), .A2(SHA1_result[70]), .A3(n13162), .ZN(n14306) );
INV_X4 U11134 ( .A(n14298), .ZN(n14299) );
NAND3_X2 U11135 ( .A1(n14299), .A2(SHA1_result[70]), .A3(n14349), .ZN(n14304) );
NOR3_X2 U11136 ( .A1(n437), .A2(n13099), .A3(n13000), .ZN(n14302) );
NOR3_X2 U11137 ( .A1(n14344), .A2(n14299), .A3(SHA1_result[70]), .ZN(n14301));
NAND3_X2 U11138 ( .A1(n14770), .A2(n14771), .A3(n13158), .ZN(n14319) );
XOR2_X2 U11139 ( .A(n14770), .B(next_C[3]), .Z(n14310) );
NAND2_X2 U11140 ( .A1(n470), .A2(n14310), .ZN(n14308) );
INV_X4 U11141 ( .A(n14310), .ZN(n14307) );
NAND2_X2 U11142 ( .A1(n14307), .A2(SHA1_result[69]), .ZN(n14313) );
NAND2_X2 U11143 ( .A1(n14308), .A2(n14313), .ZN(n14309) );
NAND2_X2 U11144 ( .A1(n14310), .A2(SHA1_result[69]), .ZN(n14314) );
NAND2_X2 U11145 ( .A1(n14311), .A2(n14314), .ZN(n14312) );
NAND2_X2 U11146 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
XOR2_X2 U11147 ( .A(SHA1_result[36]), .B(next_C[2]), .Z(n14323) );
NAND3_X2 U11148 ( .A1(n471), .A2(n14323), .A3(n14368), .ZN(n14329) );
INV_X4 U11149 ( .A(n14323), .ZN(n14320) );
NAND3_X2 U11150 ( .A1(n14323), .A2(n14322), .A3(n13117), .ZN(n14324) );
NAND3_X2 U11151 ( .A1(n14324), .A2(SHA1_result[68]), .A3(n14325), .ZN(n14328) );
NAND2_X2 U11152 ( .A1(n14326), .A2(SHA1_result[36]), .ZN(n14327) );
XOR2_X2 U11153 ( .A(SHA1_result[35]), .B(next_C[1]), .Z(n14332) );
INV_X4 U11154 ( .A(n14332), .ZN(n14333) );
NAND3_X2 U11155 ( .A1(n14333), .A2(SHA1_result[67]), .A3(n14349), .ZN(n14341) );
NAND3_X2 U11156 ( .A1(next_C[1]), .A2(SHA1_result[35]), .A3(n14330), .ZN(n14340) );
NOR3_X2 U11157 ( .A1(n472), .A2(n14360), .A3(n14757), .ZN(n14336) );
XOR2_X2 U11158 ( .A(SHA1_result[34]), .B(next_C[0]), .Z(n14348) );
INV_X4 U11159 ( .A(n14348), .ZN(n14345) );
INV_X4 U11160 ( .A(next_C[0]), .ZN(n14750) );
NAND3_X2 U11161 ( .A1(n14345), .A2(n14750), .A3(n14356), .ZN(n14346) );
NAND3_X2 U11162 ( .A1(n14347), .A2(SHA1_result[66]), .A3(n14346), .ZN(n14355) );
NAND3_X2 U11163 ( .A1(n473), .A2(n14349), .A3(n14348), .ZN(n14354) );
NOR3_X2 U11164 ( .A1(n14371), .A2(n474), .A3(n14365), .ZN(n14364) );
NOR2_X2 U11165 ( .A1(n442), .A2(n14743), .ZN(n14358) );
NOR2_X2 U11166 ( .A1(n14358), .A2(n14357), .ZN(n14359) );
NOR3_X2 U11167 ( .A1(n474), .A2(n14360), .A3(n14743), .ZN(n14361) );
NOR4_X2 U11168 ( .A1(n14364), .A2(n14363), .A3(n14362), .A4(n14361), .ZN(n14367) );
XOR2_X2 U11169 ( .A(n13084), .B(n443), .Z(n14370) );
NAND3_X2 U11170 ( .A1(n475), .A2(n14370), .A3(n14368), .ZN(n14379) );
INV_X4 U11171 ( .A(n14370), .ZN(n14372) );
NAND3_X2 U11172 ( .A1(n14374), .A2(SHA1_result[64]), .A3(n14373), .ZN(n14378) );
NAND3_X2 U11173 ( .A1(n14377), .A2(n14378), .A3(n14379), .ZN(SHA1_ft_BCD[0]));
NAND2_X2 U11174 ( .A1(n13194), .A2(n14464), .ZN(n14381) );
NAND2_X2 U11175 ( .A1(H0[31]), .A2(n13327), .ZN(n14380) );
NAND2_X2 U11176 ( .A1(n14381), .A2(n14380), .ZN(n3953) );
NAND2_X2 U11177 ( .A1(H0[30]), .A2(n13327), .ZN(n14384) );
NAND2_X2 U11178 ( .A1(n13345), .A2(n14382), .ZN(n14383) );
NAND3_X2 U11179 ( .A1(n14384), .A2(n13191), .A3(n14383), .ZN(n3954) );
NAND2_X2 U11180 ( .A1(H0[29]), .A2(n13327), .ZN(n14387) );
NAND2_X2 U11181 ( .A1(n13345), .A2(n14385), .ZN(n14386) );
NAND3_X2 U11182 ( .A1(n14387), .A2(n13191), .A3(n14386), .ZN(n3955) );
NAND2_X2 U11183 ( .A1(n13194), .A2(n14388), .ZN(n14390) );
NAND2_X2 U11184 ( .A1(H0[28]), .A2(n13327), .ZN(n14389) );
NAND2_X2 U11185 ( .A1(n14390), .A2(n14389), .ZN(n3956) );
NAND2_X2 U11186 ( .A1(n13194), .A2(n14391), .ZN(n14393) );
NAND2_X2 U11187 ( .A1(H0[27]), .A2(n13327), .ZN(n14392) );
NAND2_X2 U11188 ( .A1(n14393), .A2(n14392), .ZN(n3957) );
NAND2_X2 U11189 ( .A1(H0[26]), .A2(n13327), .ZN(n14396) );
NAND2_X2 U11190 ( .A1(n13345), .A2(n14394), .ZN(n14395) );
NAND3_X2 U11191 ( .A1(n14396), .A2(n13191), .A3(n14395), .ZN(n3958) );
NAND2_X2 U11192 ( .A1(H0[25]), .A2(n13327), .ZN(n14399) );
NAND2_X2 U11193 ( .A1(n13345), .A2(n14397), .ZN(n14398) );
NAND3_X2 U11194 ( .A1(n14399), .A2(n13191), .A3(n14398), .ZN(n3959) );
NAND2_X2 U11195 ( .A1(H0[24]), .A2(n13327), .ZN(n14402) );
NAND2_X2 U11196 ( .A1(n13346), .A2(n14400), .ZN(n14401) );
NAND3_X2 U11197 ( .A1(n14402), .A2(n13191), .A3(n14401), .ZN(n3960) );
NAND2_X2 U11198 ( .A1(n13194), .A2(SHA1_result_151), .ZN(n14404) );
NAND2_X2 U11199 ( .A1(H0[23]), .A2(n13327), .ZN(n14403) );
NAND2_X2 U11200 ( .A1(n14404), .A2(n14403), .ZN(n3961) );
NAND2_X2 U11201 ( .A1(H0[22]), .A2(n13327), .ZN(n14407) );
NAND2_X2 U11202 ( .A1(n13346), .A2(n14405), .ZN(n14406) );
NAND3_X2 U11203 ( .A1(n14407), .A2(n13191), .A3(n14406), .ZN(n3962) );
NAND2_X2 U11204 ( .A1(n13194), .A2(n14408), .ZN(n14410) );
NAND2_X2 U11205 ( .A1(H0[21]), .A2(n13327), .ZN(n14409) );
NAND2_X2 U11206 ( .A1(n14410), .A2(n14409), .ZN(n3963) );
NAND2_X2 U11207 ( .A1(n13194), .A2(SHA1_result_148), .ZN(n14412) );
NAND2_X2 U11208 ( .A1(H0[20]), .A2(n13327), .ZN(n14411) );
NAND2_X2 U11209 ( .A1(n14412), .A2(n14411), .ZN(n3964) );
NAND2_X2 U11210 ( .A1(n13195), .A2(n14413), .ZN(n14415) );
NAND2_X2 U11211 ( .A1(H0[19]), .A2(n13327), .ZN(n14414) );
NAND2_X2 U11212 ( .A1(n14415), .A2(n14414), .ZN(n3965) );
NAND2_X2 U11213 ( .A1(H0[18]), .A2(n13327), .ZN(n14418) );
NAND2_X2 U11214 ( .A1(n13346), .A2(n14416), .ZN(n14417) );
NAND3_X2 U11215 ( .A1(n14418), .A2(n13191), .A3(n14417), .ZN(n3966) );
NAND2_X2 U11216 ( .A1(n13195), .A2(n14419), .ZN(n14421) );
NAND2_X2 U11217 ( .A1(H0[17]), .A2(n13327), .ZN(n14420) );
NAND2_X2 U11218 ( .A1(n14421), .A2(n14420), .ZN(n3967) );
NAND2_X2 U11219 ( .A1(H0[16]), .A2(n13327), .ZN(n14424) );
NAND2_X2 U11220 ( .A1(n13346), .A2(n14422), .ZN(n14423) );
NAND3_X2 U11221 ( .A1(n14424), .A2(n13191), .A3(n14423), .ZN(n3968) );
NAND2_X2 U11222 ( .A1(n13195), .A2(n14425), .ZN(n14427) );
NAND2_X2 U11223 ( .A1(H0[15]), .A2(n13326), .ZN(n14426) );
NAND2_X2 U11224 ( .A1(n14427), .A2(n14426), .ZN(n3969) );
NAND2_X2 U11225 ( .A1(n13195), .A2(n14428), .ZN(n14430) );
NAND2_X2 U11226 ( .A1(H0[14]), .A2(n13326), .ZN(n14429) );
NAND2_X2 U11227 ( .A1(n14430), .A2(n14429), .ZN(n3970) );
NAND2_X2 U11228 ( .A1(H0[13]), .A2(n13326), .ZN(n14433) );
NAND2_X2 U11229 ( .A1(n13346), .A2(n14431), .ZN(n14432) );
NAND3_X2 U11230 ( .A1(n14433), .A2(n13191), .A3(n14432), .ZN(n3971) );
NAND2_X2 U11231 ( .A1(n13195), .A2(n14434), .ZN(n14436) );
NAND2_X2 U11232 ( .A1(H0[12]), .A2(n13326), .ZN(n14435) );
NAND2_X2 U11233 ( .A1(n14436), .A2(n14435), .ZN(n3972) );
NAND2_X2 U11234 ( .A1(n13195), .A2(n14437), .ZN(n14439) );
NAND2_X2 U11235 ( .A1(H0[11]), .A2(n13326), .ZN(n14438) );
NAND2_X2 U11236 ( .A1(n14439), .A2(n14438), .ZN(n3973) );
NAND2_X2 U11237 ( .A1(n13195), .A2(n14440), .ZN(n14442) );
NAND2_X2 U11238 ( .A1(H0[10]), .A2(n13326), .ZN(n14441) );
NAND2_X2 U11239 ( .A1(n14442), .A2(n14441), .ZN(n3974) );
NAND2_X2 U11240 ( .A1(H0[9]), .A2(n13326), .ZN(n14445) );
NAND2_X2 U11241 ( .A1(n13346), .A2(n14443), .ZN(n14444) );
NAND3_X2 U11242 ( .A1(n14445), .A2(n13191), .A3(n14444), .ZN(n3975) );
NAND2_X2 U11243 ( .A1(H0[8]), .A2(n13326), .ZN(n14447) );
NAND2_X2 U11244 ( .A1(n13346), .A2(SHA1_result_136), .ZN(n14446) );
NAND3_X2 U11245 ( .A1(n14447), .A2(n13190), .A3(n14446), .ZN(n3976) );
NAND2_X2 U11246 ( .A1(n13195), .A2(SHA1_result_135), .ZN(n14449) );
NAND2_X2 U11247 ( .A1(H0[7]), .A2(n13326), .ZN(n14448) );
NAND2_X2 U11248 ( .A1(n14449), .A2(n14448), .ZN(n3977) );
NAND2_X2 U11249 ( .A1(n13195), .A2(SHA1_result_134), .ZN(n14451) );
NAND2_X2 U11250 ( .A1(H0[6]), .A2(n13326), .ZN(n14450) );
NAND2_X2 U11251 ( .A1(n14451), .A2(n14450), .ZN(n3978) );
NAND2_X2 U11252 ( .A1(n13195), .A2(SHA1_result_133), .ZN(n14453) );
NAND2_X2 U11253 ( .A1(H0[5]), .A2(n13326), .ZN(n14452) );
NAND2_X2 U11254 ( .A1(n14453), .A2(n14452), .ZN(n3979) );
NAND2_X2 U11255 ( .A1(n13195), .A2(SHA1_result_132), .ZN(n14455) );
NAND2_X2 U11256 ( .A1(H0[4]), .A2(n13326), .ZN(n14454) );
NAND2_X2 U11257 ( .A1(n14455), .A2(n14454), .ZN(n3980) );
NAND2_X2 U11258 ( .A1(n13196), .A2(SHA1_result_131), .ZN(n14457) );
NAND2_X2 U11259 ( .A1(H0[3]), .A2(n13326), .ZN(n14456) );
NAND2_X2 U11260 ( .A1(n14457), .A2(n14456), .ZN(n3981) );
NAND2_X2 U11261 ( .A1(n13196), .A2(SHA1_result_130), .ZN(n14459) );
NAND2_X2 U11262 ( .A1(H0[2]), .A2(n13326), .ZN(n14458) );
NAND2_X2 U11263 ( .A1(n14459), .A2(n14458), .ZN(n3982) );
NAND2_X2 U11264 ( .A1(n13196), .A2(SHA1_result_129), .ZN(n14461) );
NAND2_X2 U11265 ( .A1(H0[1]), .A2(n13326), .ZN(n14460) );
NAND2_X2 U11266 ( .A1(n14461), .A2(n14460), .ZN(n3983) );
NAND2_X2 U11267 ( .A1(n13346), .A2(SHA1_result_128), .ZN(n14463) );
NAND2_X2 U11268 ( .A1(H0[0]), .A2(n13326), .ZN(n14462) );
NAND3_X2 U11269 ( .A1(n14463), .A2(n14462), .A3(n13186), .ZN(n3984) );
NAND2_X2 U11270 ( .A1(n13214), .A2(n14464), .ZN(n14467) );
NAND2_X2 U11271 ( .A1(next_A[31]), .A2(n13206), .ZN(n14466) );
NAND2_X2 U11272 ( .A1(N883), .A2(n13209), .ZN(n14465) );
NAND3_X2 U11273 ( .A1(n14465), .A2(n14466), .A3(n14467), .ZN(n3985) );
NAND2_X2 U11274 ( .A1(H1[31]), .A2(n13326), .ZN(n14469) );
NAND2_X2 U11275 ( .A1(n13346), .A2(next_C[29]), .ZN(n14468) );
NAND3_X2 U11276 ( .A1(n14469), .A2(n13190), .A3(n14468), .ZN(n3697) );
NAND2_X2 U11277 ( .A1(H1[30]), .A2(n13326), .ZN(n14471) );
NAND2_X2 U11278 ( .A1(n13346), .A2(next_C[28]), .ZN(n14470) );
NAND3_X2 U11279 ( .A1(n14471), .A2(n13190), .A3(n14470), .ZN(n3698) );
NAND2_X2 U11280 ( .A1(H1[29]), .A2(n13326), .ZN(n14473) );
NAND2_X2 U11281 ( .A1(n13346), .A2(next_C[27]), .ZN(n14472) );
NAND3_X2 U11282 ( .A1(n14473), .A2(n13190), .A3(n14472), .ZN(n3699) );
NAND2_X2 U11283 ( .A1(n13196), .A2(next_C[26]), .ZN(n14475) );
NAND2_X2 U11284 ( .A1(H1[28]), .A2(n13325), .ZN(n14474) );
NAND2_X2 U11285 ( .A1(n14475), .A2(n14474), .ZN(n3700) );
NAND2_X2 U11286 ( .A1(H1[27]), .A2(n13325), .ZN(n14477) );
NAND2_X2 U11287 ( .A1(n13347), .A2(next_C[25]), .ZN(n14476) );
NAND3_X2 U11288 ( .A1(n14477), .A2(n13190), .A3(n14476), .ZN(n3701) );
NAND2_X2 U11289 ( .A1(H1[26]), .A2(n13325), .ZN(n14479) );
NAND2_X2 U11290 ( .A1(n13347), .A2(next_C[24]), .ZN(n14478) );
NAND3_X2 U11291 ( .A1(n14479), .A2(n13190), .A3(n14478), .ZN(n3702) );
NAND2_X2 U11292 ( .A1(H1[25]), .A2(n13325), .ZN(n14481) );
NAND2_X2 U11293 ( .A1(n13347), .A2(next_C[23]), .ZN(n14480) );
NAND3_X2 U11294 ( .A1(n14481), .A2(n13190), .A3(n14480), .ZN(n3703) );
NAND2_X2 U11295 ( .A1(H1[24]), .A2(n13325), .ZN(n14483) );
NAND2_X2 U11296 ( .A1(n13347), .A2(next_C[22]), .ZN(n14482) );
NAND3_X2 U11297 ( .A1(n14483), .A2(n13190), .A3(n14482), .ZN(n3704) );
NAND2_X2 U11298 ( .A1(H1[23]), .A2(n13325), .ZN(n14485) );
NAND2_X2 U11299 ( .A1(n13347), .A2(next_C[21]), .ZN(n14484) );
NAND3_X2 U11300 ( .A1(n14485), .A2(n13190), .A3(n14484), .ZN(n3705) );
NAND2_X2 U11301 ( .A1(H1[22]), .A2(n13325), .ZN(n14487) );
NAND2_X2 U11302 ( .A1(n13347), .A2(next_C[20]), .ZN(n14486) );
NAND3_X2 U11303 ( .A1(n14487), .A2(n13190), .A3(n14486), .ZN(n3706) );
NAND2_X2 U11304 ( .A1(n13196), .A2(next_C[19]), .ZN(n14489) );
NAND2_X2 U11305 ( .A1(H1[21]), .A2(n13325), .ZN(n14488) );
NAND2_X2 U11306 ( .A1(n14489), .A2(n14488), .ZN(n3707) );
NAND2_X2 U11307 ( .A1(n13196), .A2(next_C[18]), .ZN(n14491) );
NAND2_X2 U11308 ( .A1(H1[20]), .A2(n13325), .ZN(n14490) );
NAND2_X2 U11309 ( .A1(n14491), .A2(n14490), .ZN(n3708) );
NAND2_X2 U11310 ( .A1(H1[19]), .A2(n13325), .ZN(n14493) );
NAND2_X2 U11311 ( .A1(n13347), .A2(next_C[17]), .ZN(n14492) );
NAND3_X2 U11312 ( .A1(n14493), .A2(n13190), .A3(n14492), .ZN(n3709) );
NAND2_X2 U11313 ( .A1(H1[18]), .A2(n13325), .ZN(n14495) );
NAND2_X2 U11314 ( .A1(n13347), .A2(next_C[16]), .ZN(n14494) );
NAND3_X2 U11315 ( .A1(n14495), .A2(n13189), .A3(n14494), .ZN(n3710) );
NAND2_X2 U11316 ( .A1(n13196), .A2(next_C[15]), .ZN(n14497) );
NAND2_X2 U11317 ( .A1(H1[17]), .A2(n13325), .ZN(n14496) );
NAND2_X2 U11318 ( .A1(n14497), .A2(n14496), .ZN(n3711) );
NAND2_X2 U11319 ( .A1(H1[16]), .A2(n13325), .ZN(n14499) );
NAND2_X2 U11320 ( .A1(n13347), .A2(next_C[14]), .ZN(n14498) );
NAND3_X2 U11321 ( .A1(n14499), .A2(n13189), .A3(n14498), .ZN(n3712) );
NAND2_X2 U11322 ( .A1(H1[15]), .A2(n13325), .ZN(n14501) );
NAND2_X2 U11323 ( .A1(n13347), .A2(next_C[13]), .ZN(n14500) );
NAND3_X2 U11324 ( .A1(n14501), .A2(n13189), .A3(n14500), .ZN(n3713) );
NAND2_X2 U11325 ( .A1(n13196), .A2(next_C[12]), .ZN(n14503) );
NAND2_X2 U11326 ( .A1(H1[14]), .A2(n13325), .ZN(n14502) );
NAND2_X2 U11327 ( .A1(n14503), .A2(n14502), .ZN(n3714) );
NAND2_X2 U11328 ( .A1(H1[13]), .A2(n13325), .ZN(n14505) );
NAND2_X2 U11329 ( .A1(n13347), .A2(next_C[11]), .ZN(n14504) );
NAND3_X2 U11330 ( .A1(n14505), .A2(n13189), .A3(n14504), .ZN(n3715) );
NAND2_X2 U11331 ( .A1(n13196), .A2(next_C[10]), .ZN(n14507) );
NAND2_X2 U11332 ( .A1(H1[12]), .A2(n13325), .ZN(n14506) );
NAND2_X2 U11333 ( .A1(n14507), .A2(n14506), .ZN(n3716) );
NAND2_X2 U11334 ( .A1(H1[11]), .A2(n13325), .ZN(n14509) );
NAND2_X2 U11335 ( .A1(n13348), .A2(next_C[9]), .ZN(n14508) );
NAND3_X2 U11336 ( .A1(n14509), .A2(n13189), .A3(n14508), .ZN(n3717) );
NAND2_X2 U11337 ( .A1(n13196), .A2(next_C[8]), .ZN(n14511) );
NAND2_X2 U11338 ( .A1(H1[10]), .A2(n13325), .ZN(n14510) );
NAND2_X2 U11339 ( .A1(n14511), .A2(n14510), .ZN(n3718) );
NAND2_X2 U11340 ( .A1(H1[9]), .A2(n13324), .ZN(n14513) );
NAND2_X2 U11341 ( .A1(n13348), .A2(next_C[7]), .ZN(n14512) );
NAND3_X2 U11342 ( .A1(n14513), .A2(n13189), .A3(n14512), .ZN(n3719) );
NAND2_X2 U11343 ( .A1(H1[8]), .A2(n13324), .ZN(n14515) );
NAND2_X2 U11344 ( .A1(n13348), .A2(next_C[6]), .ZN(n14514) );
NAND3_X2 U11345 ( .A1(n14515), .A2(n13189), .A3(n14514), .ZN(n3720) );
NAND2_X2 U11346 ( .A1(H1[7]), .A2(n13324), .ZN(n14517) );
NAND2_X2 U11347 ( .A1(n13348), .A2(next_C[5]), .ZN(n14516) );
NAND3_X2 U11348 ( .A1(n14517), .A2(n13189), .A3(n14516), .ZN(n3721) );
NAND2_X2 U11349 ( .A1(n13196), .A2(next_C[4]), .ZN(n14519) );
NAND2_X2 U11350 ( .A1(H1[6]), .A2(n13324), .ZN(n14518) );
NAND2_X2 U11351 ( .A1(n14519), .A2(n14518), .ZN(n3722) );
NAND2_X2 U11352 ( .A1(H1[5]), .A2(n13324), .ZN(n14520) );
NAND2_X2 U11353 ( .A1(n14521), .A2(n14520), .ZN(n3723) );
NAND2_X2 U11354 ( .A1(n13197), .A2(next_C[2]), .ZN(n14523) );
NAND2_X2 U11355 ( .A1(H1[4]), .A2(n13324), .ZN(n14522) );
NAND2_X2 U11356 ( .A1(n14523), .A2(n14522), .ZN(n3724) );
NAND2_X2 U11357 ( .A1(H1[3]), .A2(n13324), .ZN(n14525) );
NAND2_X2 U11358 ( .A1(n13348), .A2(next_C[1]), .ZN(n14524) );
NAND3_X2 U11359 ( .A1(n14525), .A2(n13189), .A3(n14524), .ZN(n3725) );
NAND2_X2 U11360 ( .A1(n13197), .A2(next_C[0]), .ZN(n14527) );
NAND2_X2 U11361 ( .A1(H1[2]), .A2(n13324), .ZN(n14526) );
NAND2_X2 U11362 ( .A1(n14527), .A2(n14526), .ZN(n3726) );
NAND2_X2 U11363 ( .A1(H1[1]), .A2(n13324), .ZN(n14528) );
NAND2_X2 U11364 ( .A1(n14529), .A2(n14528), .ZN(n3727) );
NAND2_X2 U11365 ( .A1(H1[0]), .A2(n13324), .ZN(n14531) );
NAND2_X2 U11366 ( .A1(n13348), .A2(next_C[30]), .ZN(n14530) );
NAND3_X2 U11367 ( .A1(n14531), .A2(n13189), .A3(n14530), .ZN(n3728) );
NAND2_X2 U11368 ( .A1(N885), .A2(n13171), .ZN(n14534) );
NAND2_X2 U11369 ( .A1(n13177), .A2(SHA1_result_129), .ZN(n14532) );
NAND3_X2 U11370 ( .A1(n14534), .A2(n14533), .A3(n14532), .ZN(n3951) );
NAND2_X2 U11371 ( .A1(H2[31]), .A2(n13324), .ZN(n14536) );
NAND2_X2 U11372 ( .A1(n13348), .A2(SHA1_result[95]), .ZN(n14535) );
NAND3_X2 U11373 ( .A1(n14536), .A2(n13188), .A3(n14535), .ZN(n3729) );
NAND2_X2 U11374 ( .A1(n13197), .A2(SHA1_result[94]), .ZN(n14538) );
NAND2_X2 U11375 ( .A1(H2[30]), .A2(n13324), .ZN(n14537) );
NAND2_X2 U11376 ( .A1(n14538), .A2(n14537), .ZN(n3730) );
NAND2_X2 U11377 ( .A1(n13197), .A2(SHA1_result[93]), .ZN(n14540) );
NAND2_X2 U11378 ( .A1(H2[29]), .A2(n13324), .ZN(n14539) );
NAND2_X2 U11379 ( .A1(n14540), .A2(n14539), .ZN(n3731) );
NAND2_X2 U11380 ( .A1(H2[28]), .A2(n13324), .ZN(n14542) );
NAND2_X2 U11381 ( .A1(n13348), .A2(SHA1_result[92]), .ZN(n14541) );
NAND3_X2 U11382 ( .A1(n14542), .A2(n13188), .A3(n14541), .ZN(n3732) );
NAND2_X2 U11383 ( .A1(H2[27]), .A2(n13324), .ZN(n14544) );
NAND2_X2 U11384 ( .A1(n13348), .A2(SHA1_result[91]), .ZN(n14543) );
NAND3_X2 U11385 ( .A1(n14544), .A2(n13188), .A3(n14543), .ZN(n3733) );
NAND2_X2 U11386 ( .A1(n13197), .A2(SHA1_result[90]), .ZN(n14546) );
NAND2_X2 U11387 ( .A1(H2[26]), .A2(n13324), .ZN(n14545) );
NAND2_X2 U11388 ( .A1(n14546), .A2(n14545), .ZN(n3734) );
NAND2_X2 U11389 ( .A1(n13197), .A2(SHA1_result[89]), .ZN(n14548) );
NAND2_X2 U11390 ( .A1(H2[25]), .A2(n13324), .ZN(n14547) );
NAND2_X2 U11391 ( .A1(n14548), .A2(n14547), .ZN(n3735) );
NAND2_X2 U11392 ( .A1(n13197), .A2(SHA1_result[88]), .ZN(n14550) );
NAND2_X2 U11393 ( .A1(H2[24]), .A2(n13324), .ZN(n14549) );
NAND2_X2 U11394 ( .A1(n14550), .A2(n14549), .ZN(n3736) );
NAND2_X2 U11395 ( .A1(H2[23]), .A2(n13324), .ZN(n14552) );
NAND2_X2 U11396 ( .A1(n13348), .A2(SHA1_result[87]), .ZN(n14551) );
NAND3_X2 U11397 ( .A1(n14552), .A2(n13188), .A3(n14551), .ZN(n3737) );
NAND2_X2 U11398 ( .A1(n13197), .A2(SHA1_result[86]), .ZN(n14554) );
NAND2_X2 U11399 ( .A1(H2[22]), .A2(n13323), .ZN(n14553) );
NAND2_X2 U11400 ( .A1(n14554), .A2(n14553), .ZN(n3738) );
NAND2_X2 U11401 ( .A1(H2[21]), .A2(n13323), .ZN(n14556) );
NAND2_X2 U11402 ( .A1(n13348), .A2(SHA1_result[85]), .ZN(n14555) );
NAND3_X2 U11403 ( .A1(n14556), .A2(n13188), .A3(n14555), .ZN(n3739) );
NAND2_X2 U11404 ( .A1(H2[20]), .A2(n13323), .ZN(n14558) );
NAND2_X2 U11405 ( .A1(n13349), .A2(SHA1_result[84]), .ZN(n14557) );
NAND3_X2 U11406 ( .A1(n14558), .A2(n13188), .A3(n14557), .ZN(n3740) );
NAND2_X2 U11407 ( .A1(H2[19]), .A2(n13323), .ZN(n14560) );
NAND2_X2 U11408 ( .A1(n13349), .A2(SHA1_result[83]), .ZN(n14559) );
NAND3_X2 U11409 ( .A1(n14560), .A2(n13188), .A3(n14559), .ZN(n3741) );
NAND2_X2 U11410 ( .A1(n13197), .A2(SHA1_result[82]), .ZN(n14562) );
NAND2_X2 U11411 ( .A1(H2[18]), .A2(n13323), .ZN(n14561) );
NAND2_X2 U11412 ( .A1(n14562), .A2(n14561), .ZN(n3742) );
NAND2_X2 U11413 ( .A1(H2[17]), .A2(n13323), .ZN(n14564) );
NAND2_X2 U11414 ( .A1(n13349), .A2(SHA1_result[81]), .ZN(n14563) );
NAND3_X2 U11415 ( .A1(n14564), .A2(n13188), .A3(n14563), .ZN(n3743) );
NAND2_X2 U11416 ( .A1(n13198), .A2(SHA1_result[80]), .ZN(n14566) );
NAND2_X2 U11417 ( .A1(H2[16]), .A2(n13323), .ZN(n14565) );
NAND2_X2 U11418 ( .A1(n14566), .A2(n14565), .ZN(n3744) );
NAND2_X2 U11419 ( .A1(H2[15]), .A2(n13323), .ZN(n14568) );
NAND2_X2 U11420 ( .A1(n13349), .A2(SHA1_result[79]), .ZN(n14567) );
NAND3_X2 U11421 ( .A1(n14568), .A2(n13188), .A3(n14567), .ZN(n3745) );
NAND2_X2 U11422 ( .A1(H2[14]), .A2(n13323), .ZN(n14570) );
NAND2_X2 U11423 ( .A1(n13349), .A2(SHA1_result[78]), .ZN(n14569) );
NAND3_X2 U11424 ( .A1(n14570), .A2(n13188), .A3(n14569), .ZN(n3746) );
NAND2_X2 U11425 ( .A1(n13198), .A2(SHA1_result[77]), .ZN(n14572) );
NAND2_X2 U11426 ( .A1(H2[13]), .A2(n13323), .ZN(n14571) );
NAND2_X2 U11427 ( .A1(n14572), .A2(n14571), .ZN(n3747) );
NAND2_X2 U11428 ( .A1(H2[12]), .A2(n13323), .ZN(n14574) );
NAND2_X2 U11429 ( .A1(n13349), .A2(SHA1_result[76]), .ZN(n14573) );
NAND3_X2 U11430 ( .A1(n14574), .A2(n13188), .A3(n14573), .ZN(n3748) );
NAND2_X2 U11431 ( .A1(H2[11]), .A2(n13323), .ZN(n14576) );
NAND2_X2 U11432 ( .A1(n13349), .A2(SHA1_result[75]), .ZN(n14575) );
NAND3_X2 U11433 ( .A1(n14576), .A2(n13187), .A3(n14575), .ZN(n3749) );
NAND2_X2 U11434 ( .A1(H2[10]), .A2(n13323), .ZN(n14578) );
NAND2_X2 U11435 ( .A1(n13349), .A2(SHA1_result[74]), .ZN(n14577) );
NAND3_X2 U11436 ( .A1(n14578), .A2(n13187), .A3(n14577), .ZN(n3750) );
NAND2_X2 U11437 ( .A1(n13198), .A2(SHA1_result[73]), .ZN(n14580) );
NAND2_X2 U11438 ( .A1(H2[9]), .A2(n13323), .ZN(n14579) );
NAND2_X2 U11439 ( .A1(n14580), .A2(n14579), .ZN(n3751) );
NAND2_X2 U11440 ( .A1(n13198), .A2(SHA1_result[72]), .ZN(n14582) );
NAND2_X2 U11441 ( .A1(H2[8]), .A2(n13323), .ZN(n14581) );
NAND2_X2 U11442 ( .A1(n14582), .A2(n14581), .ZN(n3752) );
NAND2_X2 U11443 ( .A1(H2[7]), .A2(n13323), .ZN(n14584) );
NAND2_X2 U11444 ( .A1(n13349), .A2(SHA1_result[71]), .ZN(n14583) );
NAND3_X2 U11445 ( .A1(n14584), .A2(n13187), .A3(n14583), .ZN(n3753) );
NAND2_X2 U11446 ( .A1(H2[6]), .A2(n13323), .ZN(n14586) );
NAND2_X2 U11447 ( .A1(n13349), .A2(SHA1_result[70]), .ZN(n14585) );
NAND3_X2 U11448 ( .A1(n14586), .A2(n13187), .A3(n14585), .ZN(n3754) );
NAND2_X2 U11449 ( .A1(H2[5]), .A2(n13323), .ZN(n14588) );
NAND2_X2 U11450 ( .A1(n13349), .A2(SHA1_result[69]), .ZN(n14587) );
NAND3_X2 U11451 ( .A1(n14588), .A2(n13187), .A3(n14587), .ZN(n3755) );
NAND2_X2 U11452 ( .A1(H2[4]), .A2(n13323), .ZN(n14590) );
NAND2_X2 U11453 ( .A1(n13350), .A2(SHA1_result[68]), .ZN(n14589) );
NAND3_X2 U11454 ( .A1(n14590), .A2(n13187), .A3(n14589), .ZN(n3756) );
NAND2_X2 U11455 ( .A1(H2[3]), .A2(n13322), .ZN(n14592) );
NAND2_X2 U11456 ( .A1(n13350), .A2(SHA1_result[67]), .ZN(n14591) );
NAND3_X2 U11457 ( .A1(n14592), .A2(n13187), .A3(n14591), .ZN(n3757) );
NAND2_X2 U11458 ( .A1(H2[2]), .A2(n13322), .ZN(n14594) );
NAND2_X2 U11459 ( .A1(n13350), .A2(SHA1_result[66]), .ZN(n14593) );
NAND3_X2 U11460 ( .A1(n14594), .A2(n13187), .A3(n14593), .ZN(n3758) );
NAND2_X2 U11461 ( .A1(H2[1]), .A2(n13322), .ZN(n14596) );
NAND2_X2 U11462 ( .A1(n13350), .A2(SHA1_result[65]), .ZN(n14595) );
NAND3_X2 U11463 ( .A1(n14596), .A2(n13187), .A3(n14595), .ZN(n3759) );
NAND2_X2 U11464 ( .A1(n13198), .A2(SHA1_result[64]), .ZN(n14598) );
NAND2_X2 U11465 ( .A1(H2[0]), .A2(n13322), .ZN(n14597) );
NAND2_X2 U11466 ( .A1(n14598), .A2(n14597), .ZN(n3760) );
NAND2_X2 U11467 ( .A1(N947), .A2(n13178), .ZN(n14602) );
NAND2_X2 U11468 ( .A1(n13214), .A2(SHA1_result[95]), .ZN(n14600) );
NAND4_X2 U11469 ( .A1(n14602), .A2(n13183), .A3(n14600), .A4(n14599), .ZN(n3889) );
NAND2_X2 U11470 ( .A1(n13198), .A2(SHA1_result[63]), .ZN(n14604) );
NAND2_X2 U11471 ( .A1(H3[31]), .A2(n13322), .ZN(n14603) );
NAND2_X2 U11472 ( .A1(n14604), .A2(n14603), .ZN(n3825) );
NAND2_X2 U11473 ( .A1(n13198), .A2(SHA1_result[62]), .ZN(n14606) );
NAND2_X2 U11474 ( .A1(H3[30]), .A2(n13322), .ZN(n14605) );
NAND2_X2 U11475 ( .A1(n14606), .A2(n14605), .ZN(n3826) );
NAND2_X2 U11476 ( .A1(n13198), .A2(SHA1_result[61]), .ZN(n14608) );
NAND2_X2 U11477 ( .A1(H3[29]), .A2(n13322), .ZN(n14607) );
NAND2_X2 U11478 ( .A1(n14608), .A2(n14607), .ZN(n3827) );
NAND2_X2 U11479 ( .A1(H3[28]), .A2(n13322), .ZN(n14610) );
NAND2_X2 U11480 ( .A1(n13350), .A2(SHA1_result[60]), .ZN(n14609) );
NAND3_X2 U11481 ( .A1(n14610), .A2(n13187), .A3(n14609), .ZN(n3828) );
NAND2_X2 U11482 ( .A1(n13198), .A2(SHA1_result[59]), .ZN(n14612) );
NAND2_X2 U11483 ( .A1(H3[27]), .A2(n13322), .ZN(n14611) );
NAND2_X2 U11484 ( .A1(n14612), .A2(n14611), .ZN(n3829) );
NAND2_X2 U11485 ( .A1(n13198), .A2(SHA1_result[58]), .ZN(n14614) );
NAND2_X2 U11486 ( .A1(H3[26]), .A2(n13322), .ZN(n14613) );
NAND2_X2 U11487 ( .A1(n14614), .A2(n14613), .ZN(n3830) );
NAND2_X2 U11488 ( .A1(n13198), .A2(SHA1_result[57]), .ZN(n14616) );
NAND2_X2 U11489 ( .A1(H3[25]), .A2(n13322), .ZN(n14615) );
NAND2_X2 U11490 ( .A1(n14616), .A2(n14615), .ZN(n3831) );
NAND2_X2 U11491 ( .A1(n13199), .A2(SHA1_result[56]), .ZN(n14618) );
NAND2_X2 U11492 ( .A1(H3[24]), .A2(n13322), .ZN(n14617) );
NAND2_X2 U11493 ( .A1(n14618), .A2(n14617), .ZN(n3832) );
NAND2_X2 U11494 ( .A1(n13199), .A2(SHA1_result[55]), .ZN(n14620) );
NAND2_X2 U11495 ( .A1(H3[23]), .A2(n13322), .ZN(n14619) );
NAND2_X2 U11496 ( .A1(n14620), .A2(n14619), .ZN(n3833) );
NAND2_X2 U11497 ( .A1(n13199), .A2(n14681), .ZN(n14622) );
NAND2_X2 U11498 ( .A1(H3[22]), .A2(n13322), .ZN(n14621) );
NAND2_X2 U11499 ( .A1(n14622), .A2(n14621), .ZN(n3834) );
NAND2_X2 U11500 ( .A1(H3[21]), .A2(n13322), .ZN(n14624) );
NAND2_X2 U11501 ( .A1(n13350), .A2(n14682), .ZN(n14623) );
NAND3_X2 U11502 ( .A1(n14624), .A2(n13186), .A3(n14623), .ZN(n3835) );
NAND2_X2 U11503 ( .A1(H3[20]), .A2(n13322), .ZN(n14626) );
NAND2_X2 U11504 ( .A1(n13350), .A2(n14868), .ZN(n14625) );
NAND3_X2 U11505 ( .A1(n14626), .A2(n13187), .A3(n14625), .ZN(n3836) );
NAND2_X2 U11506 ( .A1(n13199), .A2(SHA1_result[51]), .ZN(n14628) );
NAND2_X2 U11507 ( .A1(H3[19]), .A2(n13322), .ZN(n14627) );
NAND2_X2 U11508 ( .A1(n14628), .A2(n14627), .ZN(n3837) );
NAND2_X2 U11509 ( .A1(n13199), .A2(SHA1_result[50]), .ZN(n14630) );
NAND2_X2 U11510 ( .A1(H3[18]), .A2(n13322), .ZN(n14629) );
NAND2_X2 U11511 ( .A1(n14630), .A2(n14629), .ZN(n3838) );
NAND2_X2 U11512 ( .A1(H3[17]), .A2(n13322), .ZN(n14632) );
NAND2_X2 U11513 ( .A1(n13350), .A2(SHA1_result[49]), .ZN(n14631) );
NAND3_X2 U11514 ( .A1(n14632), .A2(n13186), .A3(n14631), .ZN(n3839) );
NAND2_X2 U11515 ( .A1(n13199), .A2(SHA1_result[48]), .ZN(n14634) );
NAND2_X2 U11516 ( .A1(H3[16]), .A2(n13321), .ZN(n14633) );
NAND2_X2 U11517 ( .A1(n14634), .A2(n14633), .ZN(n3840) );
NAND2_X2 U11518 ( .A1(n13199), .A2(SHA1_result[47]), .ZN(n14636) );
NAND2_X2 U11519 ( .A1(H3[15]), .A2(n13321), .ZN(n14635) );
NAND2_X2 U11520 ( .A1(n14636), .A2(n14635), .ZN(n3841) );
NAND2_X2 U11521 ( .A1(H3[14]), .A2(n13321), .ZN(n14638) );
NAND2_X2 U11522 ( .A1(n13350), .A2(n14830), .ZN(n14637) );
NAND3_X2 U11523 ( .A1(n14638), .A2(n13186), .A3(n14637), .ZN(n3842) );
NAND2_X2 U11524 ( .A1(n13199), .A2(SHA1_result[45]), .ZN(n14640) );
NAND2_X2 U11525 ( .A1(H3[13]), .A2(n13321), .ZN(n14639) );
NAND2_X2 U11526 ( .A1(n14640), .A2(n14639), .ZN(n3843) );
NAND2_X2 U11527 ( .A1(H3[12]), .A2(n13321), .ZN(n14642) );
NAND2_X2 U11528 ( .A1(n13350), .A2(n14817), .ZN(n14641) );
NAND3_X2 U11529 ( .A1(n14642), .A2(n13186), .A3(n14641), .ZN(n3844) );
NAND2_X2 U11530 ( .A1(n13199), .A2(n14810), .ZN(n14644) );
NAND2_X2 U11531 ( .A1(H3[11]), .A2(n13321), .ZN(n14643) );
NAND2_X2 U11532 ( .A1(n14644), .A2(n14643), .ZN(n3845) );
NAND2_X2 U11533 ( .A1(H3[10]), .A2(n13321), .ZN(n14646) );
NAND2_X2 U11534 ( .A1(n13350), .A2(SHA1_result[42]), .ZN(n14645) );
NAND3_X2 U11535 ( .A1(n14646), .A2(n13186), .A3(n14645), .ZN(n3846) );
NAND2_X2 U11536 ( .A1(n13199), .A2(n14797), .ZN(n14648) );
NAND2_X2 U11537 ( .A1(H3[9]), .A2(n13321), .ZN(n14647) );
NAND2_X2 U11538 ( .A1(n14648), .A2(n14647), .ZN(n3847) );
NAND2_X2 U11539 ( .A1(n13199), .A2(SHA1_result[40]), .ZN(n14650) );
NAND2_X2 U11540 ( .A1(H3[8]), .A2(n13321), .ZN(n14649) );
NAND2_X2 U11541 ( .A1(n14650), .A2(n14649), .ZN(n3848) );
NAND2_X2 U11542 ( .A1(n13195), .A2(SHA1_result[39]), .ZN(n14652) );
NAND2_X2 U11543 ( .A1(H3[7]), .A2(n13321), .ZN(n14651) );
NAND2_X2 U11544 ( .A1(n14652), .A2(n14651), .ZN(n3849) );
NAND2_X2 U11545 ( .A1(H3[6]), .A2(n13321), .ZN(n14654) );
NAND2_X2 U11546 ( .A1(n13351), .A2(n14778), .ZN(n14653) );
NAND3_X2 U11547 ( .A1(n14654), .A2(n13186), .A3(n14653), .ZN(n3850) );
NAND2_X2 U11548 ( .A1(H3[5]), .A2(n13321), .ZN(n14656) );
NAND2_X2 U11549 ( .A1(n13351), .A2(n14770), .ZN(n14655) );
NAND3_X2 U11550 ( .A1(n14656), .A2(n13186), .A3(n14655), .ZN(n3851) );
NAND2_X2 U11551 ( .A1(H3[4]), .A2(n13321), .ZN(n14658) );
NAND2_X2 U11552 ( .A1(n13351), .A2(SHA1_result[36]), .ZN(n14657) );
NAND3_X2 U11553 ( .A1(n14658), .A2(n13186), .A3(n14657), .ZN(n3852) );
NAND2_X2 U11554 ( .A1(n13194), .A2(SHA1_result[35]), .ZN(n14660) );
NAND2_X2 U11555 ( .A1(H3[3]), .A2(n13321), .ZN(n14659) );
NAND2_X2 U11556 ( .A1(n14660), .A2(n14659), .ZN(n3853) );
NAND2_X2 U11557 ( .A1(H3[2]), .A2(n13321), .ZN(n14662) );
NAND2_X2 U11558 ( .A1(n13351), .A2(SHA1_result[34]), .ZN(n14661) );
NAND3_X2 U11559 ( .A1(n14662), .A2(n13186), .A3(n14661), .ZN(n3854) );
NAND2_X2 U11560 ( .A1(H3[1]), .A2(n13321), .ZN(n14664) );
NAND2_X2 U11561 ( .A1(n13351), .A2(n14742), .ZN(n14663) );
NAND3_X2 U11562 ( .A1(n14664), .A2(n13189), .A3(n14663), .ZN(n3855) );
NAND2_X2 U11563 ( .A1(n13193), .A2(SHA1_result[32]), .ZN(n14666) );
NAND2_X2 U11564 ( .A1(H3[0]), .A2(n13321), .ZN(n14665) );
NAND2_X2 U11565 ( .A1(n14666), .A2(n14665), .ZN(n3856) );
NAND2_X2 U11566 ( .A1(n13205), .A2(SHA1_result[95]), .ZN(n14669) );
NAND2_X2 U11567 ( .A1(N979), .A2(n13209), .ZN(n14668) );
NAND2_X2 U11568 ( .A1(n13215), .A2(SHA1_result[63]), .ZN(n14667) );
NAND3_X2 U11569 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(n3857) );
NAND2_X2 U11570 ( .A1(n13332), .A2(SHA1_result[63]), .ZN(n12069) );
NAND2_X2 U11571 ( .A1(n13335), .A2(SHA1_result[31]), .ZN(n12070) );
NAND2_X2 U11572 ( .A1(n13336), .A2(SHA1_result[95]), .ZN(n12071) );
NOR2_X2 U11573 ( .A1(n13342), .A2(n12913), .ZN(n14671) );
NOR2_X2 U11574 ( .A1(n13341), .A2(n13002), .ZN(n14670) );
NOR3_X2 U11575 ( .A1(n12075), .A2(n14671), .A3(n14670), .ZN(n12072) );
NAND2_X2 U11576 ( .A1(n13332), .A2(SHA1_result[62]), .ZN(n12062) );
NAND2_X2 U11577 ( .A1(n13335), .A2(SHA1_result[30]), .ZN(n12063) );
NAND2_X2 U11578 ( .A1(n13336), .A2(SHA1_result[94]), .ZN(n12064) );
NOR2_X2 U11579 ( .A1(n13342), .A2(n12911), .ZN(n14673) );
NOR2_X2 U11580 ( .A1(n13341), .A2(n13007), .ZN(n14672) );
NOR3_X2 U11581 ( .A1(n12068), .A2(n14673), .A3(n14672), .ZN(n12065) );
NAND2_X2 U11582 ( .A1(n13332), .A2(SHA1_result[61]), .ZN(n12055) );
NAND2_X2 U11583 ( .A1(n13335), .A2(SHA1_result[29]), .ZN(n12056) );
NAND2_X2 U11584 ( .A1(n13336), .A2(SHA1_result[93]), .ZN(n12057) );
NOR2_X2 U11585 ( .A1(n13342), .A2(n12909), .ZN(n14675) );
NOR2_X2 U11586 ( .A1(n13341), .A2(n13013), .ZN(n14674) );
NOR3_X2 U11587 ( .A1(n12061), .A2(n14675), .A3(n14674), .ZN(n12058) );
NAND2_X2 U11588 ( .A1(n13332), .A2(SHA1_result[60]), .ZN(n12048) );
NAND2_X2 U11589 ( .A1(n13335), .A2(SHA1_result[28]), .ZN(n12049) );
NAND2_X2 U11590 ( .A1(n13336), .A2(SHA1_result[92]), .ZN(n12050) );
NOR2_X2 U11591 ( .A1(n13342), .A2(n12907), .ZN(n14677) );
NOR2_X2 U11592 ( .A1(n13341), .A2(n13014), .ZN(n14676) );
NOR3_X2 U11593 ( .A1(n12054), .A2(n14677), .A3(n14676), .ZN(n12051) );
NAND2_X2 U11594 ( .A1(n13332), .A2(SHA1_result[59]), .ZN(n12041) );
NAND2_X2 U11595 ( .A1(n13335), .A2(SHA1_result[27]), .ZN(n12042) );
NAND2_X2 U11596 ( .A1(n13336), .A2(SHA1_result[91]), .ZN(n12043) );
NOR2_X2 U11597 ( .A1(n13342), .A2(n12905), .ZN(n14679) );
NOR2_X2 U11598 ( .A1(n13341), .A2(n13008), .ZN(n14678) );
NOR3_X2 U11599 ( .A1(n12047), .A2(n14679), .A3(n14678), .ZN(n12044) );
NOR2_X2 U11600 ( .A1(n13341), .A2(n13003), .ZN(n12038) );
NOR2_X2 U11601 ( .A1(n13342), .A2(n12903), .ZN(n12039) );
NAND2_X2 U11602 ( .A1(n13332), .A2(SHA1_result[58]), .ZN(n12034) );
NAND2_X2 U11603 ( .A1(n13335), .A2(SHA1_result[26]), .ZN(n12035) );
NAND2_X2 U11604 ( .A1(n13336), .A2(SHA1_result[90]), .ZN(n12036) );
NOR2_X2 U11605 ( .A1(n13341), .A2(n13009), .ZN(n12031) );
NOR2_X2 U11606 ( .A1(n13342), .A2(n12901), .ZN(n12032) );
NAND2_X2 U11607 ( .A1(n13332), .A2(SHA1_result[57]), .ZN(n12027) );
NAND2_X2 U11608 ( .A1(n13335), .A2(SHA1_result[25]), .ZN(n12028) );
NAND2_X2 U11609 ( .A1(n13336), .A2(SHA1_result[89]), .ZN(n12029) );
NOR2_X2 U11610 ( .A1(n13341), .A2(n13010), .ZN(n12024) );
NOR2_X2 U11611 ( .A1(n13342), .A2(n12899), .ZN(n12025) );
NAND2_X2 U11612 ( .A1(n13332), .A2(SHA1_result[56]), .ZN(n12020) );
NAND2_X2 U11613 ( .A1(n13335), .A2(SHA1_result[24]), .ZN(n12021) );
NAND2_X2 U11614 ( .A1(n13336), .A2(SHA1_result[88]), .ZN(n12022) );
NOR2_X2 U11615 ( .A1(n13341), .A2(n14680), .ZN(n12017) );
NOR2_X2 U11616 ( .A1(n13342), .A2(n12897), .ZN(n12018) );
NAND2_X2 U11617 ( .A1(n13332), .A2(SHA1_result[55]), .ZN(n12013) );
NAND2_X2 U11618 ( .A1(n13335), .A2(SHA1_result[23]), .ZN(n12014) );
NAND2_X2 U11619 ( .A1(n13336), .A2(SHA1_result[87]), .ZN(n12015) );
NOR2_X2 U11620 ( .A1(n13341), .A2(n13006), .ZN(n12010) );
NOR2_X2 U11621 ( .A1(n13342), .A2(n12895), .ZN(n12011) );
NAND2_X2 U11622 ( .A1(n13332), .A2(n14681), .ZN(n12006) );
NAND2_X2 U11623 ( .A1(n13335), .A2(SHA1_result[22]), .ZN(n12007) );
NAND2_X2 U11624 ( .A1(n13336), .A2(SHA1_result[86]), .ZN(n12008) );
NAND2_X2 U11625 ( .A1(n13331), .A2(n14682), .ZN(n11999) );
NAND2_X2 U11626 ( .A1(n13334), .A2(SHA1_result[21]), .ZN(n12000) );
NAND2_X2 U11627 ( .A1(n13336), .A2(SHA1_result[85]), .ZN(n12001) );
NOR2_X2 U11628 ( .A1(n13342), .A2(n12893), .ZN(n14684) );
NOR2_X2 U11629 ( .A1(n13340), .A2(n13011), .ZN(n14683) );
NOR3_X2 U11630 ( .A1(n12005), .A2(n14684), .A3(n14683), .ZN(n12002) );
NAND2_X2 U11631 ( .A1(n14956), .A2(n15425), .ZN(n11845) );
NAND2_X2 U11632 ( .A1(n14954), .A2(read_counter[2]), .ZN(n11844) );
NAND2_X2 U11633 ( .A1(n14956), .A2(read_counter[0]), .ZN(n14685) );
NAND2_X2 U11634 ( .A1(n11837), .A2(n14685), .ZN(n14686) );
NAND2_X2 U11635 ( .A1(read_counter[1]), .A2(n14686), .ZN(n11838) );
NAND3_X2 U11636 ( .A1(n11837), .A2(n14956), .A3(n14952), .ZN(n11836) );
NAND2_X2 U11637 ( .A1(n14687), .A2(n14953), .ZN(n14731) );
NAND2_X2 U11638 ( .A1(n14724), .A2(n14689), .ZN(n14690) );
NAND2_X2 U11639 ( .A1(n15419), .A2(n13271), .ZN(n11006) );
NAND2_X2 U11640 ( .A1(n15404), .A2(n13271), .ZN(n11003) );
NAND2_X2 U11641 ( .A1(n15389), .A2(n13271), .ZN(n11000) );
NAND2_X2 U11642 ( .A1(n15374), .A2(n13271), .ZN(n10997) );
NAND2_X2 U11643 ( .A1(n15359), .A2(n13271), .ZN(n10994) );
NAND2_X2 U11644 ( .A1(n15344), .A2(n13271), .ZN(n10991) );
NAND2_X2 U11645 ( .A1(n15329), .A2(n13271), .ZN(n10988) );
NAND2_X2 U11646 ( .A1(n15314), .A2(n13271), .ZN(n10985) );
NAND2_X2 U11647 ( .A1(n15299), .A2(n13271), .ZN(n10982) );
NAND2_X2 U11648 ( .A1(n15284), .A2(n13271), .ZN(n10979) );
NAND2_X2 U11649 ( .A1(n15269), .A2(n13271), .ZN(n10976) );
NAND2_X2 U11650 ( .A1(n15254), .A2(n13271), .ZN(n10973) );
NAND2_X2 U11651 ( .A1(n15239), .A2(n13271), .ZN(n10970) );
NAND2_X2 U11652 ( .A1(n15224), .A2(n13271), .ZN(n10967) );
NAND2_X2 U11653 ( .A1(n15209), .A2(n13270), .ZN(n10964) );
NAND2_X2 U11654 ( .A1(n15195), .A2(n13270), .ZN(n10961) );
NAND2_X2 U11655 ( .A1(n15181), .A2(n13270), .ZN(n10958) );
NAND2_X2 U11656 ( .A1(n15167), .A2(n13270), .ZN(n10955) );
NAND2_X2 U11657 ( .A1(n15153), .A2(n13270), .ZN(n10952) );
NAND2_X2 U11658 ( .A1(n15139), .A2(n13270), .ZN(n10949) );
NAND2_X2 U11659 ( .A1(n15125), .A2(n13270), .ZN(n10946) );
NAND2_X2 U11660 ( .A1(n15111), .A2(n13270), .ZN(n10943) );
NAND2_X2 U11661 ( .A1(n15097), .A2(n13270), .ZN(n10940) );
NAND2_X2 U11662 ( .A1(n15083), .A2(n13270), .ZN(n10937) );
NAND2_X2 U11663 ( .A1(n15069), .A2(n13270), .ZN(n10934) );
NAND2_X2 U11664 ( .A1(n15055), .A2(n13270), .ZN(n10931) );
NAND2_X2 U11665 ( .A1(n15041), .A2(n13270), .ZN(n10928) );
NAND2_X2 U11666 ( .A1(n15027), .A2(n13270), .ZN(n10925) );
NAND2_X2 U11667 ( .A1(n15013), .A2(n13270), .ZN(n10922) );
NAND2_X2 U11668 ( .A1(n14999), .A2(n13270), .ZN(n10919) );
NAND2_X2 U11669 ( .A1(n14985), .A2(n13270), .ZN(n10916) );
NAND2_X2 U11670 ( .A1(n14971), .A2(n13270), .ZN(n10911) );
NAND2_X2 U11671 ( .A1(n13024), .A2(n14722), .ZN(n14692) );
NAND2_X2 U11672 ( .A1(n14724), .A2(n14693), .ZN(n14695) );
NAND2_X2 U11673 ( .A1(n14724), .A2(n14694), .ZN(n14700) );
NAND2_X2 U11674 ( .A1(n15418), .A2(n13225), .ZN(n10906) );
NAND2_X2 U11675 ( .A1(n15403), .A2(n13225), .ZN(n10903) );
NAND2_X2 U11676 ( .A1(n15388), .A2(n13225), .ZN(n10900) );
NAND2_X2 U11677 ( .A1(n15373), .A2(n13225), .ZN(n10897) );
NAND2_X2 U11678 ( .A1(n15358), .A2(n13225), .ZN(n10894) );
NAND2_X2 U11679 ( .A1(n15343), .A2(n13225), .ZN(n10891) );
NAND2_X2 U11680 ( .A1(n15328), .A2(n13225), .ZN(n10888) );
NAND2_X2 U11681 ( .A1(n15313), .A2(n13225), .ZN(n10885) );
NAND2_X2 U11682 ( .A1(n15298), .A2(n13225), .ZN(n10882) );
NAND2_X2 U11683 ( .A1(n15283), .A2(n13225), .ZN(n10879) );
NAND2_X2 U11684 ( .A1(n15268), .A2(n13225), .ZN(n10876) );
NAND2_X2 U11685 ( .A1(n15253), .A2(n13226), .ZN(n10873) );
NAND2_X2 U11686 ( .A1(n15238), .A2(n13226), .ZN(n10870) );
NAND2_X2 U11687 ( .A1(n15223), .A2(n13226), .ZN(n10867) );
NAND2_X2 U11688 ( .A1(n15208), .A2(n13226), .ZN(n10864) );
NAND2_X2 U11689 ( .A1(n15194), .A2(n13226), .ZN(n10861) );
NAND2_X2 U11690 ( .A1(n15180), .A2(n13226), .ZN(n10858) );
NAND2_X2 U11691 ( .A1(n15166), .A2(n13226), .ZN(n10855) );
NAND2_X2 U11692 ( .A1(n15152), .A2(n13226), .ZN(n10852) );
NAND2_X2 U11693 ( .A1(n15138), .A2(n13226), .ZN(n10849) );
NAND2_X2 U11694 ( .A1(n15124), .A2(n13226), .ZN(n10846) );
NAND2_X2 U11695 ( .A1(n15110), .A2(n13226), .ZN(n10843) );
NAND2_X2 U11696 ( .A1(n15096), .A2(n13227), .ZN(n10840) );
NAND2_X2 U11697 ( .A1(n15082), .A2(n13227), .ZN(n10837) );
NAND2_X2 U11698 ( .A1(n15068), .A2(n13227), .ZN(n10834) );
NAND2_X2 U11699 ( .A1(n15054), .A2(n13227), .ZN(n10831) );
NAND2_X2 U11700 ( .A1(n15040), .A2(n13227), .ZN(n10828) );
NAND2_X2 U11701 ( .A1(n15026), .A2(n13227), .ZN(n10825) );
NAND2_X2 U11702 ( .A1(n15012), .A2(n13227), .ZN(n10822) );
NAND2_X2 U11703 ( .A1(n14998), .A2(n13227), .ZN(n10819) );
NAND2_X2 U11704 ( .A1(n14984), .A2(n13227), .ZN(n10816) );
NAND2_X2 U11705 ( .A1(n14970), .A2(n13227), .ZN(n10811) );
INV_X4 U11706 ( .A(n14729), .ZN(n14727) );
NAND2_X2 U11707 ( .A1(n13024), .A2(n14727), .ZN(n14696) );
NAND2_X2 U11708 ( .A1(n14724), .A2(n14729), .ZN(n14697) );
NAND2_X2 U11709 ( .A1(n15417), .A2(n13228), .ZN(n10807) );
NAND2_X2 U11710 ( .A1(n15402), .A2(n13228), .ZN(n10804) );
NAND2_X2 U11711 ( .A1(n15387), .A2(n13228), .ZN(n10801) );
NAND2_X2 U11712 ( .A1(n15372), .A2(n13228), .ZN(n10798) );
NAND2_X2 U11713 ( .A1(n15357), .A2(n13228), .ZN(n10795) );
NAND2_X2 U11714 ( .A1(n15342), .A2(n13228), .ZN(n10792) );
NAND2_X2 U11715 ( .A1(n15327), .A2(n13228), .ZN(n10789) );
NAND2_X2 U11716 ( .A1(n15312), .A2(n13228), .ZN(n10786) );
NAND2_X2 U11717 ( .A1(n15297), .A2(n13228), .ZN(n10783) );
NAND2_X2 U11718 ( .A1(n15282), .A2(n13228), .ZN(n10780) );
NAND2_X2 U11719 ( .A1(n15267), .A2(n13228), .ZN(n10777) );
NAND2_X2 U11720 ( .A1(n15252), .A2(n13229), .ZN(n10774) );
NAND2_X2 U11721 ( .A1(n15237), .A2(n13229), .ZN(n10771) );
NAND2_X2 U11722 ( .A1(n15222), .A2(n13229), .ZN(n10768) );
NAND2_X2 U11723 ( .A1(n15207), .A2(n13229), .ZN(n10765) );
NAND2_X2 U11724 ( .A1(n15193), .A2(n13229), .ZN(n10762) );
NAND2_X2 U11725 ( .A1(n15179), .A2(n13229), .ZN(n10759) );
NAND2_X2 U11726 ( .A1(n15165), .A2(n13229), .ZN(n10756) );
NAND2_X2 U11727 ( .A1(n15151), .A2(n13229), .ZN(n10753) );
NAND2_X2 U11728 ( .A1(n15137), .A2(n13229), .ZN(n10750) );
NAND2_X2 U11729 ( .A1(n15123), .A2(n13229), .ZN(n10747) );
NAND2_X2 U11730 ( .A1(n15109), .A2(n13229), .ZN(n10744) );
NAND2_X2 U11731 ( .A1(n15095), .A2(n13230), .ZN(n10741) );
NAND2_X2 U11732 ( .A1(n15081), .A2(n13230), .ZN(n10738) );
NAND2_X2 U11733 ( .A1(n15067), .A2(n13230), .ZN(n10735) );
NAND2_X2 U11734 ( .A1(n15053), .A2(n13230), .ZN(n10732) );
NAND2_X2 U11735 ( .A1(n15039), .A2(n13230), .ZN(n10729) );
NAND2_X2 U11736 ( .A1(n15025), .A2(n13230), .ZN(n10726) );
NAND2_X2 U11737 ( .A1(n15011), .A2(n13230), .ZN(n10723) );
NAND2_X2 U11738 ( .A1(n14997), .A2(n13230), .ZN(n10720) );
NAND2_X2 U11739 ( .A1(n14983), .A2(n13230), .ZN(n10717) );
NAND2_X2 U11740 ( .A1(n14969), .A2(n13230), .ZN(n10712) );
INV_X4 U11741 ( .A(n14699), .ZN(n14704) );
NAND2_X2 U11742 ( .A1(n13024), .A2(n14704), .ZN(n14698) );
NAND2_X2 U11743 ( .A1(n14724), .A2(n14699), .ZN(n14715) );
NAND2_X2 U11744 ( .A1(n15416), .A2(n13231), .ZN(n10706) );
NAND2_X2 U11745 ( .A1(n15401), .A2(n13231), .ZN(n10703) );
NAND2_X2 U11746 ( .A1(n15386), .A2(n13231), .ZN(n10700) );
NAND2_X2 U11747 ( .A1(n15371), .A2(n13231), .ZN(n10697) );
NAND2_X2 U11748 ( .A1(n15356), .A2(n13231), .ZN(n10694) );
NAND2_X2 U11749 ( .A1(n15341), .A2(n13231), .ZN(n10691) );
NAND2_X2 U11750 ( .A1(n15326), .A2(n13231), .ZN(n10688) );
NAND2_X2 U11751 ( .A1(n15311), .A2(n13231), .ZN(n10685) );
NAND2_X2 U11752 ( .A1(n15296), .A2(n13231), .ZN(n10682) );
NAND2_X2 U11753 ( .A1(n15281), .A2(n13231), .ZN(n10679) );
NAND2_X2 U11754 ( .A1(n15266), .A2(n13231), .ZN(n10676) );
NAND2_X2 U11755 ( .A1(n15251), .A2(n13232), .ZN(n10673) );
NAND2_X2 U11756 ( .A1(n15236), .A2(n13232), .ZN(n10670) );
NAND2_X2 U11757 ( .A1(n15221), .A2(n13232), .ZN(n10667) );
NAND2_X2 U11758 ( .A1(n15206), .A2(n13232), .ZN(n10664) );
NAND2_X2 U11759 ( .A1(n15192), .A2(n13232), .ZN(n10661) );
NAND2_X2 U11760 ( .A1(n15178), .A2(n13232), .ZN(n10658) );
NAND2_X2 U11761 ( .A1(n15164), .A2(n13232), .ZN(n10655) );
NAND2_X2 U11762 ( .A1(n15150), .A2(n13232), .ZN(n10652) );
NAND2_X2 U11763 ( .A1(n15136), .A2(n13232), .ZN(n10649) );
NAND2_X2 U11764 ( .A1(n15122), .A2(n13232), .ZN(n10646) );
NAND2_X2 U11765 ( .A1(n15108), .A2(n13232), .ZN(n10643) );
NAND2_X2 U11766 ( .A1(n15094), .A2(n13233), .ZN(n10640) );
NAND2_X2 U11767 ( .A1(n15080), .A2(n13233), .ZN(n10637) );
NAND2_X2 U11768 ( .A1(n15066), .A2(n13233), .ZN(n10634) );
NAND2_X2 U11769 ( .A1(n15052), .A2(n13233), .ZN(n10631) );
NAND2_X2 U11770 ( .A1(n15038), .A2(n13233), .ZN(n10628) );
NAND2_X2 U11771 ( .A1(n15024), .A2(n13233), .ZN(n10625) );
NAND2_X2 U11772 ( .A1(n15010), .A2(n13233), .ZN(n10622) );
NAND2_X2 U11773 ( .A1(n14996), .A2(n13233), .ZN(n10619) );
NAND2_X2 U11774 ( .A1(n14982), .A2(n13233), .ZN(n10616) );
NAND2_X2 U11775 ( .A1(n14968), .A2(n13233), .ZN(n10611) );
NAND2_X2 U11776 ( .A1(n14724), .A2(n10609), .ZN(n14701) );
NAND2_X2 U11777 ( .A1(n15415), .A2(n13236), .ZN(n10607) );
NAND2_X2 U11778 ( .A1(n15400), .A2(n13236), .ZN(n10604) );
NAND2_X2 U11779 ( .A1(n15385), .A2(n13236), .ZN(n10601) );
NAND2_X2 U11780 ( .A1(n15370), .A2(n13236), .ZN(n10598) );
NAND2_X2 U11781 ( .A1(n15355), .A2(n13236), .ZN(n10595) );
NAND2_X2 U11782 ( .A1(n15340), .A2(n13236), .ZN(n10592) );
NAND2_X2 U11783 ( .A1(n15325), .A2(n13236), .ZN(n10589) );
NAND2_X2 U11784 ( .A1(n15310), .A2(n13236), .ZN(n10586) );
NAND2_X2 U11785 ( .A1(n15295), .A2(n13236), .ZN(n10583) );
NAND2_X2 U11786 ( .A1(n15280), .A2(n13236), .ZN(n10580) );
NAND2_X2 U11787 ( .A1(n15265), .A2(n13235), .ZN(n10577) );
NAND2_X2 U11788 ( .A1(n15250), .A2(n13235), .ZN(n10574) );
NAND2_X2 U11789 ( .A1(n15235), .A2(n13235), .ZN(n10571) );
NAND2_X2 U11790 ( .A1(n15220), .A2(n13235), .ZN(n10568) );
NAND2_X2 U11791 ( .A1(n15205), .A2(n13235), .ZN(n10565) );
NAND2_X2 U11792 ( .A1(n15191), .A2(n13235), .ZN(n10562) );
NAND2_X2 U11793 ( .A1(n15177), .A2(n13235), .ZN(n10559) );
NAND2_X2 U11794 ( .A1(n15163), .A2(n13235), .ZN(n10556) );
NAND2_X2 U11795 ( .A1(n15149), .A2(n13235), .ZN(n10553) );
NAND2_X2 U11796 ( .A1(n15135), .A2(n13235), .ZN(n10550) );
NAND2_X2 U11797 ( .A1(n15121), .A2(n13235), .ZN(n10547) );
NAND2_X2 U11798 ( .A1(n15107), .A2(n13234), .ZN(n10544) );
NAND2_X2 U11799 ( .A1(n15093), .A2(n13234), .ZN(n10541) );
NAND2_X2 U11800 ( .A1(n15079), .A2(n13234), .ZN(n10538) );
NAND2_X2 U11801 ( .A1(n15065), .A2(n13234), .ZN(n10535) );
NAND2_X2 U11802 ( .A1(n15051), .A2(n13234), .ZN(n10532) );
NAND2_X2 U11803 ( .A1(n15037), .A2(n13234), .ZN(n10529) );
NAND2_X2 U11804 ( .A1(n15023), .A2(n13234), .ZN(n10526) );
NAND2_X2 U11805 ( .A1(n15009), .A2(n13234), .ZN(n10523) );
NAND2_X2 U11806 ( .A1(n14995), .A2(n13234), .ZN(n10520) );
NAND2_X2 U11807 ( .A1(n14981), .A2(n13234), .ZN(n10517) );
NAND2_X2 U11808 ( .A1(n14967), .A2(n13234), .ZN(n10512) );
NAND2_X2 U11809 ( .A1(n14722), .A2(n14705), .ZN(n10510) );
NAND2_X2 U11810 ( .A1(n14724), .A2(n10510), .ZN(n14702) );
NAND2_X2 U11811 ( .A1(n15414), .A2(n13239), .ZN(n10508) );
NAND2_X2 U11812 ( .A1(n15399), .A2(n13239), .ZN(n10505) );
NAND2_X2 U11813 ( .A1(n15384), .A2(n13239), .ZN(n10502) );
NAND2_X2 U11814 ( .A1(n15369), .A2(n13239), .ZN(n10499) );
NAND2_X2 U11815 ( .A1(n15354), .A2(n13239), .ZN(n10496) );
NAND2_X2 U11816 ( .A1(n15339), .A2(n13239), .ZN(n10493) );
NAND2_X2 U11817 ( .A1(n15324), .A2(n13239), .ZN(n10490) );
NAND2_X2 U11818 ( .A1(n15309), .A2(n13239), .ZN(n10487) );
NAND2_X2 U11819 ( .A1(n15294), .A2(n13239), .ZN(n10484) );
NAND2_X2 U11820 ( .A1(n15279), .A2(n13239), .ZN(n10481) );
NAND2_X2 U11821 ( .A1(n15264), .A2(n13238), .ZN(n10478) );
NAND2_X2 U11822 ( .A1(n15249), .A2(n13238), .ZN(n10475) );
NAND2_X2 U11823 ( .A1(n15234), .A2(n13238), .ZN(n10472) );
NAND2_X2 U11824 ( .A1(n15219), .A2(n13238), .ZN(n10469) );
NAND2_X2 U11825 ( .A1(n15204), .A2(n13238), .ZN(n10466) );
NAND2_X2 U11826 ( .A1(n15190), .A2(n13238), .ZN(n10463) );
NAND2_X2 U11827 ( .A1(n15176), .A2(n13238), .ZN(n10460) );
NAND2_X2 U11828 ( .A1(n15162), .A2(n13238), .ZN(n10457) );
NAND2_X2 U11829 ( .A1(n15148), .A2(n13238), .ZN(n10454) );
NAND2_X2 U11830 ( .A1(n15134), .A2(n13238), .ZN(n10451) );
NAND2_X2 U11831 ( .A1(n15120), .A2(n13238), .ZN(n10448) );
NAND2_X2 U11832 ( .A1(n15106), .A2(n13237), .ZN(n10445) );
NAND2_X2 U11833 ( .A1(n15092), .A2(n13237), .ZN(n10442) );
NAND2_X2 U11834 ( .A1(n15078), .A2(n13237), .ZN(n10439) );
NAND2_X2 U11835 ( .A1(n15064), .A2(n13237), .ZN(n10436) );
NAND2_X2 U11836 ( .A1(n15050), .A2(n13237), .ZN(n10433) );
NAND2_X2 U11837 ( .A1(n15036), .A2(n13237), .ZN(n10430) );
NAND2_X2 U11838 ( .A1(n15022), .A2(n13237), .ZN(n10427) );
NAND2_X2 U11839 ( .A1(n15008), .A2(n13237), .ZN(n10424) );
NAND2_X2 U11840 ( .A1(n14994), .A2(n13237), .ZN(n10421) );
NAND2_X2 U11841 ( .A1(n14980), .A2(n13237), .ZN(n10418) );
NAND2_X2 U11842 ( .A1(n14966), .A2(n13237), .ZN(n10413) );
NAND2_X2 U11843 ( .A1(n14705), .A2(n14727), .ZN(n10411) );
NAND2_X2 U11844 ( .A1(n14724), .A2(n10411), .ZN(n14703) );
NAND2_X2 U11845 ( .A1(n15413), .A2(n13242), .ZN(n10409) );
NAND2_X2 U11846 ( .A1(n15398), .A2(n13242), .ZN(n10406) );
NAND2_X2 U11847 ( .A1(n15383), .A2(n13242), .ZN(n10403) );
NAND2_X2 U11848 ( .A1(n15368), .A2(n13242), .ZN(n10400) );
NAND2_X2 U11849 ( .A1(n15353), .A2(n13242), .ZN(n10397) );
NAND2_X2 U11850 ( .A1(n15338), .A2(n13242), .ZN(n10394) );
NAND2_X2 U11851 ( .A1(n15323), .A2(n13242), .ZN(n10391) );
NAND2_X2 U11852 ( .A1(n15308), .A2(n13242), .ZN(n10388) );
NAND2_X2 U11853 ( .A1(n15293), .A2(n13242), .ZN(n10385) );
NAND2_X2 U11854 ( .A1(n15278), .A2(n13242), .ZN(n10382) );
NAND2_X2 U11855 ( .A1(n15263), .A2(n13241), .ZN(n10379) );
NAND2_X2 U11856 ( .A1(n15248), .A2(n13241), .ZN(n10376) );
NAND2_X2 U11857 ( .A1(n15233), .A2(n13241), .ZN(n10373) );
NAND2_X2 U11858 ( .A1(n15218), .A2(n13241), .ZN(n10370) );
NAND2_X2 U11859 ( .A1(n15203), .A2(n13241), .ZN(n10367) );
NAND2_X2 U11860 ( .A1(n15189), .A2(n13241), .ZN(n10364) );
NAND2_X2 U11861 ( .A1(n15175), .A2(n13241), .ZN(n10361) );
NAND2_X2 U11862 ( .A1(n15161), .A2(n13241), .ZN(n10358) );
NAND2_X2 U11863 ( .A1(n15147), .A2(n13241), .ZN(n10355) );
NAND2_X2 U11864 ( .A1(n15133), .A2(n13241), .ZN(n10352) );
NAND2_X2 U11865 ( .A1(n15119), .A2(n13241), .ZN(n10349) );
NAND2_X2 U11866 ( .A1(n15105), .A2(n13240), .ZN(n10346) );
NAND2_X2 U11867 ( .A1(n15091), .A2(n13240), .ZN(n10343) );
NAND2_X2 U11868 ( .A1(n15077), .A2(n13240), .ZN(n10340) );
NAND2_X2 U11869 ( .A1(n15063), .A2(n13240), .ZN(n10337) );
NAND2_X2 U11870 ( .A1(n15049), .A2(n13240), .ZN(n10334) );
NAND2_X2 U11871 ( .A1(n15035), .A2(n13240), .ZN(n10331) );
NAND2_X2 U11872 ( .A1(n15021), .A2(n13240), .ZN(n10328) );
NAND2_X2 U11873 ( .A1(n15007), .A2(n13240), .ZN(n10325) );
NAND2_X2 U11874 ( .A1(n14993), .A2(n13240), .ZN(n10322) );
NAND2_X2 U11875 ( .A1(n14979), .A2(n13240), .ZN(n10319) );
NAND2_X2 U11876 ( .A1(n14965), .A2(n13240), .ZN(n10314) );
NAND2_X2 U11877 ( .A1(n13028), .A2(n14705), .ZN(n14706) );
NAND2_X2 U11878 ( .A1(n14724), .A2(n14707), .ZN(n14708) );
NAND2_X2 U11879 ( .A1(n15412), .A2(n13243), .ZN(n10309) );
NAND2_X2 U11880 ( .A1(n15397), .A2(n13243), .ZN(n10306) );
NAND2_X2 U11881 ( .A1(n15382), .A2(n13243), .ZN(n10303) );
NAND2_X2 U11882 ( .A1(n15367), .A2(n13243), .ZN(n10300) );
NAND2_X2 U11883 ( .A1(n15352), .A2(n13243), .ZN(n10297) );
NAND2_X2 U11884 ( .A1(n15337), .A2(n13243), .ZN(n10294) );
NAND2_X2 U11885 ( .A1(n15322), .A2(n13243), .ZN(n10291) );
NAND2_X2 U11886 ( .A1(n15307), .A2(n13243), .ZN(n10288) );
NAND2_X2 U11887 ( .A1(n15292), .A2(n13243), .ZN(n10285) );
NAND2_X2 U11888 ( .A1(n15277), .A2(n13243), .ZN(n10282) );
NAND2_X2 U11889 ( .A1(n15262), .A2(n13243), .ZN(n10279) );
NAND2_X2 U11890 ( .A1(n15247), .A2(n13244), .ZN(n10276) );
NAND2_X2 U11891 ( .A1(n15232), .A2(n13244), .ZN(n10273) );
NAND2_X2 U11892 ( .A1(n15217), .A2(n13244), .ZN(n10270) );
NAND2_X2 U11893 ( .A1(n15202), .A2(n13244), .ZN(n10267) );
NAND2_X2 U11894 ( .A1(n15188), .A2(n13244), .ZN(n10264) );
NAND2_X2 U11895 ( .A1(n15174), .A2(n13244), .ZN(n10261) );
NAND2_X2 U11896 ( .A1(n15160), .A2(n13244), .ZN(n10258) );
NAND2_X2 U11897 ( .A1(n15146), .A2(n13244), .ZN(n10255) );
NAND2_X2 U11898 ( .A1(n15132), .A2(n13244), .ZN(n10252) );
NAND2_X2 U11899 ( .A1(n15118), .A2(n13244), .ZN(n10249) );
NAND2_X2 U11900 ( .A1(n15104), .A2(n13244), .ZN(n10246) );
NAND2_X2 U11901 ( .A1(n15090), .A2(n13245), .ZN(n10243) );
NAND2_X2 U11902 ( .A1(n15076), .A2(n13245), .ZN(n10240) );
NAND2_X2 U11903 ( .A1(n15062), .A2(n13245), .ZN(n10237) );
NAND2_X2 U11904 ( .A1(n15048), .A2(n13245), .ZN(n10234) );
NAND2_X2 U11905 ( .A1(n15034), .A2(n13245), .ZN(n10231) );
NAND2_X2 U11906 ( .A1(n15020), .A2(n13245), .ZN(n10228) );
NAND2_X2 U11907 ( .A1(n15006), .A2(n13245), .ZN(n10225) );
NAND2_X2 U11908 ( .A1(n14992), .A2(n13245), .ZN(n10222) );
NAND2_X2 U11909 ( .A1(n14978), .A2(n13245), .ZN(n10219) );
NAND2_X2 U11910 ( .A1(n14964), .A2(n13245), .ZN(n10214) );
NAND2_X2 U11911 ( .A1(n14724), .A2(n10212), .ZN(n14709) );
NAND2_X2 U11912 ( .A1(n15411), .A2(n13263), .ZN(n10210) );
NAND2_X2 U11913 ( .A1(n15396), .A2(n13263), .ZN(n10207) );
NAND2_X2 U11914 ( .A1(n15381), .A2(n13263), .ZN(n10204) );
NAND2_X2 U11915 ( .A1(n15366), .A2(n13263), .ZN(n10201) );
NAND2_X2 U11916 ( .A1(n15351), .A2(n13263), .ZN(n10198) );
NAND2_X2 U11917 ( .A1(n15336), .A2(n13263), .ZN(n10195) );
NAND2_X2 U11918 ( .A1(n15321), .A2(n13263), .ZN(n10192) );
NAND2_X2 U11919 ( .A1(n15306), .A2(n13263), .ZN(n10189) );
NAND2_X2 U11920 ( .A1(n15291), .A2(n13263), .ZN(n10186) );
NAND2_X2 U11921 ( .A1(n15276), .A2(n13263), .ZN(n10183) );
NAND2_X2 U11922 ( .A1(n15261), .A2(n13262), .ZN(n10180) );
NAND2_X2 U11923 ( .A1(n15246), .A2(n13262), .ZN(n10177) );
NAND2_X2 U11924 ( .A1(n15231), .A2(n13262), .ZN(n10174) );
NAND2_X2 U11925 ( .A1(n15216), .A2(n13262), .ZN(n10171) );
NAND2_X2 U11926 ( .A1(n15201), .A2(n13262), .ZN(n10168) );
NAND2_X2 U11927 ( .A1(n15187), .A2(n13262), .ZN(n10165) );
NAND2_X2 U11928 ( .A1(n15173), .A2(n13262), .ZN(n10162) );
NAND2_X2 U11929 ( .A1(n15159), .A2(n13262), .ZN(n10159) );
NAND2_X2 U11930 ( .A1(n15145), .A2(n13262), .ZN(n10156) );
NAND2_X2 U11931 ( .A1(n15131), .A2(n13262), .ZN(n10153) );
NAND2_X2 U11932 ( .A1(n15117), .A2(n13262), .ZN(n10150) );
NAND2_X2 U11933 ( .A1(n15103), .A2(n13261), .ZN(n10147) );
NAND2_X2 U11934 ( .A1(n15089), .A2(n13261), .ZN(n10144) );
NAND2_X2 U11935 ( .A1(n15075), .A2(n13261), .ZN(n10141) );
NAND2_X2 U11936 ( .A1(n15061), .A2(n13261), .ZN(n10138) );
NAND2_X2 U11937 ( .A1(n15047), .A2(n13261), .ZN(n10135) );
NAND2_X2 U11938 ( .A1(n15033), .A2(n13261), .ZN(n10132) );
NAND2_X2 U11939 ( .A1(n15019), .A2(n13261), .ZN(n10129) );
NAND2_X2 U11940 ( .A1(n15005), .A2(n13261), .ZN(n10126) );
NAND2_X2 U11941 ( .A1(n14991), .A2(n13261), .ZN(n10123) );
NAND2_X2 U11942 ( .A1(n14977), .A2(n13261), .ZN(n10120) );
NAND2_X2 U11943 ( .A1(n14722), .A2(n14712), .ZN(n10118) );
NAND2_X2 U11944 ( .A1(n14724), .A2(n10118), .ZN(n14710) );
NAND2_X2 U11945 ( .A1(n15410), .A2(n13248), .ZN(n10116) );
NAND2_X2 U11946 ( .A1(n15395), .A2(n13248), .ZN(n10113) );
NAND2_X2 U11947 ( .A1(n15380), .A2(n13248), .ZN(n10110) );
NAND2_X2 U11948 ( .A1(n15365), .A2(n13248), .ZN(n10107) );
NAND2_X2 U11949 ( .A1(n15350), .A2(n13248), .ZN(n10104) );
NAND2_X2 U11950 ( .A1(n15335), .A2(n13248), .ZN(n10101) );
NAND2_X2 U11951 ( .A1(n15320), .A2(n13248), .ZN(n10098) );
NAND2_X2 U11952 ( .A1(n15305), .A2(n13248), .ZN(n10095) );
NAND2_X2 U11953 ( .A1(n15290), .A2(n13248), .ZN(n10092) );
NAND2_X2 U11954 ( .A1(n15275), .A2(n13248), .ZN(n10089) );
NAND2_X2 U11955 ( .A1(n15260), .A2(n13247), .ZN(n10086) );
NAND2_X2 U11956 ( .A1(n15245), .A2(n13247), .ZN(n10083) );
NAND2_X2 U11957 ( .A1(n15230), .A2(n13247), .ZN(n10080) );
NAND2_X2 U11958 ( .A1(n15215), .A2(n13247), .ZN(n10077) );
NAND2_X2 U11959 ( .A1(n15200), .A2(n13247), .ZN(n10074) );
NAND2_X2 U11960 ( .A1(n15186), .A2(n13247), .ZN(n10071) );
NAND2_X2 U11961 ( .A1(n15172), .A2(n13247), .ZN(n10068) );
NAND2_X2 U11962 ( .A1(n15158), .A2(n13247), .ZN(n10065) );
NAND2_X2 U11963 ( .A1(n15144), .A2(n13247), .ZN(n10062) );
NAND2_X2 U11964 ( .A1(n15130), .A2(n13247), .ZN(n10059) );
NAND2_X2 U11965 ( .A1(n15116), .A2(n13247), .ZN(n10056) );
NAND2_X2 U11966 ( .A1(n15102), .A2(n13246), .ZN(n10053) );
NAND2_X2 U11967 ( .A1(n15088), .A2(n13246), .ZN(n10050) );
NAND2_X2 U11968 ( .A1(n15074), .A2(n13246), .ZN(n10047) );
NAND2_X2 U11969 ( .A1(n15060), .A2(n13246), .ZN(n10044) );
NAND2_X2 U11970 ( .A1(n15046), .A2(n13246), .ZN(n10041) );
NAND2_X2 U11971 ( .A1(n15032), .A2(n13246), .ZN(n10038) );
NAND2_X2 U11972 ( .A1(n15018), .A2(n13246), .ZN(n10035) );
NAND2_X2 U11973 ( .A1(n15004), .A2(n13246), .ZN(n10032) );
NAND2_X2 U11974 ( .A1(n14990), .A2(n13246), .ZN(n10029) );
NAND2_X2 U11975 ( .A1(n14976), .A2(n13246), .ZN(n10026) );
NAND2_X2 U11976 ( .A1(n15424), .A2(n13246), .ZN(n10021) );
NAND2_X2 U11977 ( .A1(n14712), .A2(n14727), .ZN(n10019) );
NAND2_X2 U11978 ( .A1(n14724), .A2(n10019), .ZN(n14711) );
NAND2_X2 U11979 ( .A1(n15409), .A2(n13251), .ZN(n10017) );
NAND2_X2 U11980 ( .A1(n15394), .A2(n13251), .ZN(n10014) );
NAND2_X2 U11981 ( .A1(n15379), .A2(n13251), .ZN(n10011) );
NAND2_X2 U11982 ( .A1(n15364), .A2(n13251), .ZN(n10008) );
NAND2_X2 U11983 ( .A1(n15349), .A2(n13251), .ZN(n10005) );
NAND2_X2 U11984 ( .A1(n15334), .A2(n13251), .ZN(n10002) );
NAND2_X2 U11985 ( .A1(n15319), .A2(n13251), .ZN(n9999) );
NAND2_X2 U11986 ( .A1(n15304), .A2(n13251), .ZN(n9996) );
NAND2_X2 U11987 ( .A1(n15289), .A2(n13251), .ZN(n9993) );
NAND2_X2 U11988 ( .A1(n15274), .A2(n13251), .ZN(n9990) );
NAND2_X2 U11989 ( .A1(n15259), .A2(n13250), .ZN(n9987) );
NAND2_X2 U11990 ( .A1(n15244), .A2(n13250), .ZN(n9984) );
NAND2_X2 U11991 ( .A1(n15229), .A2(n13250), .ZN(n9981) );
NAND2_X2 U11992 ( .A1(n15214), .A2(n13250), .ZN(n9978) );
NAND2_X2 U11993 ( .A1(n15199), .A2(n13250), .ZN(n9975) );
NAND2_X2 U11994 ( .A1(n15185), .A2(n13250), .ZN(n9972) );
NAND2_X2 U11995 ( .A1(n15171), .A2(n13250), .ZN(n9969) );
NAND2_X2 U11996 ( .A1(n15157), .A2(n13250), .ZN(n9966) );
NAND2_X2 U11997 ( .A1(n15143), .A2(n13250), .ZN(n9963) );
NAND2_X2 U11998 ( .A1(n15129), .A2(n13250), .ZN(n9960) );
NAND2_X2 U11999 ( .A1(n15115), .A2(n13250), .ZN(n9957) );
NAND2_X2 U12000 ( .A1(n15101), .A2(n13249), .ZN(n9954) );
NAND2_X2 U12001 ( .A1(n15087), .A2(n13249), .ZN(n9951) );
NAND2_X2 U12002 ( .A1(n15073), .A2(n13249), .ZN(n9948) );
NAND2_X2 U12003 ( .A1(n15059), .A2(n13249), .ZN(n9945) );
NAND2_X2 U12004 ( .A1(n15045), .A2(n13249), .ZN(n9942) );
NAND2_X2 U12005 ( .A1(n15031), .A2(n13249), .ZN(n9939) );
NAND2_X2 U12006 ( .A1(n15017), .A2(n13249), .ZN(n9936) );
NAND2_X2 U12007 ( .A1(n15003), .A2(n13249), .ZN(n9933) );
NAND2_X2 U12008 ( .A1(n14989), .A2(n13249), .ZN(n9930) );
NAND2_X2 U12009 ( .A1(n14975), .A2(n13249), .ZN(n9927) );
NAND2_X2 U12010 ( .A1(n15423), .A2(n13249), .ZN(n9922) );
NAND2_X2 U12011 ( .A1(n13028), .A2(n14712), .ZN(n14713) );
NAND2_X2 U12012 ( .A1(n14724), .A2(n14714), .ZN(n14716) );
NAND2_X2 U12013 ( .A1(n15408), .A2(n13252), .ZN(n9916) );
NAND2_X2 U12014 ( .A1(n15393), .A2(n13252), .ZN(n9913) );
NAND2_X2 U12015 ( .A1(n15378), .A2(n13252), .ZN(n9910) );
NAND2_X2 U12016 ( .A1(n15363), .A2(n13252), .ZN(n9907) );
NAND2_X2 U12017 ( .A1(n15348), .A2(n13252), .ZN(n9904) );
NAND2_X2 U12018 ( .A1(n15333), .A2(n13252), .ZN(n9901) );
NAND2_X2 U12019 ( .A1(n15318), .A2(n13252), .ZN(n9898) );
NAND2_X2 U12020 ( .A1(n15303), .A2(n13252), .ZN(n9895) );
NAND2_X2 U12021 ( .A1(n15288), .A2(n13252), .ZN(n9892) );
NAND2_X2 U12022 ( .A1(n15273), .A2(n13252), .ZN(n9889) );
NAND2_X2 U12023 ( .A1(n15258), .A2(n13252), .ZN(n9886) );
NAND2_X2 U12024 ( .A1(n15243), .A2(n13253), .ZN(n9883) );
NAND2_X2 U12025 ( .A1(n15228), .A2(n13253), .ZN(n9880) );
NAND2_X2 U12026 ( .A1(n15213), .A2(n13253), .ZN(n9877) );
NAND2_X2 U12027 ( .A1(n15198), .A2(n13253), .ZN(n9874) );
NAND2_X2 U12028 ( .A1(n15184), .A2(n13253), .ZN(n9871) );
NAND2_X2 U12029 ( .A1(n15170), .A2(n13253), .ZN(n9868) );
NAND2_X2 U12030 ( .A1(n15156), .A2(n13253), .ZN(n9865) );
NAND2_X2 U12031 ( .A1(n15142), .A2(n13253), .ZN(n9862) );
NAND2_X2 U12032 ( .A1(n15128), .A2(n13253), .ZN(n9859) );
NAND2_X2 U12033 ( .A1(n15114), .A2(n13253), .ZN(n9856) );
NAND2_X2 U12034 ( .A1(n15100), .A2(n13253), .ZN(n9853) );
NAND2_X2 U12035 ( .A1(n15086), .A2(n13254), .ZN(n9850) );
NAND2_X2 U12036 ( .A1(n15072), .A2(n13254), .ZN(n9847) );
NAND2_X2 U12037 ( .A1(n15058), .A2(n13254), .ZN(n9844) );
NAND2_X2 U12038 ( .A1(n15044), .A2(n13254), .ZN(n9841) );
NAND2_X2 U12039 ( .A1(n15030), .A2(n13254), .ZN(n9838) );
NAND2_X2 U12040 ( .A1(n15016), .A2(n13254), .ZN(n9835) );
NAND2_X2 U12041 ( .A1(n15002), .A2(n13254), .ZN(n9832) );
NAND2_X2 U12042 ( .A1(n14988), .A2(n13254), .ZN(n9829) );
NAND2_X2 U12043 ( .A1(n14974), .A2(n13254), .ZN(n9826) );
NAND2_X2 U12044 ( .A1(n15422), .A2(n13254), .ZN(n9821) );
INV_X4 U12045 ( .A(n14719), .ZN(n14717) );
NAND2_X2 U12046 ( .A1(n14717), .A2(n14953), .ZN(n14718) );
NAND2_X2 U12047 ( .A1(n14724), .A2(n14719), .ZN(n14720) );
NAND2_X2 U12048 ( .A1(n15407), .A2(n13257), .ZN(n9817) );
NAND2_X2 U12049 ( .A1(n15392), .A2(n13257), .ZN(n9814) );
NAND2_X2 U12050 ( .A1(n15377), .A2(n13257), .ZN(n9811) );
NAND2_X2 U12051 ( .A1(n15362), .A2(n13257), .ZN(n9808) );
NAND2_X2 U12052 ( .A1(n15347), .A2(n13257), .ZN(n9805) );
NAND2_X2 U12053 ( .A1(n15332), .A2(n13257), .ZN(n9802) );
NAND2_X2 U12054 ( .A1(n15317), .A2(n13257), .ZN(n9799) );
NAND2_X2 U12055 ( .A1(n15302), .A2(n13257), .ZN(n9796) );
NAND2_X2 U12056 ( .A1(n15287), .A2(n13257), .ZN(n9793) );
NAND2_X2 U12057 ( .A1(n15272), .A2(n13257), .ZN(n9790) );
NAND2_X2 U12058 ( .A1(n15257), .A2(n13256), .ZN(n9787) );
NAND2_X2 U12059 ( .A1(n15242), .A2(n13256), .ZN(n9784) );
NAND2_X2 U12060 ( .A1(n15227), .A2(n13256), .ZN(n9781) );
NAND2_X2 U12061 ( .A1(n15212), .A2(n13256), .ZN(n9778) );
NAND2_X2 U12062 ( .A1(n15197), .A2(n13256), .ZN(n9775) );
NAND2_X2 U12063 ( .A1(n15183), .A2(n13256), .ZN(n9772) );
NAND2_X2 U12064 ( .A1(n15169), .A2(n13256), .ZN(n9769) );
NAND2_X2 U12065 ( .A1(n15155), .A2(n13256), .ZN(n9766) );
NAND2_X2 U12066 ( .A1(n15141), .A2(n13256), .ZN(n9763) );
NAND2_X2 U12067 ( .A1(n15127), .A2(n13256), .ZN(n9760) );
NAND2_X2 U12068 ( .A1(n15113), .A2(n13256), .ZN(n9757) );
NAND2_X2 U12069 ( .A1(n15099), .A2(n13255), .ZN(n9754) );
NAND2_X2 U12070 ( .A1(n15085), .A2(n13255), .ZN(n9751) );
NAND2_X2 U12071 ( .A1(n15071), .A2(n13255), .ZN(n9748) );
NAND2_X2 U12072 ( .A1(n15057), .A2(n13255), .ZN(n9745) );
NAND2_X2 U12073 ( .A1(n15043), .A2(n13255), .ZN(n9742) );
NAND2_X2 U12074 ( .A1(n15029), .A2(n13255), .ZN(n9739) );
NAND2_X2 U12075 ( .A1(n15015), .A2(n13255), .ZN(n9736) );
NAND2_X2 U12076 ( .A1(n15001), .A2(n13255), .ZN(n9733) );
NAND2_X2 U12077 ( .A1(n14987), .A2(n13255), .ZN(n9730) );
NAND2_X2 U12078 ( .A1(n14973), .A2(n13255), .ZN(n9727) );
NAND2_X2 U12079 ( .A1(n15421), .A2(n13255), .ZN(n9722) );
NAND3_X2 U12080 ( .A1(n14722), .A2(n14953), .A3(n14726), .ZN(n14721) );
NAND2_X2 U12081 ( .A1(n14722), .A2(n14726), .ZN(n14723) );
NAND2_X2 U12082 ( .A1(n14724), .A2(n14723), .ZN(n14725) );
NAND2_X2 U12083 ( .A1(n15406), .A2(n13260), .ZN(n9717) );
NAND2_X2 U12084 ( .A1(n15391), .A2(n13260), .ZN(n9714) );
NAND2_X2 U12085 ( .A1(n15376), .A2(n13260), .ZN(n9711) );
NAND2_X2 U12086 ( .A1(n15361), .A2(n13260), .ZN(n9708) );
NAND2_X2 U12087 ( .A1(n15346), .A2(n13260), .ZN(n9705) );
NAND2_X2 U12088 ( .A1(n15331), .A2(n13260), .ZN(n9702) );
NAND2_X2 U12089 ( .A1(n15316), .A2(n13260), .ZN(n9699) );
NAND2_X2 U12090 ( .A1(n15301), .A2(n13260), .ZN(n9696) );
NAND2_X2 U12091 ( .A1(n15286), .A2(n13260), .ZN(n9693) );
NAND2_X2 U12092 ( .A1(n15271), .A2(n13260), .ZN(n9690) );
NAND2_X2 U12093 ( .A1(n15256), .A2(n13259), .ZN(n9687) );
NAND2_X2 U12094 ( .A1(n15241), .A2(n13259), .ZN(n9684) );
NAND2_X2 U12095 ( .A1(n15226), .A2(n13259), .ZN(n9681) );
NAND2_X2 U12096 ( .A1(n15211), .A2(n13259), .ZN(n9678) );
NAND2_X2 U12097 ( .A1(n15196), .A2(n13259), .ZN(n9675) );
NAND2_X2 U12098 ( .A1(n15182), .A2(n13259), .ZN(n9672) );
NAND2_X2 U12099 ( .A1(n15168), .A2(n13259), .ZN(n9669) );
NAND2_X2 U12100 ( .A1(n15154), .A2(n13259), .ZN(n9666) );
NAND2_X2 U12101 ( .A1(n15140), .A2(n13259), .ZN(n9663) );
NAND2_X2 U12102 ( .A1(n15126), .A2(n13259), .ZN(n9660) );
NAND2_X2 U12103 ( .A1(n15112), .A2(n13259), .ZN(n9657) );
NAND2_X2 U12104 ( .A1(n15098), .A2(n13258), .ZN(n9654) );
NAND2_X2 U12105 ( .A1(n15084), .A2(n13258), .ZN(n9651) );
NAND2_X2 U12106 ( .A1(n15070), .A2(n13258), .ZN(n9648) );
NAND2_X2 U12107 ( .A1(n15056), .A2(n13258), .ZN(n9645) );
NAND2_X2 U12108 ( .A1(n15042), .A2(n13258), .ZN(n9642) );
NAND2_X2 U12109 ( .A1(n15028), .A2(n13258), .ZN(n9639) );
NAND2_X2 U12110 ( .A1(n15014), .A2(n13258), .ZN(n9636) );
NAND2_X2 U12111 ( .A1(n15000), .A2(n13258), .ZN(n9633) );
NAND2_X2 U12112 ( .A1(n14986), .A2(n13258), .ZN(n9630) );
NAND2_X2 U12113 ( .A1(n14972), .A2(n13258), .ZN(n9627) );
NAND2_X2 U12114 ( .A1(n15420), .A2(n13258), .ZN(n9622) );
NAND3_X2 U12115 ( .A1(n14727), .A2(n14953), .A3(n14726), .ZN(n14728) );
NAND2_X2 U12116 ( .A1(n15405), .A2(n13266), .ZN(n9615) );
NAND2_X2 U12117 ( .A1(n15390), .A2(n13266), .ZN(n9612) );
NAND2_X2 U12118 ( .A1(n15375), .A2(n13266), .ZN(n9609) );
NAND2_X2 U12119 ( .A1(n15360), .A2(n13266), .ZN(n9606) );
NAND2_X2 U12120 ( .A1(n15345), .A2(n13266), .ZN(n9603) );
NAND2_X2 U12121 ( .A1(n15330), .A2(n13266), .ZN(n9600) );
NAND2_X2 U12122 ( .A1(n15315), .A2(n13266), .ZN(n9597) );
NAND2_X2 U12123 ( .A1(n15300), .A2(n13266), .ZN(n9594) );
NAND2_X2 U12124 ( .A1(n15285), .A2(n13266), .ZN(n9591) );
NAND2_X2 U12125 ( .A1(n15270), .A2(n13266), .ZN(n9588) );
NAND2_X2 U12126 ( .A1(n15255), .A2(n13265), .ZN(n9585) );
NAND2_X2 U12127 ( .A1(n15240), .A2(n13265), .ZN(n9582) );
NAND2_X2 U12128 ( .A1(n15225), .A2(n13265), .ZN(n9579) );
NAND2_X2 U12129 ( .A1(n15210), .A2(n13265), .ZN(n9576) );
NAND2_X2 U12130 ( .A1(n14963), .A2(n13261), .ZN(n9316) );
NAND2_X2 U12131 ( .A1(n13321), .A2(n14733), .ZN(n9304) );
INV_X4 U12132 ( .A(n9304), .ZN(n14734) );
NAND2_X2 U12133 ( .A1(n14735), .A2(n14734), .ZN(n9303) );
NAND2_X2 U12134 ( .A1(n13334), .A2(SHA1_result[0]), .ZN(n14741) );
NAND2_X2 U12135 ( .A1(n13331), .A2(SHA1_result[32]), .ZN(n14740) );
NAND2_X2 U12136 ( .A1(n13337), .A2(SHA1_result[64]), .ZN(n14739) );
NOR2_X2 U12137 ( .A1(n13340), .A2(n13084), .ZN(n14737) );
NOR2_X2 U12138 ( .A1(n13343), .A2(n12851), .ZN(n14736) );
NOR3_X2 U12139 ( .A1(n11853), .A2(n14737), .A3(n14736), .ZN(n14738) );
NAND4_X2 U12140 ( .A1(n14741), .A2(n14740), .A3(n14739), .A4(n14738), .ZN(n3693) );
NAND2_X2 U12141 ( .A1(n13334), .A2(SHA1_result[1]), .ZN(n14749) );
NAND2_X2 U12142 ( .A1(n13331), .A2(n14742), .ZN(n14748) );
NAND2_X2 U12143 ( .A1(n13337), .A2(SHA1_result[65]), .ZN(n14747) );
NOR2_X2 U12144 ( .A1(n13340), .A2(n14743), .ZN(n14745) );
NOR2_X2 U12145 ( .A1(n13343), .A2(n12853), .ZN(n14744) );
NOR3_X2 U12146 ( .A1(n11865), .A2(n14745), .A3(n14744), .ZN(n14746) );
NAND4_X2 U12147 ( .A1(n14749), .A2(n14748), .A3(n14747), .A4(n14746), .ZN(n3692) );
NAND2_X2 U12148 ( .A1(n13334), .A2(SHA1_result[2]), .ZN(n14756) );
NAND2_X2 U12149 ( .A1(n13331), .A2(SHA1_result[34]), .ZN(n14755) );
NAND2_X2 U12150 ( .A1(n13337), .A2(SHA1_result[66]), .ZN(n14754) );
NOR2_X2 U12151 ( .A1(n13340), .A2(n14750), .ZN(n14752) );
NOR2_X2 U12152 ( .A1(n13343), .A2(n12855), .ZN(n14751) );
NOR3_X2 U12153 ( .A1(n11872), .A2(n14752), .A3(n14751), .ZN(n14753) );
NAND4_X2 U12154 ( .A1(n14756), .A2(n14755), .A3(n14754), .A4(n14753), .ZN(n3691) );
NAND2_X2 U12155 ( .A1(n13334), .A2(SHA1_result[3]), .ZN(n14763) );
NAND2_X2 U12156 ( .A1(n13331), .A2(SHA1_result[35]), .ZN(n14762) );
NAND2_X2 U12157 ( .A1(n13337), .A2(SHA1_result[67]), .ZN(n14761) );
NOR2_X2 U12158 ( .A1(n13340), .A2(n14757), .ZN(n14759) );
NOR2_X2 U12159 ( .A1(n13343), .A2(n12857), .ZN(n14758) );
NOR3_X2 U12160 ( .A1(n11879), .A2(n14759), .A3(n14758), .ZN(n14760) );
NAND4_X2 U12161 ( .A1(n14763), .A2(n14762), .A3(n14761), .A4(n14760), .ZN(n3690) );
NAND2_X2 U12162 ( .A1(n13334), .A2(SHA1_result[4]), .ZN(n14769) );
NAND2_X2 U12163 ( .A1(n13331), .A2(SHA1_result[36]), .ZN(n14768) );
NAND2_X2 U12164 ( .A1(n13337), .A2(SHA1_result[68]), .ZN(n14767) );
NOR2_X2 U12165 ( .A1(n13340), .A2(n13015), .ZN(n14765) );
NOR2_X2 U12166 ( .A1(n13343), .A2(n12859), .ZN(n14764) );
NOR3_X2 U12167 ( .A1(n11886), .A2(n14765), .A3(n14764), .ZN(n14766) );
NAND4_X2 U12168 ( .A1(n14769), .A2(n14768), .A3(n14767), .A4(n14766), .ZN(n3689) );
NAND2_X2 U12169 ( .A1(n13334), .A2(SHA1_result[5]), .ZN(n14777) );
NAND2_X2 U12170 ( .A1(n13331), .A2(n14770), .ZN(n14776) );
NAND2_X2 U12171 ( .A1(n13337), .A2(SHA1_result[69]), .ZN(n14775) );
NOR2_X2 U12172 ( .A1(n13340), .A2(n14771), .ZN(n14773) );
NOR2_X2 U12173 ( .A1(n13343), .A2(n12861), .ZN(n14772) );
NOR3_X2 U12174 ( .A1(n11893), .A2(n14773), .A3(n14772), .ZN(n14774) );
NAND4_X2 U12175 ( .A1(n14777), .A2(n14776), .A3(n14775), .A4(n14774), .ZN(n3688) );
NAND2_X2 U12176 ( .A1(n13334), .A2(SHA1_result[6]), .ZN(n14784) );
NAND2_X2 U12177 ( .A1(n13331), .A2(n14778), .ZN(n14783) );
NAND2_X2 U12178 ( .A1(n13337), .A2(SHA1_result[70]), .ZN(n14782) );
NOR2_X2 U12179 ( .A1(n13340), .A2(n13000), .ZN(n14780) );
NOR2_X2 U12180 ( .A1(n13343), .A2(n12863), .ZN(n14779) );
NOR3_X2 U12181 ( .A1(n11900), .A2(n14780), .A3(n14779), .ZN(n14781) );
NAND4_X2 U12182 ( .A1(n14784), .A2(n14783), .A3(n14782), .A4(n14781), .ZN(n3687) );
NAND2_X2 U12183 ( .A1(n13334), .A2(SHA1_result[7]), .ZN(n14790) );
NAND2_X2 U12184 ( .A1(n13331), .A2(SHA1_result[39]), .ZN(n14789) );
NAND2_X2 U12185 ( .A1(n13337), .A2(SHA1_result[71]), .ZN(n14788) );
NOR2_X2 U12186 ( .A1(n13340), .A2(n13019), .ZN(n14786) );
NOR2_X2 U12187 ( .A1(n13343), .A2(n12865), .ZN(n14785) );
NOR3_X2 U12188 ( .A1(n11907), .A2(n14786), .A3(n14785), .ZN(n14787) );
NAND4_X2 U12189 ( .A1(n14790), .A2(n14789), .A3(n14788), .A4(n14787), .ZN(n3686) );
NAND2_X2 U12190 ( .A1(n13334), .A2(SHA1_result[8]), .ZN(n14796) );
NAND2_X2 U12191 ( .A1(n13331), .A2(SHA1_result[40]), .ZN(n14795) );
NAND2_X2 U12192 ( .A1(n13337), .A2(SHA1_result[72]), .ZN(n14794) );
NOR2_X2 U12193 ( .A1(n13340), .A2(n13020), .ZN(n14792) );
NOR2_X2 U12194 ( .A1(n13343), .A2(n12867), .ZN(n14791) );
NOR3_X2 U12195 ( .A1(n11914), .A2(n14792), .A3(n14791), .ZN(n14793) );
NAND4_X2 U12196 ( .A1(n14796), .A2(n14795), .A3(n14794), .A4(n14793), .ZN(n3685) );
NAND2_X2 U12197 ( .A1(n13334), .A2(SHA1_result[9]), .ZN(n14803) );
NAND2_X2 U12198 ( .A1(n13331), .A2(n14797), .ZN(n14802) );
NAND2_X2 U12199 ( .A1(n13337), .A2(SHA1_result[73]), .ZN(n14801) );
NOR2_X2 U12200 ( .A1(n13340), .A2(n13079), .ZN(n14799) );
NOR2_X2 U12201 ( .A1(n13343), .A2(n12869), .ZN(n14798) );
NOR3_X2 U12202 ( .A1(n11921), .A2(n14799), .A3(n14798), .ZN(n14800) );
NAND4_X2 U12203 ( .A1(n14803), .A2(n14802), .A3(n14801), .A4(n14800), .ZN(n3684) );
NAND2_X2 U12204 ( .A1(n13333), .A2(SHA1_result[10]), .ZN(n14809) );
NAND2_X2 U12205 ( .A1(n13330), .A2(SHA1_result[42]), .ZN(n14808) );
NAND2_X2 U12206 ( .A1(n13337), .A2(SHA1_result[74]), .ZN(n14807) );
NOR2_X2 U12207 ( .A1(n13339), .A2(n13098), .ZN(n14805) );
NOR2_X2 U12208 ( .A1(n13343), .A2(n12871), .ZN(n14804) );
NOR3_X2 U12209 ( .A1(n11928), .A2(n14805), .A3(n14804), .ZN(n14806) );
NAND4_X2 U12210 ( .A1(n14809), .A2(n14808), .A3(n14807), .A4(n14806), .ZN(n3683) );
NAND2_X2 U12211 ( .A1(n13333), .A2(SHA1_result[11]), .ZN(n14816) );
NAND2_X2 U12212 ( .A1(n13330), .A2(n14810), .ZN(n14815) );
NAND2_X2 U12213 ( .A1(n13338), .A2(SHA1_result[75]), .ZN(n14814) );
NOR2_X2 U12214 ( .A1(n13339), .A2(n13001), .ZN(n14812) );
NOR2_X2 U12215 ( .A1(n13344), .A2(n12873), .ZN(n14811) );
NOR3_X2 U12216 ( .A1(n11935), .A2(n14812), .A3(n14811), .ZN(n14813) );
NAND4_X2 U12217 ( .A1(n14816), .A2(n14815), .A3(n14814), .A4(n14813), .ZN(n3682) );
NAND2_X2 U12218 ( .A1(n13333), .A2(SHA1_result[12]), .ZN(n14823) );
NAND2_X2 U12219 ( .A1(n13330), .A2(n14817), .ZN(n14822) );
NAND2_X2 U12220 ( .A1(n13338), .A2(SHA1_result[76]), .ZN(n14821) );
NOR2_X2 U12221 ( .A1(n13339), .A2(n13016), .ZN(n14819) );
NOR2_X2 U12222 ( .A1(n13344), .A2(n12875), .ZN(n14818) );
NOR3_X2 U12223 ( .A1(n11942), .A2(n14819), .A3(n14818), .ZN(n14820) );
NAND4_X2 U12224 ( .A1(n14823), .A2(n14822), .A3(n14821), .A4(n14820), .ZN(n3681) );
NAND2_X2 U12225 ( .A1(n13333), .A2(SHA1_result[13]), .ZN(n14829) );
NAND2_X2 U12226 ( .A1(n13330), .A2(SHA1_result[45]), .ZN(n14828) );
NAND2_X2 U12227 ( .A1(n13338), .A2(SHA1_result[77]), .ZN(n14827) );
NOR2_X2 U12228 ( .A1(n13339), .A2(n13022), .ZN(n14825) );
NOR2_X2 U12229 ( .A1(n13344), .A2(n12877), .ZN(n14824) );
NOR3_X2 U12230 ( .A1(n11949), .A2(n14825), .A3(n14824), .ZN(n14826) );
NAND4_X2 U12231 ( .A1(n14829), .A2(n14828), .A3(n14827), .A4(n14826), .ZN(n3680) );
NAND2_X2 U12232 ( .A1(n13333), .A2(SHA1_result[14]), .ZN(n14836) );
NAND2_X2 U12233 ( .A1(n13330), .A2(n14830), .ZN(n14835) );
NAND2_X2 U12234 ( .A1(n13338), .A2(SHA1_result[78]), .ZN(n14834) );
NOR2_X2 U12235 ( .A1(n13339), .A2(n13005), .ZN(n14832) );
NOR2_X2 U12236 ( .A1(n13344), .A2(n12879), .ZN(n14831) );
NOR3_X2 U12237 ( .A1(n11956), .A2(n14832), .A3(n14831), .ZN(n14833) );
NAND4_X2 U12238 ( .A1(n14836), .A2(n14835), .A3(n14834), .A4(n14833), .ZN(n3679) );
NAND2_X2 U12239 ( .A1(n13333), .A2(SHA1_result[15]), .ZN(n14842) );
NAND2_X2 U12240 ( .A1(n13330), .A2(SHA1_result[47]), .ZN(n14841) );
NAND2_X2 U12241 ( .A1(n13338), .A2(SHA1_result[79]), .ZN(n14840) );
NOR2_X2 U12242 ( .A1(n13339), .A2(n13021), .ZN(n14838) );
NOR2_X2 U12243 ( .A1(n13344), .A2(n12881), .ZN(n14837) );
NOR3_X2 U12244 ( .A1(n11963), .A2(n14838), .A3(n14837), .ZN(n14839) );
NAND4_X2 U12245 ( .A1(n14842), .A2(n14841), .A3(n14840), .A4(n14839), .ZN(n3678) );
NAND2_X2 U12246 ( .A1(n13333), .A2(SHA1_result[16]), .ZN(n14848) );
NAND2_X2 U12247 ( .A1(n13330), .A2(SHA1_result[48]), .ZN(n14847) );
NAND2_X2 U12248 ( .A1(n13338), .A2(SHA1_result[80]), .ZN(n14846) );
NOR2_X2 U12249 ( .A1(n13339), .A2(n13018), .ZN(n14844) );
NOR2_X2 U12250 ( .A1(n13344), .A2(n12883), .ZN(n14843) );
NOR3_X2 U12251 ( .A1(n11970), .A2(n14844), .A3(n14843), .ZN(n14845) );
NAND4_X2 U12252 ( .A1(n14848), .A2(n14847), .A3(n14846), .A4(n14845), .ZN(n3677) );
NAND2_X2 U12253 ( .A1(n13333), .A2(SHA1_result[17]), .ZN(n14854) );
NAND2_X2 U12254 ( .A1(n13330), .A2(SHA1_result[49]), .ZN(n14853) );
NAND2_X2 U12255 ( .A1(n13338), .A2(SHA1_result[81]), .ZN(n14852) );
NOR2_X2 U12256 ( .A1(n13339), .A2(n13023), .ZN(n14850) );
NOR2_X2 U12257 ( .A1(n13344), .A2(n12885), .ZN(n14849) );
NOR3_X2 U12258 ( .A1(n11977), .A2(n14850), .A3(n14849), .ZN(n14851) );
NAND4_X2 U12259 ( .A1(n14854), .A2(n14853), .A3(n14852), .A4(n14851), .ZN(n3676) );
NAND2_X2 U12260 ( .A1(n13333), .A2(SHA1_result[18]), .ZN(n14860) );
NAND2_X2 U12261 ( .A1(n13330), .A2(SHA1_result[50]), .ZN(n14859) );
NAND2_X2 U12262 ( .A1(n13338), .A2(SHA1_result[82]), .ZN(n14858) );
NOR2_X2 U12263 ( .A1(n13339), .A2(n13004), .ZN(n14856) );
NOR2_X2 U12264 ( .A1(n13344), .A2(n12887), .ZN(n14855) );
NOR3_X2 U12265 ( .A1(n11984), .A2(n14856), .A3(n14855), .ZN(n14857) );
NAND4_X2 U12266 ( .A1(n14860), .A2(n14859), .A3(n14858), .A4(n14857), .ZN(n3675) );
NAND2_X2 U12267 ( .A1(n13333), .A2(SHA1_result[19]), .ZN(n14867) );
NAND2_X2 U12268 ( .A1(n13330), .A2(SHA1_result[51]), .ZN(n14866) );
NAND2_X2 U12269 ( .A1(n13338), .A2(SHA1_result[83]), .ZN(n14865) );
NOR2_X2 U12270 ( .A1(n13339), .A2(n14861), .ZN(n14863) );
NOR2_X2 U12271 ( .A1(n13344), .A2(n12889), .ZN(n14862) );
NOR3_X2 U12272 ( .A1(n11991), .A2(n14863), .A3(n14862), .ZN(n14864) );
NAND4_X2 U12273 ( .A1(n14867), .A2(n14866), .A3(n14865), .A4(n14864), .ZN(n3674) );
NAND2_X2 U12274 ( .A1(n13333), .A2(SHA1_result[20]), .ZN(n14874) );
NAND2_X2 U12275 ( .A1(n13330), .A2(n14868), .ZN(n14873) );
NAND2_X2 U12276 ( .A1(n13338), .A2(SHA1_result[84]), .ZN(n14872) );
NOR2_X2 U12277 ( .A1(n13339), .A2(n13012), .ZN(n14870) );
NOR2_X2 U12278 ( .A1(n13344), .A2(n12891), .ZN(n14869) );
NOR3_X2 U12279 ( .A1(n11998), .A2(n14870), .A3(n14869), .ZN(n14871) );
NAND4_X2 U12280 ( .A1(n14874), .A2(n14873), .A3(n14872), .A4(n14871), .ZN(n3673) );
NAND2_X2 U12281 ( .A1(n13063), .A2(n13269), .ZN(n14877) );
NAND2_X2 U12282 ( .A1(n13265), .A2(n14951), .ZN(n14876) );
NAND2_X2 U12283 ( .A1(n13317), .A2(Wt[0]), .ZN(n14875) );
NAND3_X2 U12284 ( .A1(n14877), .A2(n14876), .A3(n14875), .ZN(n4495) );
NAND2_X2 U12285 ( .A1(n13046), .A2(n13269), .ZN(n14880) );
NAND2_X2 U12286 ( .A1(n13265), .A2(n14950), .ZN(n14879) );
NAND2_X2 U12287 ( .A1(n13317), .A2(Wt[17]), .ZN(n14878) );
NAND3_X2 U12288 ( .A1(n14880), .A2(n14879), .A3(n14878), .ZN(n4478) );
NAND2_X2 U12289 ( .A1(n13047), .A2(n13269), .ZN(n14883) );
NAND2_X2 U12290 ( .A1(n13265), .A2(n14949), .ZN(n14882) );
NAND2_X2 U12291 ( .A1(n13317), .A2(Wt[16]), .ZN(n14881) );
NAND3_X2 U12292 ( .A1(n14883), .A2(n14882), .A3(n14881), .ZN(n4479) );
NAND2_X2 U12293 ( .A1(n13048), .A2(n13269), .ZN(n14886) );
NAND2_X2 U12294 ( .A1(n13265), .A2(n14948), .ZN(n14885) );
NAND2_X2 U12295 ( .A1(n13317), .A2(Wt[15]), .ZN(n14884) );
NAND3_X2 U12296 ( .A1(n14886), .A2(n14885), .A3(n14884), .ZN(n4480) );
NAND2_X2 U12297 ( .A1(n13049), .A2(n13269), .ZN(n14889) );
NAND2_X2 U12298 ( .A1(n13265), .A2(n14947), .ZN(n14888) );
NAND2_X2 U12299 ( .A1(n13317), .A2(Wt[14]), .ZN(n14887) );
NAND3_X2 U12300 ( .A1(n14889), .A2(n14888), .A3(n14887), .ZN(n4481) );
NAND2_X2 U12301 ( .A1(n13050), .A2(n13269), .ZN(n14892) );
NAND2_X2 U12302 ( .A1(n13265), .A2(n14946), .ZN(n14891) );
NAND2_X2 U12303 ( .A1(n13317), .A2(Wt[13]), .ZN(n14890) );
NAND3_X2 U12304 ( .A1(n14892), .A2(n14891), .A3(n14890), .ZN(n4482) );
NAND2_X2 U12305 ( .A1(n13051), .A2(n13269), .ZN(n14895) );
NAND2_X2 U12306 ( .A1(n13265), .A2(n14945), .ZN(n14894) );
NAND2_X2 U12307 ( .A1(n13314), .A2(Wt[12]), .ZN(n14893) );
NAND3_X2 U12308 ( .A1(n14895), .A2(n14894), .A3(n14893), .ZN(n4483) );
NAND2_X2 U12309 ( .A1(n13052), .A2(n13269), .ZN(n14898) );
NAND2_X2 U12310 ( .A1(n13264), .A2(n14944), .ZN(n14897) );
NAND2_X2 U12311 ( .A1(n13273), .A2(Wt[11]), .ZN(n14896) );
NAND3_X2 U12312 ( .A1(n14898), .A2(n14897), .A3(n14896), .ZN(n4484) );
NAND2_X2 U12313 ( .A1(n13053), .A2(n13269), .ZN(n14901) );
NAND2_X2 U12314 ( .A1(n13264), .A2(n14943), .ZN(n14900) );
NAND2_X2 U12315 ( .A1(n13272), .A2(Wt[10]), .ZN(n14899) );
NAND3_X2 U12316 ( .A1(n14901), .A2(n14900), .A3(n14899), .ZN(n4485) );
NAND2_X2 U12317 ( .A1(n13054), .A2(n13269), .ZN(n14904) );
NAND2_X2 U12318 ( .A1(n13264), .A2(n14942), .ZN(n14903) );
NAND2_X2 U12319 ( .A1(n13315), .A2(Wt[9]), .ZN(n14902) );
NAND3_X2 U12320 ( .A1(n14904), .A2(n14903), .A3(n14902), .ZN(n4486) );
NAND2_X2 U12321 ( .A1(n13055), .A2(n13268), .ZN(n14907) );
NAND2_X2 U12322 ( .A1(n13264), .A2(n14941), .ZN(n14906) );
NAND2_X2 U12323 ( .A1(n13315), .A2(Wt[8]), .ZN(n14905) );
NAND3_X2 U12324 ( .A1(n14907), .A2(n14906), .A3(n14905), .ZN(n4487) );
NAND2_X2 U12325 ( .A1(n13056), .A2(n13268), .ZN(n14910) );
NAND2_X2 U12326 ( .A1(n13264), .A2(n14940), .ZN(n14909) );
NAND2_X2 U12327 ( .A1(n13315), .A2(Wt[7]), .ZN(n14908) );
NAND3_X2 U12328 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(n4488) );
NAND2_X2 U12329 ( .A1(n13057), .A2(n13268), .ZN(n14913) );
NAND2_X2 U12330 ( .A1(n13264), .A2(n14939), .ZN(n14912) );
NAND2_X2 U12331 ( .A1(n13315), .A2(Wt[6]), .ZN(n14911) );
NAND3_X2 U12332 ( .A1(n14913), .A2(n14912), .A3(n14911), .ZN(n4489) );
NAND2_X2 U12333 ( .A1(n13058), .A2(n13268), .ZN(n14916) );
NAND2_X2 U12334 ( .A1(n13264), .A2(n14938), .ZN(n14915) );
NAND2_X2 U12335 ( .A1(n13315), .A2(Wt[5]), .ZN(n14914) );
NAND3_X2 U12336 ( .A1(n14916), .A2(n14915), .A3(n14914), .ZN(n4490) );
NAND2_X2 U12337 ( .A1(n13059), .A2(n13268), .ZN(n14919) );
NAND2_X2 U12338 ( .A1(n13264), .A2(n14937), .ZN(n14918) );
NAND2_X2 U12339 ( .A1(n13315), .A2(Wt[4]), .ZN(n14917) );
NAND3_X2 U12340 ( .A1(n14919), .A2(n14918), .A3(n14917), .ZN(n4491) );
NAND2_X2 U12341 ( .A1(n13060), .A2(n13268), .ZN(n14922) );
NAND2_X2 U12342 ( .A1(n13264), .A2(n14936), .ZN(n14921) );
NAND2_X2 U12343 ( .A1(n13315), .A2(Wt[3]), .ZN(n14920) );
NAND3_X2 U12344 ( .A1(n14922), .A2(n14921), .A3(n14920), .ZN(n4492) );
NAND2_X2 U12345 ( .A1(n13061), .A2(n13268), .ZN(n14925) );
NAND2_X2 U12346 ( .A1(n13264), .A2(n14935), .ZN(n14924) );
NAND2_X2 U12347 ( .A1(n13315), .A2(Wt[2]), .ZN(n14923) );
NAND3_X2 U12348 ( .A1(n14925), .A2(n14924), .A3(n14923), .ZN(n4493) );
NAND2_X2 U12349 ( .A1(n13062), .A2(n13268), .ZN(n14928) );
NAND2_X2 U12350 ( .A1(n13264), .A2(n14934), .ZN(n14927) );
NAND2_X2 U12351 ( .A1(n13315), .A2(Wt[1]), .ZN(n14926) );
NAND3_X2 U12352 ( .A1(n14928), .A2(n14927), .A3(n14926), .ZN(n4494) );
INV_X4 U12353 ( .A(n11837), .ZN(n14954) );
INV_X4 U12354 ( .A(n12076), .ZN(n14956) );
INV_X4 U12355 ( .A(n12077), .ZN(n14957) );
INV_X4 U12356 ( .A(n9309), .ZN(n14958) );
INV_X4 U12357 ( .A(n11840), .ZN(n15425) );
INV_X4 U12358 ( .A(cmd_w_i), .ZN(n15426) );
NAND2_X2 _add_3_root_add_136_4_U427  ( .A1(SHA1_ft_BCD[10]), .A2(SHA1_result_133), .ZN(_add_3_root_add_136_4_n357 ) );
NOR2_X4 _add_3_root_add_136_4_U426  ( .A1(_add_3_root_add_136_4_n30 ), .A2(_add_3_root_add_136_4_n401 ), .ZN(_add_3_root_add_136_4_n394 ) );
INV_X4 _add_3_root_add_136_4_U425  ( .A(n14930), .ZN(_add_3_root_add_136_4_n398 ) );
INV_X4 _add_3_root_add_136_4_U424  ( .A(SHA1_result_128), .ZN(_add_3_root_add_136_4_n399 ) );
INV_X4 _add_3_root_add_136_4_U423  ( .A(_add_3_root_add_136_4_n112 ), .ZN(_add_3_root_add_136_4_n387 ) );
INV_X4 _add_3_root_add_136_4_U422  ( .A(SHA1_result_131), .ZN(_add_3_root_add_136_4_n393 ) );
INV_X4 _add_3_root_add_136_4_U421  ( .A(SHA1_ft_BCD[9]), .ZN(_add_3_root_add_136_4_n390 ) );
INV_X4 _add_3_root_add_136_4_U420  ( .A(SHA1_result_132), .ZN(_add_3_root_add_136_4_n391 ) );
NAND3_X4 _add_3_root_add_136_4_U419  ( .A1(_add_3_root_add_136_4_n108 ),.A2(_add_3_root_add_136_4_n386 ), .A3(_add_3_root_add_136_4_n111 ),.ZN(_add_3_root_add_136_4_n102 ) );
INV_X4 _add_3_root_add_136_4_U418  ( .A(_add_3_root_add_136_4_n315 ), .ZN(_add_3_root_add_136_4_n381 ) );
INV_X4 _add_3_root_add_136_4_U417  ( .A(n14385), .ZN(_add_3_root_add_136_4_n385 ) );
INV_X4 _add_3_root_add_136_4_U416  ( .A(SHA1_ft_BCD[3]), .ZN(_add_3_root_add_136_4_n382 ) );
INV_X4 _add_3_root_add_136_4_U415  ( .A(n14382), .ZN(_add_3_root_add_136_4_n383 ) );
NAND3_X4 _add_3_root_add_136_4_U414  ( .A1(_add_3_root_add_136_4_n378 ),.A2(_add_3_root_add_136_4_n164 ), .A3(_add_3_root_add_136_4_n380 ),.ZN(_add_3_root_add_136_4_n316 ) );
NOR2_X4 _add_3_root_add_136_4_U413  ( .A1(_add_3_root_add_136_4_n381 ), .A2(_add_3_root_add_136_4_n316 ), .ZN(_add_3_root_add_136_4_n377 ) );
NOR2_X4 _add_3_root_add_136_4_U412  ( .A1(_add_3_root_add_136_4_n123 ), .A2(_add_3_root_add_136_4_n162 ), .ZN(_add_3_root_add_136_4_n317 ) );
NAND3_X4 _add_3_root_add_136_4_U411  ( .A1(_add_3_root_add_136_4_n189 ),.A2(_add_3_root_add_136_4_n376 ), .A3(_add_3_root_add_136_4_n375 ),.ZN(_add_3_root_add_136_4_n374 ) );
NAND3_X4 _add_3_root_add_136_4_U410  ( .A1(_add_3_root_add_136_4_n373 ),.A2(_add_3_root_add_136_4_n93 ), .A3(_add_3_root_add_136_4_n374 ),.ZN(_add_3_root_add_136_4_n371 ) );
INV_X4 _add_3_root_add_136_4_U409  ( .A(SHA1_ft_BCD[11]), .ZN(_add_3_root_add_136_4_n368 ) );
INV_X4 _add_3_root_add_136_4_U408  ( .A(SHA1_result_134), .ZN(_add_3_root_add_136_4_n369 ) );
NAND2_X2 _add_3_root_add_136_4_U407  ( .A1(SHA1_ft_BCD[11]), .A2(SHA1_result_134), .ZN(_add_3_root_add_136_4_n356 ) );
NAND2_X2 _add_3_root_add_136_4_U406  ( .A1(_add_3_root_add_136_4_n327 ),.A2(_add_3_root_add_136_4_n356 ), .ZN(_add_3_root_add_136_4_n367 ) );
XNOR2_X2 _add_3_root_add_136_4_U405  ( .A(_add_3_root_add_136_4_n366 ), .B(_add_3_root_add_136_4_n367 ), .ZN(N75) );
NAND2_X2 _add_3_root_add_136_4_U404  ( .A1(_add_3_root_add_136_4_n95 ), .A2(_add_3_root_add_136_4_n93 ), .ZN(_add_3_root_add_136_4_n360 ) );
INV_X4 _add_3_root_add_136_4_U403  ( .A(SHA1_result_135), .ZN(_add_3_root_add_136_4_n354 ) );
NOR3_X4 _add_3_root_add_136_4_U402  ( .A1(_add_3_root_add_136_4_n105 ), .A2(_add_3_root_add_136_4_n100 ), .A3(_add_3_root_add_136_4_n352 ), .ZN(_add_3_root_add_136_4_n342 ) );
NAND2_X2 _add_3_root_add_136_4_U401  ( .A1(_add_3_root_add_136_4_n5 ), .A2(_add_3_root_add_136_4_n322 ), .ZN(_add_3_root_add_136_4_n349 ) );
NAND2_X2 _add_3_root_add_136_4_U400  ( .A1(_add_3_root_add_136_4_n34 ), .A2(n14443), .ZN(_add_3_root_add_136_4_n340 ) );
INV_X4 _add_3_root_add_136_4_U399  ( .A(_add_3_root_add_136_4_n340 ), .ZN(_add_3_root_add_136_4_n324 ) );
XNOR2_X2 _add_3_root_add_136_4_U398  ( .A(_add_3_root_add_136_4_n344 ), .B(_add_3_root_add_136_4_n345 ), .ZN(N78) );
NAND2_X2 _add_3_root_add_136_4_U397  ( .A1(_add_3_root_add_136_4_n76 ), .A2(_add_3_root_add_136_4_n341 ), .ZN(_add_3_root_add_136_4_n339 ) );
NAND2_X2 _add_3_root_add_136_4_U396  ( .A1(_add_3_root_add_136_4_n339 ),.A2(_add_3_root_add_136_4_n340 ), .ZN(_add_3_root_add_136_4_n338 ) );
NOR2_X4 _add_3_root_add_136_4_U395  ( .A1(_add_3_root_add_136_4_n337 ), .A2(_add_3_root_add_136_4_n338 ), .ZN(_add_3_root_add_136_4_n333 ) );
INV_X4 _add_3_root_add_136_4_U394  ( .A(SHA1_ft_BCD[15]), .ZN(_add_3_root_add_136_4_n335 ) );
INV_X4 _add_3_root_add_136_4_U393  ( .A(n14440), .ZN(_add_3_root_add_136_4_n336 ) );
NAND2_X2 _add_3_root_add_136_4_U392  ( .A1(_add_3_root_add_136_4_n335 ),.A2(_add_3_root_add_136_4_n336 ), .ZN(_add_3_root_add_136_4_n320 ) );
INV_X4 _add_3_root_add_136_4_U391  ( .A(_add_3_root_add_136_4_n320 ), .ZN(_add_3_root_add_136_4_n331 ) );
XNOR2_X2 _add_3_root_add_136_4_U390  ( .A(_add_3_root_add_136_4_n333 ), .B(_add_3_root_add_136_4_n334 ), .ZN(N79) );
NAND2_X2 _add_3_root_add_136_4_U389  ( .A1(SHA1_ft_BCD[16]), .A2(n14437),.ZN(_add_3_root_add_136_4_n305 ) );
NOR2_X4 _add_3_root_add_136_4_U388  ( .A1(n14437), .A2(SHA1_ft_BCD[16]),.ZN(_add_3_root_add_136_4_n297 ) );
INV_X4 _add_3_root_add_136_4_U387  ( .A(_add_3_root_add_136_4_n297 ), .ZN(_add_3_root_add_136_4_n332 ) );
NAND2_X2 _add_3_root_add_136_4_U386  ( .A1(_add_3_root_add_136_4_n305 ),.A2(_add_3_root_add_136_4_n332 ), .ZN(_add_3_root_add_136_4_n307 ) );
NOR3_X4 _add_3_root_add_136_4_U385  ( .A1(_add_3_root_add_136_4_n323 ), .A2(_add_3_root_add_136_4_n324 ), .A3(_add_3_root_add_136_4_n85 ), .ZN(_add_3_root_add_136_4_n321 ) );
INV_X4 _add_3_root_add_136_4_U384  ( .A(_add_3_root_add_136_4_n183 ), .ZN(_add_3_root_add_136_4_n318 ) );
NOR2_X4 _add_3_root_add_136_4_U383  ( .A1(_add_3_root_add_136_4_n37 ), .A2(_add_3_root_add_136_4_n318 ), .ZN(_add_3_root_add_136_4_n308 ) );
NAND2_X2 _add_3_root_add_136_4_U382  ( .A1(_add_3_root_add_136_4_n314 ),.A2(_add_3_root_add_136_4_n315 ), .ZN(_add_3_root_add_136_4_n313 ) );
NAND2_X2 _add_3_root_add_136_4_U381  ( .A1(_add_3_root_add_136_4_n312 ),.A2(_add_3_root_add_136_4_n313 ), .ZN(_add_3_root_add_136_4_n188 ) );
NAND3_X2 _add_3_root_add_136_4_U380  ( .A1(_add_3_root_add_136_4_n189 ),.A2(_add_3_root_add_136_4_n188 ), .A3(_add_3_root_add_136_4_n311 ),.ZN(_add_3_root_add_136_4_n309 ) );
NAND3_X4 _add_3_root_add_136_4_U379  ( .A1(_add_3_root_add_136_4_n308 ),.A2(_add_3_root_add_136_4_n309 ), .A3(_add_3_root_add_136_4_n185 ),.ZN(_add_3_root_add_136_4_n241 ) );
XNOR2_X2 _add_3_root_add_136_4_U378  ( .A(_add_3_root_add_136_4_n241 ), .B(_add_3_root_add_136_4_n307 ), .ZN(N80) );
NAND2_X2 _add_3_root_add_136_4_U377  ( .A1(_add_3_root_add_136_4_n305 ),.A2(_add_3_root_add_136_4_n306 ), .ZN(_add_3_root_add_136_4_n301 ) );
INV_X4 _add_3_root_add_136_4_U376  ( .A(SHA1_ft_BCD[17]), .ZN(_add_3_root_add_136_4_n303 ) );
INV_X4 _add_3_root_add_136_4_U375  ( .A(n14434), .ZN(_add_3_root_add_136_4_n304 ) );
XNOR2_X2 _add_3_root_add_136_4_U374  ( .A(_add_3_root_add_136_4_n301 ), .B(_add_3_root_add_136_4_n302 ), .ZN(N81) );
NAND2_X2 _add_3_root_add_136_4_U373  ( .A1(_add_3_root_add_136_4_n299 ),.A2(_add_3_root_add_136_4_n300 ), .ZN(_add_3_root_add_136_4_n290 ) );
NAND2_X2 _add_3_root_add_136_4_U372  ( .A1(_add_3_root_add_136_4_n286 ),.A2(_add_3_root_add_136_4_n241 ), .ZN(_add_3_root_add_136_4_n295 ) );
INV_X4 _add_3_root_add_136_4_U371  ( .A(SHA1_ft_BCD[18]), .ZN(_add_3_root_add_136_4_n293 ) );
INV_X4 _add_3_root_add_136_4_U370  ( .A(n14431), .ZN(_add_3_root_add_136_4_n294 ) );
XNOR2_X2 _add_3_root_add_136_4_U369  ( .A(_add_3_root_add_136_4_n291 ), .B(_add_3_root_add_136_4_n292 ), .ZN(N82) );
NAND2_X2 _add_3_root_add_136_4_U368  ( .A1(_add_3_root_add_136_4_n288 ),.A2(_add_3_root_add_136_4_n289 ), .ZN(_add_3_root_add_136_4_n278 ) );
NAND2_X2 _add_3_root_add_136_4_U367  ( .A1(_add_3_root_add_136_4_n78 ), .A2(_add_3_root_add_136_4_n241 ), .ZN(_add_3_root_add_136_4_n285 ) );
NAND2_X2 _add_3_root_add_136_4_U366  ( .A1(SHA1_ft_BCD[19]), .A2(n14428),.ZN(_add_3_root_add_136_4_n179 ) );
INV_X4 _add_3_root_add_136_4_U365  ( .A(SHA1_ft_BCD[19]), .ZN(_add_3_root_add_136_4_n283 ) );
INV_X4 _add_3_root_add_136_4_U364  ( .A(n14428), .ZN(_add_3_root_add_136_4_n284 ) );
NAND2_X2 _add_3_root_add_136_4_U363  ( .A1(_add_3_root_add_136_4_n283 ),.A2(_add_3_root_add_136_4_n284 ), .ZN(_add_3_root_add_136_4_n277 ) );
NAND2_X2 _add_3_root_add_136_4_U362  ( .A1(_add_3_root_add_136_4_n179 ),.A2(_add_3_root_add_136_4_n277 ), .ZN(_add_3_root_add_136_4_n282 ) );
XNOR2_X2 _add_3_root_add_136_4_U361  ( .A(_add_3_root_add_136_4_n281 ), .B(_add_3_root_add_136_4_n282 ), .ZN(N83) );
INV_X4 _add_3_root_add_136_4_U360  ( .A(_add_3_root_add_136_4_n280 ), .ZN(_add_3_root_add_136_4_n279 ) );
INV_X4 _add_3_root_add_136_4_U359  ( .A(_add_3_root_add_136_4_n179 ), .ZN(_add_3_root_add_136_4_n239 ) );
NAND2_X2 _add_3_root_add_136_4_U358  ( .A1(_add_3_root_add_136_4_n278 ),.A2(_add_3_root_add_136_4_n277 ), .ZN(_add_3_root_add_136_4_n192 ) );
INV_X4 _add_3_root_add_136_4_U357  ( .A(_add_3_root_add_136_4_n192 ), .ZN(_add_3_root_add_136_4_n240 ) );
INV_X4 _add_3_root_add_136_4_U356  ( .A(SHA1_ft_BCD[20]), .ZN(_add_3_root_add_136_4_n273 ) );
INV_X4 _add_3_root_add_136_4_U355  ( .A(n14425), .ZN(_add_3_root_add_136_4_n274 ) );
XNOR2_X2 _add_3_root_add_136_4_U354  ( .A(_add_3_root_add_136_4_n52 ), .B(_add_3_root_add_136_4_n272 ), .ZN(N84) );
INV_X4 _add_3_root_add_136_4_U353  ( .A(_add_3_root_add_136_4_n271 ), .ZN(_add_3_root_add_136_4_n265 ) );
INV_X4 _add_3_root_add_136_4_U352  ( .A(_add_3_root_add_136_4_n266 ), .ZN(_add_3_root_add_136_4_n270 ) );
XNOR2_X2 _add_3_root_add_136_4_U351  ( .A(_add_3_root_add_136_4_n267 ), .B(_add_3_root_add_136_4_n268 ), .ZN(N85) );
NOR2_X4 _add_3_root_add_136_4_U350  ( .A1(_add_3_root_add_136_4_n81 ), .A2(_add_3_root_add_136_4_n266 ), .ZN(_add_3_root_add_136_4_n252 ) );
NOR2_X4 _add_3_root_add_136_4_U349  ( .A1(_add_3_root_add_136_4_n81 ), .A2(_add_3_root_add_136_4_n265 ), .ZN(_add_3_root_add_136_4_n257 ) );
NAND2_X2 _add_3_root_add_136_4_U348  ( .A1(_add_3_root_add_136_4_n257 ),.A2(_add_3_root_add_136_4_n52 ), .ZN(_add_3_root_add_136_4_n263 ) );
NAND2_X2 _add_3_root_add_136_4_U347  ( .A1(SHA1_ft_BCD[22]), .A2(n14419),.ZN(_add_3_root_add_136_4_n254 ) );
INV_X4 _add_3_root_add_136_4_U346  ( .A(SHA1_ft_BCD[22]), .ZN(_add_3_root_add_136_4_n260 ) );
INV_X4 _add_3_root_add_136_4_U345  ( .A(n14419), .ZN(_add_3_root_add_136_4_n261 ) );
NAND2_X2 _add_3_root_add_136_4_U344  ( .A1(_add_3_root_add_136_4_n260 ),.A2(_add_3_root_add_136_4_n261 ), .ZN(_add_3_root_add_136_4_n255 ) );
NAND2_X2 _add_3_root_add_136_4_U343  ( .A1(_add_3_root_add_136_4_n254 ),.A2(_add_3_root_add_136_4_n255 ), .ZN(_add_3_root_add_136_4_n259 ) );
XNOR2_X2 _add_3_root_add_136_4_U342  ( .A(_add_3_root_add_136_4_n258 ), .B(_add_3_root_add_136_4_n259 ), .ZN(N86) );
NAND2_X2 _add_3_root_add_136_4_U341  ( .A1(_add_3_root_add_136_4_n257 ),.A2(_add_3_root_add_136_4_n255 ), .ZN(_add_3_root_add_136_4_n245 ) );
INV_X4 _add_3_root_add_136_4_U340  ( .A(_add_3_root_add_136_4_n255 ), .ZN(_add_3_root_add_136_4_n238 ) );
INV_X4 _add_3_root_add_136_4_U339  ( .A(_add_3_root_add_136_4_n254 ), .ZN(_add_3_root_add_136_4_n253 ) );
NOR3_X4 _add_3_root_add_136_4_U338  ( .A1(_add_3_root_add_136_4_n252 ), .A2(_add_3_root_add_136_4_n9 ), .A3(_add_3_root_add_136_4_n253 ), .ZN(_add_3_root_add_136_4_n236 ) );
NAND2_X2 _add_3_root_add_136_4_U337  ( .A1(SHA1_ft_BCD[23]), .A2(n14416),.ZN(_add_3_root_add_136_4_n235 ) );
INV_X4 _add_3_root_add_136_4_U336  ( .A(_add_3_root_add_136_4_n235 ), .ZN(_add_3_root_add_136_4_n173 ) );
INV_X4 _add_3_root_add_136_4_U335  ( .A(SHA1_ft_BCD[23]), .ZN(_add_3_root_add_136_4_n248 ) );
INV_X4 _add_3_root_add_136_4_U334  ( .A(n14416), .ZN(_add_3_root_add_136_4_n249 ) );
NAND2_X2 _add_3_root_add_136_4_U333  ( .A1(_add_3_root_add_136_4_n248 ),.A2(_add_3_root_add_136_4_n249 ), .ZN(_add_3_root_add_136_4_n244 ) );
INV_X4 _add_3_root_add_136_4_U332  ( .A(_add_3_root_add_136_4_n244 ), .ZN(_add_3_root_add_136_4_n237 ) );
XNOR2_X2 _add_3_root_add_136_4_U331  ( .A(_add_3_root_add_136_4_n246 ), .B(_add_3_root_add_136_4_n247 ), .ZN(N87) );
NAND2_X2 _add_3_root_add_136_4_U330  ( .A1(SHA1_ft_BCD[24]), .A2(n14413),.ZN(_add_3_root_add_136_4_n226 ) );
NOR2_X4 _add_3_root_add_136_4_U329  ( .A1(n14413), .A2(SHA1_ft_BCD[24]),.ZN(_add_3_root_add_136_4_n208 ) );
NAND2_X2 _add_3_root_add_136_4_U328  ( .A1(_add_3_root_add_136_4_n226 ),.A2(_add_3_root_add_136_4_n229 ), .ZN(_add_3_root_add_136_4_n232 ) );
INV_X4 _add_3_root_add_136_4_U327  ( .A(_add_3_root_add_136_4_n245 ), .ZN(_add_3_root_add_136_4_n243 ) );
INV_X4 _add_3_root_add_136_4_U326  ( .A(_add_3_root_add_136_4_n242 ), .ZN(_add_3_root_add_136_4_n134 ) );
INV_X4 _add_3_root_add_136_4_U325  ( .A(_add_3_root_add_136_4_n175 ), .ZN(_add_3_root_add_136_4_n234 ) );
NAND2_X2 _add_3_root_add_136_4_U324  ( .A1(_add_3_root_add_136_4_n233 ),.A2(_add_3_root_add_136_4_n230 ), .ZN(_add_3_root_add_136_4_n207 ) );
XNOR2_X2 _add_3_root_add_136_4_U323  ( .A(_add_3_root_add_136_4_n207 ), .B(_add_3_root_add_136_4_n232 ), .ZN(N88) );
NAND2_X2 _add_3_root_add_136_4_U322  ( .A1(_add_3_root_add_136_4_n230 ),.A2(_add_3_root_add_136_4_n233 ), .ZN(_add_3_root_add_136_4_n228 ) );
NAND2_X2 _add_3_root_add_136_4_U321  ( .A1(_add_3_root_add_136_4_n228 ),.A2(_add_3_root_add_136_4_n229 ), .ZN(_add_3_root_add_136_4_n227 ) );
NAND2_X2 _add_3_root_add_136_4_U320  ( .A1(SHA1_ft_BCD[25]), .A2(SHA1_result_148), .ZN(_add_3_root_add_136_4_n215 ) );
INV_X4 _add_3_root_add_136_4_U319  ( .A(SHA1_ft_BCD[25]), .ZN(_add_3_root_add_136_4_n224 ) );
INV_X4 _add_3_root_add_136_4_U318  ( .A(SHA1_result_148), .ZN(_add_3_root_add_136_4_n225 ) );
NAND2_X2 _add_3_root_add_136_4_U317  ( .A1(_add_3_root_add_136_4_n224 ),.A2(_add_3_root_add_136_4_n225 ), .ZN(_add_3_root_add_136_4_n221 ) );
NAND2_X2 _add_3_root_add_136_4_U316  ( .A1(_add_3_root_add_136_4_n215 ),.A2(_add_3_root_add_136_4_n221 ), .ZN(_add_3_root_add_136_4_n223 ) );
XNOR2_X2 _add_3_root_add_136_4_U315  ( .A(_add_3_root_add_136_4_n222 ), .B(_add_3_root_add_136_4_n223 ), .ZN(N89) );
INV_X4 _add_3_root_add_136_4_U314  ( .A(_add_3_root_add_136_4_n207 ), .ZN(_add_3_root_add_136_4_n201 ) );
INV_X4 _add_3_root_add_136_4_U313  ( .A(_add_3_root_add_136_4_n221 ), .ZN(_add_3_root_add_136_4_n210 ) );
NOR3_X4 _add_3_root_add_136_4_U312  ( .A1(_add_3_root_add_136_4_n201 ), .A2(_add_3_root_add_136_4_n210 ), .A3(_add_3_root_add_136_4_n208 ), .ZN(_add_3_root_add_136_4_n219 ) );
NAND2_X2 _add_3_root_add_136_4_U311  ( .A1(_add_3_root_add_136_4_n214 ),.A2(_add_3_root_add_136_4_n215 ), .ZN(_add_3_root_add_136_4_n220 ) );
NAND2_X2 _add_3_root_add_136_4_U310  ( .A1(SHA1_ft_BCD[26]), .A2(n14408),.ZN(_add_3_root_add_136_4_n200 ) );
INV_X4 _add_3_root_add_136_4_U309  ( .A(SHA1_ft_BCD[26]), .ZN(_add_3_root_add_136_4_n217 ) );
INV_X4 _add_3_root_add_136_4_U308  ( .A(n14408), .ZN(_add_3_root_add_136_4_n218 ) );
NAND2_X2 _add_3_root_add_136_4_U307  ( .A1(_add_3_root_add_136_4_n217 ),.A2(_add_3_root_add_136_4_n218 ), .ZN(_add_3_root_add_136_4_n211 ) );
XNOR2_X2 _add_3_root_add_136_4_U306  ( .A(_add_3_root_add_136_4_n216 ), .B(_add_3_root_add_136_4_n11 ), .ZN(N90) );
INV_X4 _add_3_root_add_136_4_U305  ( .A(_add_3_root_add_136_4_n200 ), .ZN(_add_3_root_add_136_4_n212 ) );
NAND2_X2 _add_3_root_add_136_4_U304  ( .A1(_add_3_root_add_136_4_n220 ),.A2(_add_3_root_add_136_4_n211 ), .ZN(_add_3_root_add_136_4_n199 ) );
INV_X4 _add_3_root_add_136_4_U303  ( .A(_add_3_root_add_136_4_n199 ), .ZN(_add_3_root_add_136_4_n213 ) );
INV_X4 _add_3_root_add_136_4_U302  ( .A(_add_3_root_add_136_4_n211 ), .ZN(_add_3_root_add_136_4_n209 ) );
NAND2_X2 _add_3_root_add_136_4_U301  ( .A1(_add_3_root_add_136_4_n202 ),.A2(_add_3_root_add_136_4_n207 ), .ZN(_add_3_root_add_136_4_n206 ) );
NAND2_X2 _add_3_root_add_136_4_U300  ( .A1(_add_3_root_add_136_4_n205 ),.A2(_add_3_root_add_136_4_n206 ), .ZN(_add_3_root_add_136_4_n203 ) );
NAND2_X2 _add_3_root_add_136_4_U299  ( .A1(SHA1_ft_BCD[27]), .A2(n14405),.ZN(_add_3_root_add_136_4_n196 ) );
NAND2_X2 _add_3_root_add_136_4_U298  ( .A1(_add_3_root_add_136_4_n196 ),.A2(_add_3_root_add_136_4_n198 ), .ZN(_add_3_root_add_136_4_n204 ) );
XNOR2_X2 _add_3_root_add_136_4_U297  ( .A(_add_3_root_add_136_4_n203 ), .B(_add_3_root_add_136_4_n204 ), .ZN(N91) );
NAND2_X2 _add_3_root_add_136_4_U296  ( .A1(_add_3_root_add_136_4_n202 ),.A2(_add_3_root_add_136_4_n198 ), .ZN(_add_3_root_add_136_4_n178 ) );
NAND2_X2 _add_3_root_add_136_4_U295  ( .A1(_add_3_root_add_136_4_n199 ),.A2(_add_3_root_add_136_4_n200 ), .ZN(_add_3_root_add_136_4_n197 ) );
NAND2_X2 _add_3_root_add_136_4_U294  ( .A1(_add_3_root_add_136_4_n197 ),.A2(_add_3_root_add_136_4_n198 ), .ZN(_add_3_root_add_136_4_n195 ) );
NAND2_X2 _add_3_root_add_136_4_U293  ( .A1(_add_3_root_add_136_4_n195 ),.A2(_add_3_root_add_136_4_n196 ), .ZN(_add_3_root_add_136_4_n171 ) );
NAND2_X2 _add_3_root_add_136_4_U292  ( .A1(SHA1_ft_BCD[28]), .A2(SHA1_result_151), .ZN(_add_3_root_add_136_4_n148 ) );
XNOR2_X2 _add_3_root_add_136_4_U291  ( .A(_add_3_root_add_136_4_n193 ), .B(_add_3_root_add_136_4_n17 ), .ZN(N92) );
INV_X4 _add_3_root_add_136_4_U290  ( .A(_add_3_root_add_136_4_n190 ), .ZN(_add_3_root_add_136_4_n187 ) );
NAND4_X2 _add_3_root_add_136_4_U289  ( .A1(_add_3_root_add_136_4_n182 ),.A2(_add_3_root_add_136_4_n32 ), .A3(_add_3_root_add_136_4_n184 ),.A4(_add_3_root_add_136_4_n185 ), .ZN(_add_3_root_add_136_4_n181 ) );
NAND2_X2 _add_3_root_add_136_4_U288  ( .A1(_add_3_root_add_136_4_n14 ), .A2(_add_3_root_add_136_4_n181 ), .ZN(_add_3_root_add_136_4_n180 ) );
INV_X4 _add_3_root_add_136_4_U287  ( .A(_add_3_root_add_136_4_n178 ), .ZN(_add_3_root_add_136_4_n177 ) );
NAND2_X2 _add_3_root_add_136_4_U286  ( .A1(_add_3_root_add_136_4_n177 ),.A2(_add_3_root_add_136_4_n172 ), .ZN(_add_3_root_add_136_4_n133 ) );
INV_X4 _add_3_root_add_136_4_U285  ( .A(_add_3_root_add_136_4_n133 ), .ZN(_add_3_root_add_136_4_n174 ) );
NAND2_X2 _add_3_root_add_136_4_U284  ( .A1(_add_3_root_add_136_4_n174 ),.A2(_add_3_root_add_136_4_n25 ), .ZN(_add_3_root_add_136_4_n176 ) );
NAND2_X2 _add_3_root_add_136_4_U283  ( .A1(_add_3_root_add_136_4_n36 ), .A2(_add_3_root_add_136_4_n174 ), .ZN(_add_3_root_add_136_4_n143 ) );
NAND2_X2 _add_3_root_add_136_4_U282  ( .A1(_add_3_root_add_136_4_n173 ),.A2(_add_3_root_add_136_4_n174 ), .ZN(_add_3_root_add_136_4_n144 ) );
NAND2_X2 _add_3_root_add_136_4_U281  ( .A1(_add_3_root_add_136_4_n143 ),.A2(_add_3_root_add_136_4_n144 ), .ZN(_add_3_root_add_136_4_n169 ) );
NAND2_X2 _add_3_root_add_136_4_U280  ( .A1(_add_3_root_add_136_4_n171 ),.A2(_add_3_root_add_136_4_n172 ), .ZN(_add_3_root_add_136_4_n159 ) );
NAND2_X2 _add_3_root_add_136_4_U279  ( .A1(_add_3_root_add_136_4_n159 ),.A2(_add_3_root_add_136_4_n148 ), .ZN(_add_3_root_add_136_4_n170 ) );
INV_X4 _add_3_root_add_136_4_U278  ( .A(_add_3_root_add_136_4_n156 ), .ZN(_add_3_root_add_136_4_n149 ) );
NAND2_X2 _add_3_root_add_136_4_U277  ( .A1(SHA1_ft_BCD[29]), .A2(n14400),.ZN(_add_3_root_add_136_4_n145 ) );
INV_X4 _add_3_root_add_136_4_U276  ( .A(_add_3_root_add_136_4_n145 ), .ZN(_add_3_root_add_136_4_n157 ) );
XNOR2_X2 _add_3_root_add_136_4_U275  ( .A(_add_3_root_add_136_4_n166 ), .B(_add_3_root_add_136_4_n167 ), .ZN(N93) );
INV_X4 _add_3_root_add_136_4_U274  ( .A(_add_3_root_add_136_4_n159 ), .ZN(_add_3_root_add_136_4_n146 ) );
NAND2_X2 _add_3_root_add_136_4_U273  ( .A1(_add_3_root_add_136_4_n146 ),.A2(_add_3_root_add_136_4_n156 ), .ZN(_add_3_root_add_136_4_n152 ) );
INV_X4 _add_3_root_add_136_4_U272  ( .A(_add_3_root_add_136_4_n131 ), .ZN(_add_3_root_add_136_4_n155 ) );
NAND4_X2 _add_3_root_add_136_4_U271  ( .A1(_add_3_root_add_136_4_n174 ),.A2(_add_3_root_add_136_4_n155 ), .A3(_add_3_root_add_136_4_n25 ),.A4(_add_3_root_add_136_4_n156 ), .ZN(_add_3_root_add_136_4_n154 ) );
NAND4_X2 _add_3_root_add_136_4_U270  ( .A1(_add_3_root_add_136_4_n151 ),.A2(_add_3_root_add_136_4_n152 ), .A3(_add_3_root_add_136_4_n153 ),.A4(_add_3_root_add_136_4_n154 ), .ZN(_add_3_root_add_136_4_n150 ) );
INV_X4 _add_3_root_add_136_4_U269  ( .A(_add_3_root_add_136_4_n135 ), .ZN(_add_3_root_add_136_4_n142 ) );
NAND2_X2 _add_3_root_add_136_4_U268  ( .A1(_add_3_root_add_136_4_n146 ),.A2(_add_3_root_add_136_4_n135 ), .ZN(_add_3_root_add_136_4_n137 ) );
NAND3_X2 _add_3_root_add_136_4_U267  ( .A1(_add_3_root_add_136_4_n136 ),.A2(_add_3_root_add_136_4_n137 ), .A3(_add_3_root_add_136_4_n138 ),.ZN(_add_3_root_add_136_4_n129 ) );
NAND2_X2 _add_3_root_add_136_4_U266  ( .A1(_add_3_root_add_136_4_n25 ), .A2(_add_3_root_add_136_4_n135 ), .ZN(_add_3_root_add_136_4_n132 ) );
XNOR2_X2 _add_3_root_add_136_4_U265  ( .A(_add_3_root_add_136_4_n127 ), .B(_add_3_root_add_136_4_n128 ), .ZN(N95) );
NOR2_X4 _add_3_root_add_136_4_U264  ( .A1(_add_3_root_add_136_4_n120 ), .A2(_add_3_root_add_136_4_n121 ), .ZN(_add_3_root_add_136_4_n119 ) );
INV_X4 _add_3_root_add_136_4_U263  ( .A(_add_3_root_add_136_4_n117 ), .ZN(_add_3_root_add_136_4_n116 ) );
XNOR2_X2 _add_3_root_add_136_4_U262  ( .A(_add_3_root_add_136_4_n103 ), .B(_add_3_root_add_136_4_n16 ), .ZN(N72) );
INV_X4 _add_3_root_add_136_4_U261  ( .A(_add_3_root_add_136_4_n96 ), .ZN(_add_3_root_add_136_4_n94 ) );
NAND2_X4 _add_3_root_add_136_4_U260  ( .A1(_add_3_root_add_136_4_n394 ),.A2(_add_3_root_add_136_4_n395 ), .ZN(_add_3_root_add_136_4_n310 ) );
NAND2_X4 _add_3_root_add_136_4_U259  ( .A1(_add_3_root_add_136_4_n310 ),.A2(_add_3_root_add_136_4_n108 ), .ZN(_add_3_root_add_136_4_n365 ) );
NAND2_X4 _add_3_root_add_136_4_U258  ( .A1(_add_3_root_add_136_4_n326 ),.A2(_add_3_root_add_136_4_n327 ), .ZN(_add_3_root_add_136_4_n351 ) );
NOR3_X2 _add_3_root_add_136_4_U257  ( .A1(_add_3_root_add_136_4_n342 ), .A2(_add_3_root_add_136_4_n348 ), .A3(_add_3_root_add_136_4_n70 ), .ZN(_add_3_root_add_136_4_n346 ) );
NAND3_X2 _add_3_root_add_136_4_U256  ( .A1(_add_3_root_add_136_4_n310 ),.A2(_add_3_root_add_136_4_n108 ), .A3(_add_3_root_add_136_4_n311 ),.ZN(_add_3_root_add_136_4_n185 ) );
NAND2_X4 _add_3_root_add_136_4_U255  ( .A1(_add_3_root_add_136_4_n110 ),.A2(_add_3_root_add_136_4_n38 ), .ZN(_add_3_root_add_136_4_n106 ) );
NAND2_X4 _add_3_root_add_136_4_U254  ( .A1(_add_3_root_add_136_4_n359 ),.A2(_add_3_root_add_136_4_n360 ), .ZN(_add_3_root_add_136_4_n358 ) );
NAND2_X4 _add_3_root_add_136_4_U253  ( .A1(_add_3_root_add_136_4_n382 ),.A2(_add_3_root_add_136_4_n383 ), .ZN(_add_3_root_add_136_4_n380 ) );
NAND2_X4 _add_3_root_add_136_4_U252  ( .A1(SHA1_ft_BCD[4]), .A2(n14464),.ZN(_add_3_root_add_136_4_n114 ) );
NAND2_X4 _add_3_root_add_136_4_U251  ( .A1(_add_3_root_add_136_4_n353 ),.A2(_add_3_root_add_136_4_n354 ), .ZN(_add_3_root_add_136_4_n328 ) );
NAND2_X1 _add_3_root_add_136_4_U250  ( .A1(_add_3_root_add_136_4_n328 ),.A2(_add_3_root_add_136_4_n329 ), .ZN(_add_3_root_add_136_4_n348 ) );
NOR3_X2 _add_3_root_add_136_4_U249  ( .A1(_add_3_root_add_136_4_n342 ), .A2(_add_3_root_add_136_4_n70 ), .A3(_add_3_root_add_136_4_n343 ), .ZN(_add_3_root_add_136_4_n337 ) );
NAND2_X4 _add_3_root_add_136_4_U248  ( .A1(_add_3_root_add_136_4_n368 ),.A2(_add_3_root_add_136_4_n369 ), .ZN(_add_3_root_add_136_4_n327 ) );
NOR2_X2 _add_3_root_add_136_4_U247  ( .A1(_add_3_root_add_136_4_n101 ), .A2(_add_3_root_add_136_4_n102 ), .ZN(_add_3_root_add_136_4_n99 ) );
INV_X4 _add_3_root_add_136_4_U246  ( .A(_add_3_root_add_136_4_n279 ), .ZN(_add_3_root_add_136_4_n163 ) );
INV_X4 _add_3_root_add_136_4_U245  ( .A(_add_3_root_add_136_4_n37 ), .ZN(_add_3_root_add_136_4_n184 ) );
AND2_X2 _add_3_root_add_136_4_U244  ( .A1(SHA1_ft_BCD[15]), .A2(n14440),.ZN(_add_3_root_add_136_4_n85 ) );
AND2_X2 _add_3_root_add_136_4_U243  ( .A1(SHA1_ft_BCD[30]), .A2(n14397),.ZN(_add_3_root_add_136_4_n84 ) );
NOR2_X4 _add_3_root_add_136_4_U242  ( .A1(SHA1_ft_BCD[21]), .A2(n14422),.ZN(_add_3_root_add_136_4_n81 ) );
NOR2_X2 _add_3_root_add_136_4_U241  ( .A1(SHA1_ft_BCD[30]), .A2(n14397),.ZN(_add_3_root_add_136_4_n80 ) );
OR2_X2 _add_3_root_add_136_4_U240  ( .A1(SHA1_ft_BCD[28]), .A2(SHA1_result_151), .ZN(_add_3_root_add_136_4_n172 ) );
OR2_X2 _add_3_root_add_136_4_U239  ( .A1(SHA1_ft_BCD[27]), .A2(n14405), .ZN(_add_3_root_add_136_4_n198 ) );
NAND2_X2 _add_3_root_add_136_4_U238  ( .A1(n14930), .A2(SHA1_result_128),.ZN(_add_3_root_add_136_4_n115 ) );
XOR2_X2 _add_3_root_add_136_4_U237  ( .A(n14394), .B(SHA1_ft_BCD[31]), .Z(_add_3_root_add_136_4_n128 ) );
OR2_X2 _add_3_root_add_136_4_U236  ( .A1(SHA1_ft_BCD[29]), .A2(n14400), .ZN(_add_3_root_add_136_4_n156 ) );
NOR2_X4 _add_3_root_add_136_4_U235  ( .A1(SHA1_ft_BCD[14]), .A2(n14443),.ZN(_add_3_root_add_136_4_n79 ) );
INV_X4 _add_3_root_add_136_4_U234  ( .A(_add_3_root_add_136_4_n380 ), .ZN(_add_3_root_add_136_4_n123 ) );
NOR2_X1 _add_3_root_add_136_4_U233  ( .A1(_add_3_root_add_136_4_n149 ), .A2(_add_3_root_add_136_4_n148 ), .ZN(_add_3_root_add_136_4_n158 ) );
NOR2_X2 _add_3_root_add_136_4_U232  ( .A1(_add_3_root_add_136_4_n157 ), .A2(_add_3_root_add_136_4_n158 ), .ZN(_add_3_root_add_136_4_n153 ) );
AND2_X2 _add_3_root_add_136_4_U231  ( .A1(_add_3_root_add_136_4_n347 ), .A2(_add_3_root_add_136_4_n329 ), .ZN(_add_3_root_add_136_4_n76 ) );
NOR2_X1 _add_3_root_add_136_4_U230  ( .A1(_add_3_root_add_136_4_n142 ), .A2(_add_3_root_add_136_4_n148 ), .ZN(_add_3_root_add_136_4_n147 ) );
NOR2_X1 _add_3_root_add_136_4_U229  ( .A1(_add_3_root_add_136_4_n79 ), .A2(_add_3_root_add_136_4_n28 ), .ZN(_add_3_root_add_136_4_n341 ) );
NOR2_X2 _add_3_root_add_136_4_U228  ( .A1(_add_3_root_add_136_4_n296 ), .A2(_add_3_root_add_136_4_n297 ), .ZN(_add_3_root_add_136_4_n286 ) );
NOR3_X1 _add_3_root_add_136_4_U227  ( .A1(_add_3_root_add_136_4_n208 ), .A2(_add_3_root_add_136_4_n209 ), .A3(_add_3_root_add_136_4_n210 ), .ZN(_add_3_root_add_136_4_n202 ) );
NOR2_X1 _add_3_root_add_136_4_U226  ( .A1(_add_3_root_add_136_4_n324 ), .A2(_add_3_root_add_136_4_n79 ), .ZN(_add_3_root_add_136_4_n345 ) );
NOR2_X2 _add_3_root_add_136_4_U225  ( .A1(_add_3_root_add_136_4_n84 ), .A2(_add_3_root_add_136_4_n147 ), .ZN(_add_3_root_add_136_4_n136 ) );
AND2_X2 _add_3_root_add_136_4_U224  ( .A1(_add_3_root_add_136_4_n192 ), .A2(_add_3_root_add_136_4_n72 ), .ZN(_add_3_root_add_136_4_n131 ) );
NOR2_X1 _add_3_root_add_136_4_U223  ( .A1(_add_3_root_add_136_4_n81 ), .A2(_add_3_root_add_136_4_n9 ), .ZN(_add_3_root_add_136_4_n268 ) );
NOR3_X2 _add_3_root_add_136_4_U222  ( .A1(_add_3_root_add_136_4_n168 ), .A2(_add_3_root_add_136_4_n169 ), .A3(_add_3_root_add_136_4_n170 ), .ZN(_add_3_root_add_136_4_n166 ) );
NOR2_X2 _add_3_root_add_136_4_U221  ( .A1(_add_3_root_add_136_4_n149 ), .A2(_add_3_root_add_136_4_n157 ), .ZN(_add_3_root_add_136_4_n167 ) );
NOR2_X2 _add_3_root_add_136_4_U220  ( .A1(_add_3_root_add_136_4_n194 ), .A2(_add_3_root_add_136_4_n171 ), .ZN(_add_3_root_add_136_4_n193 ) );
NOR2_X2 _add_3_root_add_136_4_U219  ( .A1(_add_3_root_add_136_4_n212 ), .A2(_add_3_root_add_136_4_n213 ), .ZN(_add_3_root_add_136_4_n205 ) );
NOR2_X1 _add_3_root_add_136_4_U218  ( .A1(_add_3_root_add_136_4_n9 ), .A2(_add_3_root_add_136_4_n252 ), .ZN(_add_3_root_add_136_4_n262 ) );
NOR2_X1 _add_3_root_add_136_4_U217  ( .A1(_add_3_root_add_136_4_n331 ), .A2(_add_3_root_add_136_4_n85 ), .ZN(_add_3_root_add_136_4_n334 ) );
INV_X8 _add_3_root_add_136_4_U216  ( .A(_add_3_root_add_136_4_n86 ), .ZN(_add_3_root_add_136_4_n87 ) );
NOR2_X1 _add_3_root_add_136_4_U215  ( .A1(_add_3_root_add_136_4_n149 ), .A2(_add_3_root_add_136_4_n144 ), .ZN(_add_3_root_add_136_4_n161 ) );
NOR2_X1 _add_3_root_add_136_4_U214  ( .A1(_add_3_root_add_136_4_n149 ), .A2(_add_3_root_add_136_4_n143 ), .ZN(_add_3_root_add_136_4_n160 ) );
NOR2_X2 _add_3_root_add_136_4_U213  ( .A1(_add_3_root_add_136_4_n160 ), .A2(_add_3_root_add_136_4_n161 ), .ZN(_add_3_root_add_136_4_n151 ) );
INV_X2 _add_3_root_add_136_4_U212  ( .A(_add_3_root_add_136_4_n102 ), .ZN(_add_3_root_add_136_4_n189 ) );
NAND3_X1 _add_3_root_add_136_4_U211  ( .A1(_add_3_root_add_136_4_n14 ), .A2(_add_3_root_add_136_4_n134 ), .A3(_add_3_root_add_136_4_n241 ), .ZN(_add_3_root_add_136_4_n230 ) );
NOR2_X1 _add_3_root_add_136_4_U210  ( .A1(_add_3_root_add_136_4_n256 ), .A2(_add_3_root_add_136_4_n245 ), .ZN(_add_3_root_add_136_4_n250 ) );
NOR2_X1 _add_3_root_add_136_4_U209  ( .A1(_add_3_root_add_136_4_n201 ), .A2(_add_3_root_add_136_4_n178 ), .ZN(_add_3_root_add_136_4_n194 ) );
AND2_X2 _add_3_root_add_136_4_U208  ( .A1(_add_3_root_add_136_4_n240 ), .A2(_add_3_root_add_136_4_n134 ), .ZN(_add_3_root_add_136_4_n68 ) );
NOR2_X2 _add_3_root_add_136_4_U207  ( .A1(_add_3_root_add_136_4_n131 ), .A2(_add_3_root_add_136_4_n176 ), .ZN(_add_3_root_add_136_4_n168 ) );
NOR3_X1 _add_3_root_add_136_4_U206  ( .A1(_add_3_root_add_136_4_n131 ), .A2(_add_3_root_add_136_4_n132 ), .A3(_add_3_root_add_136_4_n133 ), .ZN(_add_3_root_add_136_4_n130 ) );
NOR2_X1 _add_3_root_add_136_4_U205  ( .A1(_add_3_root_add_136_4_n142 ), .A2(_add_3_root_add_136_4_n143 ), .ZN(_add_3_root_add_136_4_n141 ) );
NOR2_X1 _add_3_root_add_136_4_U204  ( .A1(_add_3_root_add_136_4_n142 ), .A2(_add_3_root_add_136_4_n144 ), .ZN(_add_3_root_add_136_4_n140 ) );
NAND2_X2 _add_3_root_add_136_4_U203  ( .A1(_add_3_root_add_136_4_n327 ),.A2(_add_3_root_add_136_4_n326 ), .ZN(_add_3_root_add_136_4_n67 ) );
NOR2_X2 _add_3_root_add_136_4_U202  ( .A1(_add_3_root_add_136_4_n129 ), .A2(_add_3_root_add_136_4_n130 ), .ZN(_add_3_root_add_136_4_n127 ) );
INV_X1 _add_3_root_add_136_4_U201  ( .A(n14391), .ZN(_add_3_root_add_136_4_n403 ) );
OR2_X4 _add_3_root_add_136_4_U200  ( .A1(SHA1_ft_BCD[7]), .A2(SHA1_result_130), .ZN(_add_3_root_add_136_4_n108 ) );
AND2_X2 _add_3_root_add_136_4_U199  ( .A1(_add_3_root_add_136_4_n179 ), .A2(_add_3_root_add_136_4_n180 ), .ZN(_add_3_root_add_136_4_n72 ) );
NOR2_X1 _add_3_root_add_136_4_U198  ( .A1(_add_3_root_add_136_4_n80 ), .A2(_add_3_root_add_136_4_n145 ), .ZN(_add_3_root_add_136_4_n139 ) );
NOR3_X1 _add_3_root_add_136_4_U197  ( .A1(_add_3_root_add_136_4_n139 ), .A2(_add_3_root_add_136_4_n140 ), .A3(_add_3_root_add_136_4_n141 ), .ZN(_add_3_root_add_136_4_n138 ) );
NOR2_X2 _add_3_root_add_136_4_U196  ( .A1(_add_3_root_add_136_4_n80 ), .A2(_add_3_root_add_136_4_n84 ), .ZN(_add_3_root_add_136_4_n66 ) );
XOR2_X2 _add_3_root_add_136_4_U195  ( .A(_add_3_root_add_136_4_n150 ), .B(_add_3_root_add_136_4_n66 ), .Z(N94) );
NOR2_X1 _add_3_root_add_136_4_U194  ( .A1(_add_3_root_add_136_4_n80 ), .A2(_add_3_root_add_136_4_n149 ), .ZN(_add_3_root_add_136_4_n135 ) );
NOR2_X1 _add_3_root_add_136_4_U193  ( .A1(_add_3_root_add_136_4_n30 ), .A2(_add_3_root_add_136_4_n21 ), .ZN(_add_3_root_add_136_4_n64 ) );
NOR2_X1 _add_3_root_add_136_4_U192  ( .A1(_add_3_root_add_136_4_n105 ), .A2(_add_3_root_add_136_4_n100 ), .ZN(_add_3_root_add_136_4_n363 ) );
INV_X1 _add_3_root_add_136_4_U191  ( .A(_add_3_root_add_136_4_n316 ), .ZN(_add_3_root_add_136_4_n314 ) );
NOR2_X2 _add_3_root_add_136_4_U190  ( .A1(_add_3_root_add_136_4_n10 ), .A2(_add_3_root_add_136_4_n317 ), .ZN(_add_3_root_add_136_4_n312 ) );
NOR2_X2 _add_3_root_add_136_4_U189  ( .A1(_add_3_root_add_136_4_n250 ), .A2(_add_3_root_add_136_4_n251 ), .ZN(_add_3_root_add_136_4_n246 ) );
NOR2_X1 _add_3_root_add_136_4_U188  ( .A1(_add_3_root_add_136_4_n238 ), .A2(_add_3_root_add_136_4_n236 ), .ZN(_add_3_root_add_136_4_n251 ) );
NAND3_X2 _add_3_root_add_136_4_U187  ( .A1(n14437), .A2(SHA1_ft_BCD[16]),.A3(_add_3_root_add_136_4_n298 ), .ZN(_add_3_root_add_136_4_n299 ) );
NAND3_X1 _add_3_root_add_136_4_U186  ( .A1(n14413), .A2(SHA1_ft_BCD[24]),.A3(_add_3_root_add_136_4_n221 ), .ZN(_add_3_root_add_136_4_n214 ) );
INV_X8 _add_3_root_add_136_4_U185  ( .A(_add_3_root_add_136_4_n365 ), .ZN(_add_3_root_add_136_4_n100 ) );
NAND2_X4 _add_3_root_add_136_4_U184  ( .A1(_add_3_root_add_136_4_n62 ), .A2(_add_3_root_add_136_4_n63 ), .ZN(N74) );
NAND2_X4 _add_3_root_add_136_4_U183  ( .A1(_add_3_root_add_136_4_n60 ), .A2(_add_3_root_add_136_4_n61 ), .ZN(_add_3_root_add_136_4_n63 ) );
NAND2_X2 _add_3_root_add_136_4_U182  ( .A1(_add_3_root_add_136_4_n371 ),.A2(_add_3_root_add_136_4_n372 ), .ZN(_add_3_root_add_136_4_n62 ) );
INV_X2 _add_3_root_add_136_4_U181  ( .A(_add_3_root_add_136_4_n372 ), .ZN(_add_3_root_add_136_4_n60 ) );
NAND2_X4 _add_3_root_add_136_4_U180  ( .A1(_add_3_root_add_136_4_n58 ), .A2(_add_3_root_add_136_4_n59 ), .ZN(N70) );
NOR2_X4 _add_3_root_add_136_4_U179  ( .A1(_add_3_root_add_136_4_n18 ), .A2(_add_3_root_add_136_4_n361 ), .ZN(_add_3_root_add_136_4_n359 ) );
INV_X2 _add_3_root_add_136_4_U178  ( .A(_add_3_root_add_136_4_n64 ), .ZN(_add_3_root_add_136_4_n57 ) );
NAND2_X1 _add_3_root_add_136_4_U177  ( .A1(_add_3_root_add_136_4_n108 ),.A2(_add_3_root_add_136_4_n8 ), .ZN(_add_3_root_add_136_4_n107 ) );
INV_X4 _add_3_root_add_136_4_U176  ( .A(_add_3_root_add_136_4_n106 ), .ZN(_add_3_root_add_136_4_n53 ) );
NAND2_X4 _add_3_root_add_136_4_U175  ( .A1(_add_3_root_add_136_4_n56 ), .A2(_add_3_root_add_136_4_n55 ), .ZN(N71) );
NAND2_X4 _add_3_root_add_136_4_U174  ( .A1(_add_3_root_add_136_4_n53 ), .A2(_add_3_root_add_136_4_n54 ), .ZN(_add_3_root_add_136_4_n56 ) );
NAND2_X4 _add_3_root_add_136_4_U173  ( .A1(SHA1_ft_BCD[0]), .A2(n14391),.ZN(_add_3_root_add_136_4_n280 ) );
AND2_X2 _add_3_root_add_136_4_U172  ( .A1(_add_3_root_add_136_4_n379 ), .A2(_add_3_root_add_136_4_n163 ), .ZN(N64) );
INV_X2 _add_3_root_add_136_4_U171  ( .A(_add_3_root_add_136_4_n107 ), .ZN(_add_3_root_add_136_4_n54 ) );
NAND2_X2 _add_3_root_add_136_4_U170  ( .A1(_add_3_root_add_136_4_n275 ),.A2(_add_3_root_add_136_4_n276 ), .ZN(_add_3_root_add_136_4_n52 ) );
INV_X8 _add_3_root_add_136_4_U169  ( .A(_add_3_root_add_136_4_n6 ), .ZN(N77));
INV_X1 _add_3_root_add_136_4_U168  ( .A(_add_3_root_add_136_4_n41 ), .ZN(_add_3_root_add_136_4_n402 ) );
NAND2_X4 _add_3_root_add_136_4_U167  ( .A1(_add_3_root_add_136_4_n398 ),.A2(_add_3_root_add_136_4_n399 ), .ZN(_add_3_root_add_136_4_n112 ) );
NAND2_X4 _add_3_root_add_136_4_U166  ( .A1(_add_3_root_add_136_4_n293 ),.A2(_add_3_root_add_136_4_n294 ), .ZN(_add_3_root_add_136_4_n287 ) );
INV_X1 _add_3_root_add_136_4_U165  ( .A(_add_3_root_add_136_4_n328 ), .ZN(_add_3_root_add_136_4_n350 ) );
NAND2_X1 _add_3_root_add_136_4_U164  ( .A1(_add_3_root_add_136_4_n341 ),.A2(_add_3_root_add_136_4_n328 ), .ZN(_add_3_root_add_136_4_n343 ) );
NOR2_X4 _add_3_root_add_136_4_U163  ( .A1(_add_3_root_add_136_4_n239 ), .A2(_add_3_root_add_136_4_n240 ), .ZN(_add_3_root_add_136_4_n275 ) );
NAND2_X4 _add_3_root_add_136_4_U162  ( .A1(_add_3_root_add_136_4_n303 ),.A2(_add_3_root_add_136_4_n304 ), .ZN(_add_3_root_add_136_4_n298 ) );
NAND2_X1 _add_3_root_add_136_4_U161  ( .A1(_add_3_root_add_136_4_n298 ),.A2(_add_3_root_add_136_4_n300 ), .ZN(_add_3_root_add_136_4_n302 ) );
INV_X1 _add_3_root_add_136_4_U160  ( .A(_add_3_root_add_136_4_n298 ), .ZN(_add_3_root_add_136_4_n296 ) );
NAND2_X4 _add_3_root_add_136_4_U159  ( .A1(SHA1_ft_BCD[7]), .A2(SHA1_result_130), .ZN(_add_3_root_add_136_4_n109 ) );
NAND2_X4 _add_3_root_add_136_4_U158  ( .A1(_add_3_root_add_136_4_n273 ),.A2(_add_3_root_add_136_4_n274 ), .ZN(_add_3_root_add_136_4_n271 ) );
NAND2_X1 _add_3_root_add_136_4_U157  ( .A1(_add_3_root_add_136_4_n271 ),.A2(_add_3_root_add_136_4_n266 ), .ZN(_add_3_root_add_136_4_n272 ) );
NOR2_X4 _add_3_root_add_136_4_U156  ( .A1(_add_3_root_add_136_4_n269 ), .A2(_add_3_root_add_136_4_n270 ), .ZN(_add_3_root_add_136_4_n267 ) );
NAND2_X4 _add_3_root_add_136_4_U155  ( .A1(_add_3_root_add_136_4_n263 ),.A2(_add_3_root_add_136_4_n262 ), .ZN(_add_3_root_add_136_4_n258 ) );
NOR2_X1 _add_3_root_add_136_4_U154  ( .A1(_add_3_root_add_136_4_n10 ), .A2(_add_3_root_add_136_4_n123 ), .ZN(_add_3_root_add_136_4_n50 ) );
XNOR2_X2 _add_3_root_add_136_4_U153  ( .A(_add_3_root_add_136_4_n122 ), .B(_add_3_root_add_136_4_n50 ), .ZN(N67) );
NAND2_X2 _add_3_root_add_136_4_U152  ( .A1(_add_3_root_add_136_4_n357 ),.A2(_add_3_root_add_136_4_n362 ), .ZN(_add_3_root_add_136_4_n372 ) );
NAND2_X2 _add_3_root_add_136_4_U151  ( .A1(_add_3_root_add_136_4_n371 ),.A2(_add_3_root_add_136_4_n362 ), .ZN(_add_3_root_add_136_4_n370 ) );
NAND3_X4 _add_3_root_add_136_4_U150  ( .A1(_add_3_root_add_136_4_n327 ),.A2(_add_3_root_add_136_4_n362 ), .A3(_add_3_root_add_136_4_n364 ),.ZN(_add_3_root_add_136_4_n191 ) );
NOR2_X4 _add_3_root_add_136_4_U149  ( .A1(_add_3_root_add_136_4_n388 ), .A2(_add_3_root_add_136_4_n389 ), .ZN(_add_3_root_add_136_4_n373 ) );
NOR2_X2 _add_3_root_add_136_4_U148  ( .A1(_add_3_root_add_136_4_n365 ), .A2(_add_3_root_add_136_4_n19 ), .ZN(_add_3_root_add_136_4_n388 ) );
NAND2_X4 _add_3_root_add_136_4_U147  ( .A1(_add_3_root_add_136_4_n384 ),.A2(_add_3_root_add_136_4_n385 ), .ZN(_add_3_root_add_136_4_n378 ) );
NOR2_X4 _add_3_root_add_136_4_U146  ( .A1(_add_3_root_add_136_4_n99 ), .A2(_add_3_root_add_136_4_n100 ), .ZN(_add_3_root_add_136_4_n97 ) );
AND2_X2 _add_3_root_add_136_4_U145  ( .A1(_add_3_root_add_136_4_n114 ), .A2(_add_3_root_add_136_4_n115 ), .ZN(_add_3_root_add_136_4_n48 ) );
INV_X1 _add_3_root_add_136_4_U144  ( .A(_add_3_root_add_136_4_n115 ), .ZN(_add_3_root_add_136_4_n47 ) );
OR2_X1 _add_3_root_add_136_4_U143  ( .A1(_add_3_root_add_136_4_n47 ), .A2(_add_3_root_add_136_4_n112 ), .ZN(_add_3_root_add_136_4_n46 ) );
NAND2_X2 _add_3_root_add_136_4_U142  ( .A1(_add_3_root_add_136_4_n116 ),.A2(_add_3_root_add_136_4_n48 ), .ZN(_add_3_root_add_136_4_n45 ) );
NAND3_X2 _add_3_root_add_136_4_U141  ( .A1(_add_3_root_add_136_4_n358 ),.A2(_add_3_root_add_136_4_n357 ), .A3(_add_3_root_add_136_4_n356 ),.ZN(_add_3_root_add_136_4_n326 ) );
INV_X4 _add_3_root_add_136_4_U140  ( .A(_add_3_root_add_136_4_n71 ), .ZN(N66) );
INV_X4 _add_3_root_add_136_4_U139  ( .A(_add_3_root_add_136_4_n44 ), .ZN(_add_3_root_add_136_4_n118 ) );
NAND2_X4 _add_3_root_add_136_4_U138  ( .A1(_add_3_root_add_136_4_n45 ), .A2(_add_3_root_add_136_4_n46 ), .ZN(_add_3_root_add_136_4_n44 ) );
NAND2_X4 _add_3_root_add_136_4_U137  ( .A1(_add_3_root_add_136_4_n397 ),.A2(_add_3_root_add_136_4_n396 ), .ZN(_add_3_root_add_136_4_n395 ) );
INV_X4 _add_3_root_add_136_4_U136  ( .A(_add_3_root_add_136_4_n191 ), .ZN(_add_3_root_add_136_4_n186 ) );
NOR2_X2 _add_3_root_add_136_4_U135  ( .A1(_add_3_root_add_136_4_n331 ), .A2(_add_3_root_add_136_4_n79 ), .ZN(_add_3_root_add_136_4_n330 ) );
NAND3_X4 _add_3_root_add_136_4_U134  ( .A1(_add_3_root_add_136_4_n330 ),.A2(_add_3_root_add_136_4_n329 ), .A3(_add_3_root_add_136_4_n328 ),.ZN(_add_3_root_add_136_4_n190 ) );
NAND2_X4 _add_3_root_add_136_4_U133  ( .A1(SHA1_ft_BCD[9]), .A2(SHA1_result_132), .ZN(_add_3_root_add_136_4_n93 ) );
INV_X8 _add_3_root_add_136_4_U132  ( .A(_add_3_root_add_136_4_n87 ), .ZN(_add_3_root_add_136_4_n376 ) );
OR2_X1 _add_3_root_add_136_4_U131  ( .A1(_add_3_root_add_136_4_n121 ), .A2(_add_3_root_add_136_4_n83 ), .ZN(_add_3_root_add_136_4_n43 ) );
XNOR2_X2 _add_3_root_add_136_4_U130  ( .A(_add_3_root_add_136_4_n376 ), .B(_add_3_root_add_136_4_n43 ), .ZN(N68) );
OR2_X2 _add_3_root_add_136_4_U129  ( .A1(_add_3_root_add_136_4_n125 ), .A2(_add_3_root_add_136_4_n15 ), .ZN(_add_3_root_add_136_4_n42 ) );
XNOR2_X1 _add_3_root_add_136_4_U128  ( .A(_add_3_root_add_136_4_n126 ), .B(_add_3_root_add_136_4_n42 ), .ZN(_add_3_root_add_136_4_n71 ) );
INV_X2 _add_3_root_add_136_4_U127  ( .A(_add_3_root_add_136_4_n162 ), .ZN(_add_3_root_add_136_4_n125 ) );
BUF_X16 _add_3_root_add_136_4_U126  ( .A(SHA1_ft_BCD[0]), .Z(_add_3_root_add_136_4_n41 ) );
NAND3_X2 _add_3_root_add_136_4_U125  ( .A1(_add_3_root_add_136_4_n116 ),.A2(_add_3_root_add_136_4_n115 ), .A3(_add_3_root_add_136_4_n39 ),.ZN(_add_3_root_add_136_4_n113 ) );
OR2_X4 _add_3_root_add_136_4_U124  ( .A1(_add_3_root_add_136_4_n273 ), .A2(_add_3_root_add_136_4_n274 ), .ZN(_add_3_root_add_136_4_n266 ) );
NAND2_X4 _add_3_root_add_136_4_U123  ( .A1(SHA1_ft_BCD[8]), .A2(SHA1_result_131), .ZN(_add_3_root_add_136_4_n95 ) );
NAND2_X2 _add_3_root_add_136_4_U122  ( .A1(_add_3_root_add_136_4_n370 ),.A2(_add_3_root_add_136_4_n357 ), .ZN(_add_3_root_add_136_4_n366 ) );
NOR2_X4 _add_3_root_add_136_4_U121  ( .A1(n14929), .A2(n14388), .ZN(_add_3_root_add_136_4_n90 ) );
INV_X8 _add_3_root_add_136_4_U120  ( .A(_add_3_root_add_136_4_n90 ), .ZN(_add_3_root_add_136_4_n164 ) );
INV_X8 _add_3_root_add_136_4_U119  ( .A(_add_3_root_add_136_4_n351 ), .ZN(_add_3_root_add_136_4_n352 ) );
NOR2_X4 _add_3_root_add_136_4_U118  ( .A1(_add_3_root_add_136_4_n352 ), .A2(_add_3_root_add_136_4_n186 ), .ZN(_add_3_root_add_136_4_n70 ) );
NOR2_X4 _add_3_root_add_136_4_U117  ( .A1(_add_3_root_add_136_4_n219 ), .A2(_add_3_root_add_136_4_n220 ), .ZN(_add_3_root_add_136_4_n216 ) );
NAND2_X4 _add_3_root_add_136_4_U116  ( .A1(_add_3_root_add_136_4_n234 ),.A2(_add_3_root_add_136_4_n235 ), .ZN(_add_3_root_add_136_4_n231 ) );
AND2_X2 _add_3_root_add_136_4_U115  ( .A1(_add_3_root_add_136_4_n239 ), .A2(_add_3_root_add_136_4_n134 ), .ZN(_add_3_root_add_136_4_n69 ) );
NOR3_X4 _add_3_root_add_136_4_U114  ( .A1(_add_3_root_add_136_4_n68 ), .A2(_add_3_root_add_136_4_n69 ), .A3(_add_3_root_add_136_4_n231 ), .ZN(_add_3_root_add_136_4_n233 ) );
BUF_X16 _add_3_root_add_136_4_U113  ( .A(_add_3_root_add_136_4_n114 ), .Z(_add_3_root_add_136_4_n39 ) );
NOR2_X4 _add_3_root_add_136_4_U112  ( .A1(_add_3_root_add_136_4_n346 ), .A2(_add_3_root_add_136_4_n76 ), .ZN(_add_3_root_add_136_4_n344 ) );
NAND2_X2 _add_3_root_add_136_4_U111  ( .A1(_add_3_root_add_136_4_n106 ),.A2(_add_3_root_add_136_4_n107 ), .ZN(_add_3_root_add_136_4_n55 ) );
NOR3_X4 _add_3_root_add_136_4_U110  ( .A1(_add_3_root_add_136_4_n236 ), .A2(_add_3_root_add_136_4_n237 ), .A3(_add_3_root_add_136_4_n238 ), .ZN(_add_3_root_add_136_4_n175 ) );
INV_X1 _add_3_root_add_136_4_U109  ( .A(_add_3_root_add_136_4_n234 ), .ZN(_add_3_root_add_136_4_n36 ) );
NAND2_X4 _add_3_root_add_136_4_U108  ( .A1(SHA1_ft_BCD[2]), .A2(n14385),.ZN(_add_3_root_add_136_4_n162 ) );
NOR2_X4 _add_3_root_add_136_4_U107  ( .A1(SHA1_ft_BCD[6]), .A2(SHA1_result_129), .ZN(_add_3_root_add_136_4_n35 ) );
INV_X2 _add_3_root_add_136_4_U106  ( .A(_add_3_root_add_136_4_n33 ), .ZN(_add_3_root_add_136_4_n34 ) );
INV_X1 _add_3_root_add_136_4_U105  ( .A(_add_3_root_add_136_4_n318 ), .ZN(_add_3_root_add_136_4_n32 ) );
INV_X2 _add_3_root_add_136_4_U104  ( .A(SHA1_ft_BCD[6]), .ZN(_add_3_root_add_136_4_n400 ) );
NAND2_X2 _add_3_root_add_136_4_U103  ( .A1(_add_3_root_add_136_4_n44 ), .A2(_add_3_root_add_136_4_n64 ), .ZN(_add_3_root_add_136_4_n59 ) );
NOR2_X4 _add_3_root_add_136_4_U102  ( .A1(_add_3_root_add_136_4_n190 ), .A2(_add_3_root_add_136_4_n191 ), .ZN(_add_3_root_add_136_4_n311 ) );
NAND2_X4 _add_3_root_add_136_4_U101  ( .A1(_add_3_root_add_136_4_n390 ),.A2(_add_3_root_add_136_4_n391 ), .ZN(_add_3_root_add_136_4_n92 ) );
INV_X1 _add_3_root_add_136_4_U100  ( .A(_add_3_root_add_136_4_n361 ), .ZN(_add_3_root_add_136_4_n29 ) );
XNOR2_X2 _add_3_root_add_136_4_U99  ( .A(_add_3_root_add_136_4_n65 ), .B(_add_3_root_add_136_4_n3 ), .ZN(N76) );
NAND2_X1 _add_3_root_add_136_4_U98  ( .A1(_add_3_root_add_136_4_n402 ), .A2(_add_3_root_add_136_4_n403 ), .ZN(_add_3_root_add_136_4_n379 ) );
INV_X4 _add_3_root_add_136_4_U97  ( .A(_add_3_root_add_136_4_n28 ), .ZN(_add_3_root_add_136_4_n329 ) );
NOR2_X4 _add_3_root_add_136_4_U96  ( .A1(SHA1_ft_BCD[13]), .A2(SHA1_result_136), .ZN(_add_3_root_add_136_4_n28 ) );
NAND2_X1 _add_3_root_add_136_4_U95  ( .A1(n14434), .A2(SHA1_ft_BCD[17]),.ZN(_add_3_root_add_136_4_n300 ) );
AND2_X2 _add_3_root_add_136_4_U94  ( .A1(_add_3_root_add_136_4_n299 ), .A2(_add_3_root_add_136_4_n300 ), .ZN(_add_3_root_add_136_4_n27 ) );
NAND2_X4 _add_3_root_add_136_4_U93  ( .A1(SHA1_ft_BCD[12]), .A2(SHA1_result_135), .ZN(_add_3_root_add_136_4_n322 ) );
NOR2_X4 _add_3_root_add_136_4_U92  ( .A1(_add_3_root_add_136_4_n124 ), .A2(_add_3_root_add_136_4_n125 ), .ZN(_add_3_root_add_136_4_n122 ) );
NOR2_X1 _add_3_root_add_136_4_U91  ( .A1(_add_3_root_add_136_4_n361 ), .A2(_add_3_root_add_136_4_n95 ), .ZN(_add_3_root_add_136_4_n389 ) );
NAND2_X4 _add_3_root_add_136_4_U90  ( .A1(SHA1_ft_BCD[13]), .A2(SHA1_result_136), .ZN(_add_3_root_add_136_4_n325 ) );
NAND2_X1 _add_3_root_add_136_4_U89  ( .A1(_add_3_root_add_136_4_n322 ), .A2(_add_3_root_add_136_4_n325 ), .ZN(_add_3_root_add_136_4_n347 ) );
NOR2_X2 _add_3_root_add_136_4_U88  ( .A1(_add_3_root_add_136_4_n98 ), .A2(_add_3_root_add_136_4_n361 ), .ZN(_add_3_root_add_136_4_n375 ) );
INV_X2 _add_3_root_add_136_4_U87  ( .A(SHA1_ft_BCD[8]), .ZN(_add_3_root_add_136_4_n392 ) );
NAND2_X4 _add_3_root_add_136_4_U86  ( .A1(_add_3_root_add_136_4_n392 ), .A2(_add_3_root_add_136_4_n393 ), .ZN(_add_3_root_add_136_4_n104 ) );
INV_X8 _add_3_root_add_136_4_U85  ( .A(_add_3_root_add_136_4_n104 ), .ZN(_add_3_root_add_136_4_n98 ) );
NOR2_X2 _add_3_root_add_136_4_U84  ( .A1(_add_3_root_add_136_4_n105 ), .A2(_add_3_root_add_136_4_n100 ), .ZN(_add_3_root_add_136_4_n103 ) );
BUF_X8 _add_3_root_add_136_4_U83  ( .A(_add_3_root_add_136_4_n352 ), .Z(_add_3_root_add_136_4_n26 ) );
INV_X8 _add_3_root_add_136_4_U82  ( .A(_add_3_root_add_136_4_n92 ), .ZN(_add_3_root_add_136_4_n361 ) );
NOR2_X4 _add_3_root_add_136_4_U81  ( .A1(_add_3_root_add_136_4_n126 ), .A2(_add_3_root_add_136_4_n15 ), .ZN(_add_3_root_add_136_4_n124 ) );
NAND2_X4 _add_3_root_add_136_4_U80  ( .A1(_add_3_root_add_136_4_n243 ), .A2(_add_3_root_add_136_4_n244 ), .ZN(_add_3_root_add_136_4_n242 ) );
INV_X1 _add_3_root_add_136_4_U79  ( .A(_add_3_root_add_136_4_n242 ), .ZN(_add_3_root_add_136_4_n25 ) );
NOR2_X4 _add_3_root_add_136_4_U78  ( .A1(_add_3_root_add_136_4_n98 ), .A2(_add_3_root_add_136_4_n361 ), .ZN(_add_3_root_add_136_4_n364 ) );
AND2_X4 _add_3_root_add_136_4_U77  ( .A1(_add_3_root_add_136_4_n165 ), .A2(_add_3_root_add_136_4_n73 ), .ZN(_add_3_root_add_136_4_n126 ) );
NAND2_X2 _add_3_root_add_136_4_U76  ( .A1(_add_3_root_add_136_4_n290 ), .A2(_add_3_root_add_136_4_n287 ), .ZN(_add_3_root_add_136_4_n288 ) );
AND2_X2 _add_3_root_add_136_4_U75  ( .A1(_add_3_root_add_136_4_n165 ), .A2(_add_3_root_add_136_4_n164 ), .ZN(_add_3_root_add_136_4_n22 ) );
XNOR2_X2 _add_3_root_add_136_4_U74  ( .A(_add_3_root_add_136_4_n22 ), .B(_add_3_root_add_136_4_n163 ), .ZN(N65) );
INV_X8 _add_3_root_add_136_4_U73  ( .A(SHA1_ft_BCD[2]), .ZN(_add_3_root_add_136_4_n384 ) );
NOR2_X2 _add_3_root_add_136_4_U72  ( .A1(_add_3_root_add_136_4_n363 ), .A2(_add_3_root_add_136_4_n191 ), .ZN(_add_3_root_add_136_4_n355 ) );
INV_X4 _add_3_root_add_136_4_U71  ( .A(_add_3_root_add_136_4_n20 ), .ZN(_add_3_root_add_136_4_n21 ) );
INV_X4 _add_3_root_add_136_4_U70  ( .A(_add_3_root_add_136_4_n35 ), .ZN(_add_3_root_add_136_4_n20 ) );
NAND2_X2 _add_3_root_add_136_4_U69  ( .A1(_add_3_root_add_136_4_n285 ), .A2(_add_3_root_add_136_4_n23 ), .ZN(_add_3_root_add_136_4_n281 ) );
INV_X4 _add_3_root_add_136_4_U68  ( .A(_add_3_root_add_136_4_n18 ), .ZN(_add_3_root_add_136_4_n362 ) );
NOR2_X4 _add_3_root_add_136_4_U67  ( .A1(SHA1_ft_BCD[10]), .A2(SHA1_result_133), .ZN(_add_3_root_add_136_4_n18 ) );
NAND2_X2 _add_3_root_add_136_4_U66  ( .A1(_add_3_root_add_136_4_n226 ), .A2(_add_3_root_add_136_4_n227 ), .ZN(_add_3_root_add_136_4_n222 ) );
NAND2_X2 _add_3_root_add_136_4_U65  ( .A1(SHA1_ft_BCD[18]), .A2(n14431),.ZN(_add_3_root_add_136_4_n289 ) );
NAND2_X1 _add_3_root_add_136_4_U64  ( .A1(_add_3_root_add_136_4_n287 ), .A2(_add_3_root_add_136_4_n289 ), .ZN(_add_3_root_add_136_4_n292 ) );
AND2_X2 _add_3_root_add_136_4_U63  ( .A1(_add_3_root_add_136_4_n288 ), .A2(_add_3_root_add_136_4_n289 ), .ZN(_add_3_root_add_136_4_n23 ) );
INV_X2 _add_3_root_add_136_4_U62  ( .A(_add_3_root_add_136_4_n364 ), .ZN(_add_3_root_add_136_4_n19 ) );
AND2_X2 _add_3_root_add_136_4_U61  ( .A1(_add_3_root_add_136_4_n286 ), .A2(_add_3_root_add_136_4_n287 ), .ZN(_add_3_root_add_136_4_n78 ) );
AND2_X4 _add_3_root_add_136_4_U60  ( .A1(_add_3_root_add_136_4_n148 ), .A2(_add_3_root_add_136_4_n172 ), .ZN(_add_3_root_add_136_4_n17 ) );
AND2_X2 _add_3_root_add_136_4_U59  ( .A1(_add_3_root_add_136_4_n95 ), .A2(_add_3_root_add_136_4_n104 ), .ZN(_add_3_root_add_136_4_n16 ) );
INV_X1 _add_3_root_add_136_4_U58  ( .A(_add_3_root_add_136_4_n208 ), .ZN(_add_3_root_add_136_4_n229 ) );
AND2_X4 _add_3_root_add_136_4_U57  ( .A1(_add_3_root_add_136_4_n384 ), .A2(_add_3_root_add_136_4_n385 ), .ZN(_add_3_root_add_136_4_n15 ) );
AND2_X2 _add_3_root_add_136_4_U56  ( .A1(_add_3_root_add_136_4_n78 ), .A2(_add_3_root_add_136_4_n277 ), .ZN(_add_3_root_add_136_4_n14 ) );
BUF_X4 _add_3_root_add_136_4_U55  ( .A(_add_3_root_add_136_4_n83 ), .Z(_add_3_root_add_136_4_n40 ) );
INV_X4 _add_3_root_add_136_4_U54  ( .A(_add_3_root_add_136_4_n101 ), .ZN(_add_3_root_add_136_4_n86 ) );
NAND2_X4 _add_3_root_add_136_4_U53  ( .A1(_add_3_root_add_136_4_n280 ), .A2(_add_3_root_add_136_4_n165 ), .ZN(_add_3_root_add_136_4_n315 ) );
NAND4_X1 _add_3_root_add_136_4_U52  ( .A1(_add_3_root_add_136_4_n186 ), .A2(_add_3_root_add_136_4_n187 ), .A3(_add_3_root_add_136_4_n188 ), .A4(_add_3_root_add_136_4_n189 ), .ZN(_add_3_root_add_136_4_n182 ) );
NOR2_X1 _add_3_root_add_136_4_U51  ( .A1(_add_3_root_add_136_4_n173 ), .A2(_add_3_root_add_136_4_n237 ), .ZN(_add_3_root_add_136_4_n247 ) );
NAND2_X2 _add_3_root_add_136_4_U50  ( .A1(_add_3_root_add_136_4_n27 ), .A2(_add_3_root_add_136_4_n295 ), .ZN(_add_3_root_add_136_4_n291 ) );
INV_X4 _add_3_root_add_136_4_U49  ( .A(SHA1_result_129), .ZN(_add_3_root_add_136_4_n31 ) );
INV_X4 _add_3_root_add_136_4_U48  ( .A(_add_3_root_add_136_4_n371 ), .ZN(_add_3_root_add_136_4_n61 ) );
NAND2_X2 _add_3_root_add_136_4_U47  ( .A1(_add_3_root_add_136_4_n321 ), .A2(_add_3_root_add_136_4_n24 ), .ZN(_add_3_root_add_136_4_n319 ) );
NAND2_X2 _add_3_root_add_136_4_U46  ( .A1(_add_3_root_add_136_4_n241 ), .A2(_add_3_root_add_136_4_n14 ), .ZN(_add_3_root_add_136_4_n276 ) );
NAND2_X2 _add_3_root_add_136_4_U45  ( .A1(_add_3_root_add_136_4_n276 ), .A2(_add_3_root_add_136_4_n275 ), .ZN(_add_3_root_add_136_4_n264 ) );
INV_X4 _add_3_root_add_136_4_U44  ( .A(_add_3_root_add_136_4_n264 ), .ZN(_add_3_root_add_136_4_n256 ) );
NOR2_X2 _add_3_root_add_136_4_U43  ( .A1(_add_3_root_add_136_4_n89 ), .A2(_add_3_root_add_136_4_n40 ), .ZN(_add_3_root_add_136_4_n117 ) );
NOR2_X4 _add_3_root_add_136_4_U42  ( .A1(SHA1_ft_BCD[4]), .A2(n14464), .ZN(_add_3_root_add_136_4_n83 ) );
NOR2_X4 _add_3_root_add_136_4_U41  ( .A1(_add_3_root_add_136_4_n97 ), .A2(_add_3_root_add_136_4_n98 ), .ZN(_add_3_root_add_136_4_n96 ) );
NAND2_X4 _add_3_root_add_136_4_U40  ( .A1(_add_3_root_add_136_4_n114 ), .A2(_add_3_root_add_136_4_n115 ), .ZN(_add_3_root_add_136_4_n397 ) );
INV_X1 _add_3_root_add_136_4_U39  ( .A(_add_3_root_add_136_4_n114 ), .ZN(_add_3_root_add_136_4_n121 ) );
NAND2_X2 _add_3_root_add_136_4_U38  ( .A1(_add_3_root_add_136_4_n241 ), .A2(_add_3_root_add_136_4_n332 ), .ZN(_add_3_root_add_136_4_n306 ) );
XNOR2_X2 _add_3_root_add_136_4_U37  ( .A(_add_3_root_add_136_4_n91 ), .B(_add_3_root_add_136_4_n12 ), .ZN(N73) );
NOR2_X4 _add_3_root_add_136_4_U36  ( .A1(_add_3_root_add_136_4_n87 ), .A2(_add_3_root_add_136_4_n102 ), .ZN(_add_3_root_add_136_4_n105 ) );
NAND2_X1 _add_3_root_add_136_4_U35  ( .A1(_add_3_root_add_136_4_n29 ), .A2(_add_3_root_add_136_4_n93 ), .ZN(_add_3_root_add_136_4_n12 ) );
AND2_X4 _add_3_root_add_136_4_U34  ( .A1(_add_3_root_add_136_4_n200 ), .A2(_add_3_root_add_136_4_n211 ), .ZN(_add_3_root_add_136_4_n11 ) );
AND2_X4 _add_3_root_add_136_4_U33  ( .A1(SHA1_ft_BCD[3]), .A2(n14382), .ZN(_add_3_root_add_136_4_n10 ) );
AND2_X2 _add_3_root_add_136_4_U32  ( .A1(SHA1_ft_BCD[21]), .A2(n14422), .ZN(_add_3_root_add_136_4_n9 ) );
NAND2_X2 _add_3_root_add_136_4_U31  ( .A1(_add_3_root_add_136_4_n94 ), .A2(_add_3_root_add_136_4_n95 ), .ZN(_add_3_root_add_136_4_n91 ) );
NOR2_X2 _add_3_root_add_136_4_U30  ( .A1(_add_3_root_add_136_4_n355 ), .A2(_add_3_root_add_136_4_n26 ), .ZN(_add_3_root_add_136_4_n65 ) );
NOR2_X2 _add_3_root_add_136_4_U29  ( .A1(_add_3_root_add_136_4_n67 ), .A2(_add_3_root_add_136_4_n190 ), .ZN(_add_3_root_add_136_4_n37 ) );
NAND2_X2 _add_3_root_add_136_4_U28  ( .A1(_add_3_root_add_136_4_n319 ), .A2(_add_3_root_add_136_4_n320 ), .ZN(_add_3_root_add_136_4_n183 ) );
NAND2_X4 _add_3_root_add_136_4_U27  ( .A1(_add_3_root_add_136_4_n118 ), .A2(_add_3_root_add_136_4_n57 ), .ZN(_add_3_root_add_136_4_n58 ) );
NOR2_X4 _add_3_root_add_136_4_U26  ( .A1(_add_3_root_add_136_4_n87 ), .A2(_add_3_root_add_136_4_n40 ), .ZN(_add_3_root_add_136_4_n120 ) );
INV_X8 _add_3_root_add_136_4_U25  ( .A(_add_3_root_add_136_4_n109 ), .ZN(_add_3_root_add_136_4_n401 ) );
INV_X1 _add_3_root_add_136_4_U24  ( .A(_add_3_root_add_136_4_n401 ), .ZN(_add_3_root_add_136_4_n8 ) );
INV_X8 _add_3_root_add_136_4_U23  ( .A(_add_3_root_add_136_4_n21 ), .ZN(_add_3_root_add_136_4_n111 ) );
OR3_X4 _add_3_root_add_136_4_U22  ( .A1(_add_3_root_add_136_4_n322 ), .A2(_add_3_root_add_136_4_n79 ), .A3(_add_3_root_add_136_4_n28 ), .ZN(_add_3_root_add_136_4_n24 ) );
NOR2_X4 _add_3_root_add_136_4_U21  ( .A1(_add_3_root_add_136_4_n265 ), .A2(_add_3_root_add_136_4_n256 ), .ZN(_add_3_root_add_136_4_n269 ) );
NOR2_X2 _add_3_root_add_136_4_U20  ( .A1(_add_3_root_add_136_4_n35 ), .A2(_add_3_root_add_136_4_n387 ), .ZN(_add_3_root_add_136_4_n396 ) );
AND2_X2 _add_3_root_add_136_4_U19  ( .A1(_add_3_root_add_136_4_n329 ), .A2(_add_3_root_add_136_4_n325 ), .ZN(_add_3_root_add_136_4_n7 ) );
XNOR2_X2 _add_3_root_add_136_4_U18  ( .A(_add_3_root_add_136_4_n349 ), .B(_add_3_root_add_136_4_n7 ), .ZN(_add_3_root_add_136_4_n6 ) );
NOR2_X4 _add_3_root_add_136_4_U17  ( .A1(_add_3_root_add_136_4_n83 ), .A2(_add_3_root_add_136_4_n387 ), .ZN(_add_3_root_add_136_4_n386 ) );
OR3_X2 _add_3_root_add_136_4_U16  ( .A1(_add_3_root_add_136_4_n342 ), .A2(_add_3_root_add_136_4_n350 ), .A3(_add_3_root_add_136_4_n70 ), .ZN(_add_3_root_add_136_4_n5 ) );
AND2_X2 _add_3_root_add_136_4_U15  ( .A1(_add_3_root_add_136_4_n112 ), .A2(_add_3_root_add_136_4_n111 ), .ZN(_add_3_root_add_136_4_n4 ) );
AND2_X2 _add_3_root_add_136_4_U14  ( .A1(_add_3_root_add_136_4_n322 ), .A2(_add_3_root_add_136_4_n328 ), .ZN(_add_3_root_add_136_4_n3 ) );
NOR2_X4 _add_3_root_add_136_4_U13  ( .A1(_add_3_root_add_136_4_n400 ), .A2(_add_3_root_add_136_4_n31 ), .ZN(_add_3_root_add_136_4_n30 ) );
INV_X4 _add_3_root_add_136_4_U12  ( .A(_add_3_root_add_136_4_n30 ), .ZN(_add_3_root_add_136_4_n38 ) );
NAND2_X2 _add_3_root_add_136_4_U11  ( .A1(_add_3_root_add_136_4_n113 ), .A2(_add_3_root_add_136_4_n4 ), .ZN(_add_3_root_add_136_4_n110 ) );
NAND2_X2 _add_3_root_add_136_4_U10  ( .A1(_add_3_root_add_136_4_n279 ), .A2(_add_3_root_add_136_4_n164 ), .ZN(_add_3_root_add_136_4_n73 ) );
AND2_X2 _add_3_root_add_136_4_U9  ( .A1(_add_3_root_add_136_4_n115 ), .A2(_add_3_root_add_136_4_n112 ), .ZN(_add_3_root_add_136_4_n2 ) );
XNOR2_X2 _add_3_root_add_136_4_U8  ( .A(_add_3_root_add_136_4_n119 ), .B(_add_3_root_add_136_4_n2 ), .ZN(N69) );
INV_X1 _add_3_root_add_136_4_U7  ( .A(SHA1_ft_BCD[14]), .ZN(_add_3_root_add_136_4_n33 ) );
NOR2_X1 _add_3_root_add_136_4_U6  ( .A1(_add_3_root_add_136_4_n79 ), .A2(_add_3_root_add_136_4_n325 ), .ZN(_add_3_root_add_136_4_n323 ) );
NAND2_X2 _add_3_root_add_136_4_U5  ( .A1(n14929), .A2(n14388), .ZN(_add_3_root_add_136_4_n165 ) );
INV_X2 _add_3_root_add_136_4_U4  ( .A(SHA1_ft_BCD[12]), .ZN(_add_3_root_add_136_4_n353 ) );
NOR3_X2 _add_3_root_add_136_4_U3  ( .A1(_add_3_root_add_136_4_n377 ), .A2(_add_3_root_add_136_4_n317 ), .A3(_add_3_root_add_136_4_n10 ), .ZN(_add_3_root_add_136_4_n89 ) );
NOR3_X4 _add_3_root_add_136_4_U2  ( .A1(_add_3_root_add_136_4_n377 ), .A2(_add_3_root_add_136_4_n317 ), .A3(_add_3_root_add_136_4_n10 ), .ZN(_add_3_root_add_136_4_n101 ) );
NAND2_X2 _add_2_root_add_136_4_U468  ( .A1(Kt[0]), .A2(SHA1_result[0]), .ZN(_add_2_root_add_136_4_n327 ) );
NAND2_X2 _add_2_root_add_136_4_U467  ( .A1(Kt[10]), .A2(SHA1_result[10]),.ZN(_add_2_root_add_136_4_n418 ) );
INV_X4 _add_2_root_add_136_4_U466  ( .A(_add_2_root_add_136_4_n418 ), .ZN(_add_2_root_add_136_4_n406 ) );
NAND2_X2 _add_2_root_add_136_4_U465  ( .A1(Kt[9]), .A2(SHA1_result[9]), .ZN(_add_2_root_add_136_4_n420 ) );
INV_X4 _add_2_root_add_136_4_U464  ( .A(_add_2_root_add_136_4_n420 ), .ZN(_add_2_root_add_136_4_n46 ) );
NAND2_X2 _add_2_root_add_136_4_U463  ( .A1(Kt[0]), .A2(SHA1_result[0]), .ZN(_add_2_root_add_136_4_n436 ) );
NAND2_X2 _add_2_root_add_136_4_U462  ( .A1(Kt[1]), .A2(SHA1_result[1]), .ZN(_add_2_root_add_136_4_n437 ) );
NAND2_X2 _add_2_root_add_136_4_U461  ( .A1(_add_2_root_add_136_4_n436 ),.A2(_add_2_root_add_136_4_n437 ), .ZN(_add_2_root_add_136_4_n434 ) );
INV_X4 _add_2_root_add_136_4_U460  ( .A(_add_2_root_add_136_4_n155 ), .ZN(_add_2_root_add_136_4_n354 ) );
INV_X4 _add_2_root_add_136_4_U459  ( .A(_add_2_root_add_136_4_n353 ), .ZN(_add_2_root_add_136_4_n84 ) );
NAND2_X2 _add_2_root_add_136_4_U458  ( .A1(Kt[3]), .A2(SHA1_result[3]), .ZN(_add_2_root_add_136_4_n241 ) );
INV_X4 _add_2_root_add_136_4_U457  ( .A(_add_2_root_add_136_4_n241 ), .ZN(_add_2_root_add_136_4_n83 ) );
INV_X4 _add_2_root_add_136_4_U456  ( .A(_add_2_root_add_136_4_n394 ), .ZN(_add_2_root_add_136_4_n53 ) );
NAND2_X2 _add_2_root_add_136_4_U455  ( .A1(Kt[7]), .A2(SHA1_result[7]), .ZN(_add_2_root_add_136_4_n62 ) );
NAND2_X2 _add_2_root_add_136_4_U454  ( .A1(Kt[4]), .A2(SHA1_result[4]), .ZN(_add_2_root_add_136_4_n429 ) );
NAND2_X2 _add_2_root_add_136_4_U453  ( .A1(Kt[5]), .A2(SHA1_result[5]), .ZN(_add_2_root_add_136_4_n69 ) );
NAND2_X2 _add_2_root_add_136_4_U452  ( .A1(_add_2_root_add_136_4_n429 ),.A2(_add_2_root_add_136_4_n69 ), .ZN(_add_2_root_add_136_4_n428 ) );
NAND2_X2 _add_2_root_add_136_4_U451  ( .A1(_add_2_root_add_136_4_n427 ),.A2(_add_2_root_add_136_4_n428 ), .ZN(_add_2_root_add_136_4_n426 ) );
XNOR2_X2 _add_2_root_add_136_4_U450  ( .A(_add_2_root_add_136_4_n422 ), .B(_add_2_root_add_136_4_n423 ), .ZN(N106) );
NAND2_X2 _add_2_root_add_136_4_U449  ( .A1(_add_2_root_add_136_4_n31 ), .A2(_add_2_root_add_136_4_n418 ), .ZN(_add_2_root_add_136_4_n417 ) );
XNOR2_X2 _add_2_root_add_136_4_U448  ( .A(_add_2_root_add_136_4_n414 ), .B(_add_2_root_add_136_4_n415 ), .ZN(N107) );
NAND2_X2 _add_2_root_add_136_4_U447  ( .A1(_add_2_root_add_136_4_n185 ),.A2(_add_2_root_add_136_4_n52 ), .ZN(_add_2_root_add_136_4_n400 ) );
NAND2_X2 _add_2_root_add_136_4_U446  ( .A1(_add_2_root_add_136_4_n407 ),.A2(_add_2_root_add_136_4_n408 ), .ZN(_add_2_root_add_136_4_n403 ) );
INV_X4 _add_2_root_add_136_4_U445  ( .A(_add_2_root_add_136_4_n402 ), .ZN(_add_2_root_add_136_4_n362 ) );
NAND2_X2 _add_2_root_add_136_4_U444  ( .A1(_add_2_root_add_136_4_n363 ),.A2(_add_2_root_add_136_4_n362 ), .ZN(_add_2_root_add_136_4_n392 ) );
INV_X4 _add_2_root_add_136_4_U443  ( .A(_add_2_root_add_136_4_n54 ), .ZN(_add_2_root_add_136_4_n242 ) );
NAND2_X2 _add_2_root_add_136_4_U442  ( .A1(_add_2_root_add_136_4_n242 ),.A2(_add_2_root_add_136_4_n185 ), .ZN(_add_2_root_add_136_4_n401 ) );
NAND2_X2 _add_2_root_add_136_4_U441  ( .A1(Kt[12]), .A2(SHA1_result[12]),.ZN(_add_2_root_add_136_4_n393 ) );
INV_X4 _add_2_root_add_136_4_U440  ( .A(_add_2_root_add_136_4_n393 ), .ZN(_add_2_root_add_136_4_n360 ) );
XNOR2_X2 _add_2_root_add_136_4_U439  ( .A(_add_2_root_add_136_4_n24 ), .B(_add_2_root_add_136_4_n399 ), .ZN(N108) );
NAND2_X2 _add_2_root_add_136_4_U438  ( .A1(_add_2_root_add_136_4_n37 ), .A2(_add_2_root_add_136_4_n393 ), .ZN(_add_2_root_add_136_4_n396 ) );
NAND2_X2 _add_2_root_add_136_4_U437  ( .A1(Kt[13]), .A2(SHA1_result[13]),.ZN(_add_2_root_add_136_4_n370 ) );
INV_X4 _add_2_root_add_136_4_U436  ( .A(_add_2_root_add_136_4_n370 ), .ZN(_add_2_root_add_136_4_n398 ) );
INV_X4 _add_2_root_add_136_4_U435  ( .A(_add_2_root_add_136_4_n52 ), .ZN(_add_2_root_add_136_4_n395 ) );
NAND2_X2 _add_2_root_add_136_4_U434  ( .A1(_add_2_root_add_136_4_n392 ),.A2(_add_2_root_add_136_4_n393 ), .ZN(_add_2_root_add_136_4_n391 ) );
NAND2_X2 _add_2_root_add_136_4_U433  ( .A1(Kt[14]), .A2(SHA1_result[14]),.ZN(_add_2_root_add_136_4_n371 ) );
INV_X4 _add_2_root_add_136_4_U432  ( .A(_add_2_root_add_136_4_n371 ), .ZN(_add_2_root_add_136_4_n388 ) );
XNOR2_X2 _add_2_root_add_136_4_U431  ( .A(_add_2_root_add_136_4_n386 ), .B(_add_2_root_add_136_4_n387 ), .ZN(N110) );
NAND2_X2 _add_2_root_add_136_4_U430  ( .A1(_add_2_root_add_136_4_n36 ), .A2(_add_2_root_add_136_4_n371 ), .ZN(_add_2_root_add_136_4_n382 ) );
NAND2_X2 _add_2_root_add_136_4_U429  ( .A1(Kt[15]), .A2(SHA1_result[15]),.ZN(_add_2_root_add_136_4_n132 ) );
INV_X4 _add_2_root_add_136_4_U428  ( .A(_add_2_root_add_136_4_n132 ), .ZN(_add_2_root_add_136_4_n252 ) );
XNOR2_X2 _add_2_root_add_136_4_U427  ( .A(_add_2_root_add_136_4_n379 ), .B(_add_2_root_add_136_4_n380 ), .ZN(N111) );
NAND2_X2 _add_2_root_add_136_4_U426  ( .A1(Kt[4]), .A2(SHA1_result[4]), .ZN(_add_2_root_add_136_4_n68 ) );
NAND2_X2 _add_2_root_add_136_4_U425  ( .A1(_add_2_root_add_136_4_n68 ), .A2(_add_2_root_add_136_4_n69 ), .ZN(_add_2_root_add_136_4_n238 ) );
INV_X4 _add_2_root_add_136_4_U424  ( .A(_add_2_root_add_136_4_n65 ), .ZN(_add_2_root_add_136_4_n373 ) );
INV_X4 _add_2_root_add_136_4_U423  ( .A(_add_2_root_add_136_4_n61 ), .ZN(_add_2_root_add_136_4_n374 ) );
INV_X4 _add_2_root_add_136_4_U422  ( .A(_add_2_root_add_136_4_n64 ), .ZN(_add_2_root_add_136_4_n375 ) );
INV_X4 _add_2_root_add_136_4_U421  ( .A(_add_2_root_add_136_4_n278 ), .ZN(_add_2_root_add_136_4_n127 ) );
NAND2_X2 _add_2_root_add_136_4_U420  ( .A1(_add_2_root_add_136_4_n370 ),.A2(_add_2_root_add_136_4_n371 ), .ZN(_add_2_root_add_136_4_n366 ) );
INV_X4 _add_2_root_add_136_4_U419  ( .A(_add_2_root_add_136_4_n368 ), .ZN(_add_2_root_add_136_4_n367 ) );
AND3_X2 _add_2_root_add_136_4_U418  ( .A1(_add_2_root_add_136_4_n366 ), .A2(_add_2_root_add_136_4_n42 ), .A3(_add_2_root_add_136_4_n367 ), .ZN(_add_2_root_add_136_4_n128 ) );
NAND2_X2 _add_2_root_add_136_4_U417  ( .A1(_add_2_root_add_136_4_n364 ),.A2(_add_2_root_add_136_4_n365 ), .ZN(_add_2_root_add_136_4_n123 ) );
INV_X4 _add_2_root_add_136_4_U416  ( .A(_add_2_root_add_136_4_n123 ), .ZN(_add_2_root_add_136_4_n355 ) );
INV_X4 _add_2_root_add_136_4_U415  ( .A(_add_2_root_add_136_4_n1 ), .ZN(_add_2_root_add_136_4_n237 ) );
NAND2_X2 _add_2_root_add_136_4_U414  ( .A1(_add_2_root_add_136_4_n361 ),.A2(_add_2_root_add_136_4_n185 ), .ZN(_add_2_root_add_136_4_n130 ) );
NAND2_X2 _add_2_root_add_136_4_U413  ( .A1(_add_2_root_add_136_4_n360 ),.A2(_add_2_root_add_136_4_n237 ), .ZN(_add_2_root_add_136_4_n131 ) );
NAND4_X2 _add_2_root_add_136_4_U412  ( .A1(_add_2_root_add_136_4_n129 ),.A2(_add_2_root_add_136_4_n130 ), .A3(_add_2_root_add_136_4_n131 ),.A4(_add_2_root_add_136_4_n132 ), .ZN(_add_2_root_add_136_4_n356 ) );
NAND2_X2 _add_2_root_add_136_4_U411  ( .A1(_add_2_root_add_136_4_n358 ),.A2(_add_2_root_add_136_4_n359 ), .ZN(_add_2_root_add_136_4_n122 ) );
INV_X4 _add_2_root_add_136_4_U410  ( .A(_add_2_root_add_136_4_n122 ), .ZN(_add_2_root_add_136_4_n357 ) );
INV_X4 _add_2_root_add_136_4_U409  ( .A(_add_2_root_add_136_4_n86 ), .ZN(_add_2_root_add_136_4_n352 ) );
NAND2_X2 _add_2_root_add_136_4_U408  ( .A1(Kt[1]), .A2(SHA1_result[1]), .ZN(_add_2_root_add_136_4_n156 ) );
NAND2_X2 _add_2_root_add_136_4_U407  ( .A1(_add_2_root_add_136_4_n327 ),.A2(_add_2_root_add_136_4_n156 ), .ZN(_add_2_root_add_136_4_n250 ) );
INV_X4 _add_2_root_add_136_4_U406  ( .A(_add_2_root_add_136_4_n250 ), .ZN(_add_2_root_add_136_4_n351 ) );
NAND4_X2 _add_2_root_add_136_4_U405  ( .A1(_add_2_root_add_136_4_n34 ), .A2(_add_2_root_add_136_4_n185 ), .A3(_add_2_root_add_136_4_n350 ), .A4(_add_2_root_add_136_4_n237 ), .ZN(_add_2_root_add_136_4_n125 ) );
NAND2_X2 _add_2_root_add_136_4_U404  ( .A1(Kt[16]), .A2(SHA1_result[16]),.ZN(_add_2_root_add_136_4_n345 ) );
NAND2_X2 _add_2_root_add_136_4_U403  ( .A1(_add_2_root_add_136_4_n43 ), .A2(_add_2_root_add_136_4_n345 ), .ZN(_add_2_root_add_136_4_n347 ) );
XNOR2_X2 _add_2_root_add_136_4_U402  ( .A(_add_2_root_add_136_4_n306 ), .B(_add_2_root_add_136_4_n347 ), .ZN(N112) );
NAND2_X2 _add_2_root_add_136_4_U401  ( .A1(_add_2_root_add_136_4_n306 ),.A2(_add_2_root_add_136_4_n43 ), .ZN(_add_2_root_add_136_4_n346 ) );
NAND2_X2 _add_2_root_add_136_4_U400  ( .A1(_add_2_root_add_136_4_n345 ),.A2(_add_2_root_add_136_4_n346 ), .ZN(_add_2_root_add_136_4_n343 ) );
NAND2_X2 _add_2_root_add_136_4_U399  ( .A1(Kt[17]), .A2(SHA1_result[17]),.ZN(_add_2_root_add_136_4_n340 ) );
NAND2_X2 _add_2_root_add_136_4_U398  ( .A1(_add_2_root_add_136_4_n340 ),.A2(_add_2_root_add_136_4_n342 ), .ZN(_add_2_root_add_136_4_n344 ) );
XNOR2_X2 _add_2_root_add_136_4_U397  ( .A(_add_2_root_add_136_4_n343 ), .B(_add_2_root_add_136_4_n344 ), .ZN(N113) );
INV_X4 _add_2_root_add_136_4_U396  ( .A(_add_2_root_add_136_4_n336 ), .ZN(_add_2_root_add_136_4_n342 ) );
INV_X4 _add_2_root_add_136_4_U395  ( .A(SHA1_result[18]), .ZN(_add_2_root_add_136_4_n338 ) );
NAND2_X2 _add_2_root_add_136_4_U394  ( .A1(_add_2_root_add_136_4_n324 ),.A2(_add_2_root_add_136_4_n306 ), .ZN(_add_2_root_add_136_4_n332 ) );
NAND2_X2 _add_2_root_add_136_4_U393  ( .A1(_add_2_root_add_136_4_n263 ),.A2(_add_2_root_add_136_4_n332 ), .ZN(_add_2_root_add_136_4_n328 ) );
NAND2_X2 _add_2_root_add_136_4_U392  ( .A1(Kt[19]), .A2(SHA1_result[19]),.ZN(_add_2_root_add_136_4_n116 ) );
INV_X4 _add_2_root_add_136_4_U391  ( .A(Kt[19]), .ZN(_add_2_root_add_136_4_n330 ) );
INV_X4 _add_2_root_add_136_4_U390  ( .A(SHA1_result[19]), .ZN(_add_2_root_add_136_4_n331 ) );
NAND2_X2 _add_2_root_add_136_4_U389  ( .A1(_add_2_root_add_136_4_n330 ),.A2(_add_2_root_add_136_4_n331 ), .ZN(_add_2_root_add_136_4_n265 ) );
NAND2_X2 _add_2_root_add_136_4_U388  ( .A1(_add_2_root_add_136_4_n116 ),.A2(_add_2_root_add_136_4_n265 ), .ZN(_add_2_root_add_136_4_n329 ) );
XNOR2_X2 _add_2_root_add_136_4_U387  ( .A(_add_2_root_add_136_4_n328 ), .B(_add_2_root_add_136_4_n329 ), .ZN(N115) );
INV_X4 _add_2_root_add_136_4_U386  ( .A(_add_2_root_add_136_4_n156 ), .ZN(_add_2_root_add_136_4_n326 ) );
XNOR2_X2 _add_2_root_add_136_4_U385  ( .A(_add_2_root_add_136_4_n436 ), .B(_add_2_root_add_136_4_n325 ), .ZN(N97) );
INV_X4 _add_2_root_add_136_4_U384  ( .A(_add_2_root_add_136_4_n306 ), .ZN(_add_2_root_add_136_4_n153 ) );
NAND2_X2 _add_2_root_add_136_4_U383  ( .A1(_add_2_root_add_136_4_n264 ),.A2(_add_2_root_add_136_4_n265 ), .ZN(_add_2_root_add_136_4_n112 ) );
NAND2_X2 _add_2_root_add_136_4_U382  ( .A1(_add_2_root_add_136_4_n112 ),.A2(_add_2_root_add_136_4_n116 ), .ZN(_add_2_root_add_136_4_n296 ) );
XNOR2_X2 _add_2_root_add_136_4_U381  ( .A(_add_2_root_add_136_4_n321 ), .B(_add_2_root_add_136_4_n322 ), .ZN(N116) );
NAND4_X2 _add_2_root_add_136_4_U380  ( .A1(_add_2_root_add_136_4_n129 ),.A2(_add_2_root_add_136_4_n130 ), .A3(_add_2_root_add_136_4_n131 ),.A4(_add_2_root_add_136_4_n132 ), .ZN(_add_2_root_add_136_4_n317 ) );
NAND2_X2 _add_2_root_add_136_4_U379  ( .A1(_add_2_root_add_136_4_n122 ),.A2(_add_2_root_add_136_4_n123 ), .ZN(_add_2_root_add_136_4_n319 ) );
NAND2_X2 _add_2_root_add_136_4_U378  ( .A1(Kt[21]), .A2(SHA1_result[21]),.ZN(_add_2_root_add_136_4_n309 ) );
INV_X4 _add_2_root_add_136_4_U377  ( .A(_add_2_root_add_136_4_n309 ), .ZN(_add_2_root_add_136_4_n312 ) );
XNOR2_X2 _add_2_root_add_136_4_U376  ( .A(_add_2_root_add_136_4_n310 ), .B(_add_2_root_add_136_4_n311 ), .ZN(N117) );
NAND2_X2 _add_2_root_add_136_4_U375  ( .A1(_add_2_root_add_136_4_n296 ),.A2(_add_2_root_add_136_4_n305 ), .ZN(_add_2_root_add_136_4_n301 ) );
NAND2_X2 _add_2_root_add_136_4_U374  ( .A1(Kt[20]), .A2(SHA1_result[20]),.ZN(_add_2_root_add_136_4_n308 ) );
NAND2_X2 _add_2_root_add_136_4_U373  ( .A1(_add_2_root_add_136_4_n308 ),.A2(_add_2_root_add_136_4_n309 ), .ZN(_add_2_root_add_136_4_n307 ) );
NAND2_X2 _add_2_root_add_136_4_U372  ( .A1(_add_2_root_add_136_4_n307 ),.A2(_add_2_root_add_136_4_n289 ), .ZN(_add_2_root_add_136_4_n302 ) );
INV_X4 _add_2_root_add_136_4_U371  ( .A(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n304 ) );
NAND2_X2 _add_2_root_add_136_4_U370  ( .A1(Kt[22]), .A2(SHA1_result[22]),.ZN(_add_2_root_add_136_4_n287 ) );
INV_X4 _add_2_root_add_136_4_U369  ( .A(Kt[22]), .ZN(_add_2_root_add_136_4_n299 ) );
INV_X4 _add_2_root_add_136_4_U368  ( .A(SHA1_result[22]), .ZN(_add_2_root_add_136_4_n300 ) );
NAND2_X2 _add_2_root_add_136_4_U367  ( .A1(_add_2_root_add_136_4_n299 ),.A2(_add_2_root_add_136_4_n300 ), .ZN(_add_2_root_add_136_4_n163 ) );
NAND2_X2 _add_2_root_add_136_4_U366  ( .A1(_add_2_root_add_136_4_n287 ),.A2(_add_2_root_add_136_4_n163 ), .ZN(_add_2_root_add_136_4_n298 ) );
XNOR2_X2 _add_2_root_add_136_4_U365  ( .A(_add_2_root_add_136_4_n297 ), .B(_add_2_root_add_136_4_n298 ), .ZN(N118) );
INV_X4 _add_2_root_add_136_4_U364  ( .A(_add_2_root_add_136_4_n163 ), .ZN(_add_2_root_add_136_4_n293 ) );
NAND2_X2 _add_2_root_add_136_4_U363  ( .A1(Kt[21]), .A2(SHA1_result[21]),.ZN(_add_2_root_add_136_4_n286 ) );
INV_X4 _add_2_root_add_136_4_U362  ( .A(_add_2_root_add_136_4_n290 ), .ZN(_add_2_root_add_136_4_n289 ) );
NAND2_X2 _add_2_root_add_136_4_U361  ( .A1(_add_2_root_add_136_4_n165 ),.A2(_add_2_root_add_136_4_n163 ), .ZN(_add_2_root_add_136_4_n261 ) );
INV_X4 _add_2_root_add_136_4_U360  ( .A(_add_2_root_add_136_4_n261 ), .ZN(_add_2_root_add_136_4_n285 ) );
INV_X4 _add_2_root_add_136_4_U359  ( .A(Kt[23]), .ZN(_add_2_root_add_136_4_n282 ) );
INV_X4 _add_2_root_add_136_4_U358  ( .A(SHA1_result[23]), .ZN(_add_2_root_add_136_4_n283 ) );
NAND2_X2 _add_2_root_add_136_4_U357  ( .A1(_add_2_root_add_136_4_n282 ),.A2(_add_2_root_add_136_4_n283 ), .ZN(_add_2_root_add_136_4_n164 ) );
NAND2_X2 _add_2_root_add_136_4_U356  ( .A1(Kt[23]), .A2(SHA1_result[23]),.ZN(_add_2_root_add_136_4_n167 ) );
NAND2_X2 _add_2_root_add_136_4_U355  ( .A1(_add_2_root_add_136_4_n164 ),.A2(_add_2_root_add_136_4_n167 ), .ZN(_add_2_root_add_136_4_n281 ) );
INV_X4 _add_2_root_add_136_4_U354  ( .A(_add_2_root_add_136_4_n280 ), .ZN(_add_2_root_add_136_4_n279 ) );
NAND2_X2 _add_2_root_add_136_4_U353  ( .A1(_add_2_root_add_136_4_n277 ),.A2(_add_2_root_add_136_4_n278 ), .ZN(_add_2_root_add_136_4_n275 ) );
NAND2_X2 _add_2_root_add_136_4_U352  ( .A1(_add_2_root_add_136_4_n130 ),.A2(_add_2_root_add_136_4_n122 ), .ZN(_add_2_root_add_136_4_n276 ) );
NOR2_X2 _add_2_root_add_136_4_U351  ( .A1(_add_2_root_add_136_4_n275 ), .A2(_add_2_root_add_136_4_n276 ), .ZN(_add_2_root_add_136_4_n268 ) );
NAND3_X2 _add_2_root_add_136_4_U350  ( .A1(_add_2_root_add_136_4_n242 ),.A2(_add_2_root_add_136_4_n250 ), .A3(_add_2_root_add_136_4_n237 ),.ZN(_add_2_root_add_136_4_n273 ) );
NAND2_X2 _add_2_root_add_136_4_U349  ( .A1(_add_2_root_add_136_4_n123 ),.A2(_add_2_root_add_136_4_n131 ), .ZN(_add_2_root_add_136_4_n272 ) );
NAND2_X2 _add_2_root_add_136_4_U348  ( .A1(_add_2_root_add_136_4_n268 ),.A2(_add_2_root_add_136_4_n269 ), .ZN(_add_2_root_add_136_4_n267 ) );
NAND2_X2 _add_2_root_add_136_4_U347  ( .A1(_add_2_root_add_136_4_n266 ),.A2(_add_2_root_add_136_4_n267 ), .ZN(_add_2_root_add_136_4_n255 ) );
INV_X4 _add_2_root_add_136_4_U346  ( .A(_add_2_root_add_136_4_n265 ), .ZN(_add_2_root_add_136_4_n262 ) );
INV_X4 _add_2_root_add_136_4_U345  ( .A(_add_2_root_add_136_4_n264 ), .ZN(_add_2_root_add_136_4_n263 ) );
NAND2_X2 _add_2_root_add_136_4_U344  ( .A1(_add_2_root_add_136_4_n261 ),.A2(_add_2_root_add_136_4_n167 ), .ZN(_add_2_root_add_136_4_n260 ) );
NAND2_X2 _add_2_root_add_136_4_U343  ( .A1(_add_2_root_add_136_4_n260 ),.A2(_add_2_root_add_136_4_n164 ), .ZN(_add_2_root_add_136_4_n223 ) );
INV_X4 _add_2_root_add_136_4_U342  ( .A(_add_2_root_add_136_4_n223 ), .ZN(_add_2_root_add_136_4_n259 ) );
NAND2_X2 _add_2_root_add_136_4_U341  ( .A1(_add_2_root_add_136_4_n255 ),.A2(_add_2_root_add_136_4_n256 ), .ZN(_add_2_root_add_136_4_n192 ) );
INV_X4 _add_2_root_add_136_4_U340  ( .A(_add_2_root_add_136_4_n192 ), .ZN(_add_2_root_add_136_4_n215 ) );
XNOR2_X2 _add_2_root_add_136_4_U339  ( .A(_add_2_root_add_136_4_n215 ), .B(_add_2_root_add_136_4_n254 ), .ZN(N120) );
INV_X4 _add_2_root_add_136_4_U338  ( .A(_add_2_root_add_136_4_n131 ), .ZN(_add_2_root_add_136_4_n253 ) );
NAND3_X2 _add_2_root_add_136_4_U337  ( .A1(_add_2_root_add_136_4_n242 ),.A2(_add_2_root_add_136_4_n250 ), .A3(_add_2_root_add_136_4_n237 ),.ZN(_add_2_root_add_136_4_n248 ) );
NAND2_X2 _add_2_root_add_136_4_U336  ( .A1(_add_2_root_add_136_4_n34 ), .A2(_add_2_root_add_136_4_n185 ), .ZN(_add_2_root_add_136_4_n249 ) );
NAND3_X2 _add_2_root_add_136_4_U335  ( .A1(_add_2_root_add_136_4_n237 ),.A2(_add_2_root_add_136_4_n242 ), .A3(_add_2_root_add_136_4_n243 ),.ZN(_add_2_root_add_136_4_n227 ) );
NAND2_X2 _add_2_root_add_136_4_U334  ( .A1(_add_2_root_add_136_4_n239 ),.A2(_add_2_root_add_136_4_n240 ), .ZN(_add_2_root_add_136_4_n228 ) );
NAND2_X2 _add_2_root_add_136_4_U333  ( .A1(_add_2_root_add_136_4_n237 ),.A2(_add_2_root_add_136_4_n238 ), .ZN(_add_2_root_add_136_4_n235 ) );
NAND2_X2 _add_2_root_add_136_4_U332  ( .A1(_add_2_root_add_136_4_n223 ),.A2(_add_2_root_add_136_4_n28 ), .ZN(_add_2_root_add_136_4_n221 ) );
XNOR2_X2 _add_2_root_add_136_4_U331  ( .A(_add_2_root_add_136_4_n216 ), .B(_add_2_root_add_136_4_n217 ), .ZN(N121) );
NAND2_X2 _add_2_root_add_136_4_U330  ( .A1(Kt[25]), .A2(SHA1_result[25]),.ZN(_add_2_root_add_136_4_n213 ) );
NAND2_X2 _add_2_root_add_136_4_U329  ( .A1(Kt[24]), .A2(SHA1_result[24]),.ZN(_add_2_root_add_136_4_n214 ) );
NAND2_X2 _add_2_root_add_136_4_U328  ( .A1(_add_2_root_add_136_4_n213 ),.A2(_add_2_root_add_136_4_n214 ), .ZN(_add_2_root_add_136_4_n198 ) );
INV_X4 _add_2_root_add_136_4_U327  ( .A(_add_2_root_add_136_4_n199 ), .ZN(_add_2_root_add_136_4_n207 ) );
INV_X4 _add_2_root_add_136_4_U326  ( .A(Kt[26]), .ZN(_add_2_root_add_136_4_n210 ) );
INV_X4 _add_2_root_add_136_4_U325  ( .A(SHA1_result[26]), .ZN(_add_2_root_add_136_4_n211 ) );
NAND2_X2 _add_2_root_add_136_4_U324  ( .A1(_add_2_root_add_136_4_n210 ),.A2(_add_2_root_add_136_4_n211 ), .ZN(_add_2_root_add_136_4_n197 ) );
NAND2_X2 _add_2_root_add_136_4_U323  ( .A1(Kt[26]), .A2(SHA1_result[26]),.ZN(_add_2_root_add_136_4_n195 ) );
NAND2_X2 _add_2_root_add_136_4_U322  ( .A1(_add_2_root_add_136_4_n197 ),.A2(_add_2_root_add_136_4_n195 ), .ZN(_add_2_root_add_136_4_n209 ) );
NAND2_X2 _add_2_root_add_136_4_U321  ( .A1(_add_2_root_add_136_4_n13 ), .A2(_add_2_root_add_136_4_n197 ), .ZN(_add_2_root_add_136_4_n204 ) );
INV_X4 _add_2_root_add_136_4_U320  ( .A(_add_2_root_add_136_4_n208 ), .ZN(_add_2_root_add_136_4_n206 ) );
NAND2_X2 _add_2_root_add_136_4_U319  ( .A1(_add_2_root_add_136_4_n193 ),.A2(_add_2_root_add_136_4_n192 ), .ZN(_add_2_root_add_136_4_n205 ) );
NAND2_X2 _add_2_root_add_136_4_U318  ( .A1(Kt[27]), .A2(SHA1_result[27]),.ZN(_add_2_root_add_136_4_n194 ) );
INV_X4 _add_2_root_add_136_4_U317  ( .A(Kt[27]), .ZN(_add_2_root_add_136_4_n202 ) );
INV_X4 _add_2_root_add_136_4_U316  ( .A(SHA1_result[27]), .ZN(_add_2_root_add_136_4_n203 ) );
NAND2_X2 _add_2_root_add_136_4_U315  ( .A1(_add_2_root_add_136_4_n202 ),.A2(_add_2_root_add_136_4_n203 ), .ZN(_add_2_root_add_136_4_n170 ) );
NAND2_X2 _add_2_root_add_136_4_U314  ( .A1(_add_2_root_add_136_4_n194 ),.A2(_add_2_root_add_136_4_n170 ), .ZN(_add_2_root_add_136_4_n201 ) );
XNOR2_X2 _add_2_root_add_136_4_U313  ( .A(_add_2_root_add_136_4_n200 ), .B(_add_2_root_add_136_4_n201 ), .ZN(N123) );
NAND2_X2 _add_2_root_add_136_4_U312  ( .A1(_add_2_root_add_136_4_n172 ),.A2(_add_2_root_add_136_4_n170 ), .ZN(_add_2_root_add_136_4_n189 ) );
INV_X4 _add_2_root_add_136_4_U311  ( .A(_add_2_root_add_136_4_n176 ), .ZN(_add_2_root_add_136_4_n193 ) );
NAND2_X2 _add_2_root_add_136_4_U310  ( .A1(_add_2_root_add_136_4_n193 ),.A2(_add_2_root_add_136_4_n170 ), .ZN(_add_2_root_add_136_4_n108 ) );
INV_X4 _add_2_root_add_136_4_U309  ( .A(_add_2_root_add_136_4_n108 ), .ZN(_add_2_root_add_136_4_n191 ) );
NAND2_X2 _add_2_root_add_136_4_U308  ( .A1(_add_2_root_add_136_4_n191 ),.A2(_add_2_root_add_136_4_n192 ), .ZN(_add_2_root_add_136_4_n190 ) );
NAND2_X2 _add_2_root_add_136_4_U307  ( .A1(_add_2_root_add_136_4_n189 ),.A2(_add_2_root_add_136_4_n190 ), .ZN(_add_2_root_add_136_4_n186 ) );
NAND2_X2 _add_2_root_add_136_4_U306  ( .A1(Kt[28]), .A2(SHA1_result[28]),.ZN(_add_2_root_add_136_4_n106 ) );
INV_X4 _add_2_root_add_136_4_U305  ( .A(Kt[28]), .ZN(_add_2_root_add_136_4_n187 ) );
INV_X4 _add_2_root_add_136_4_U304  ( .A(SHA1_result[28]), .ZN(_add_2_root_add_136_4_n188 ) );
NAND2_X2 _add_2_root_add_136_4_U303  ( .A1(_add_2_root_add_136_4_n187 ),.A2(_add_2_root_add_136_4_n188 ), .ZN(_add_2_root_add_136_4_n171 ) );
NAND4_X2 _add_2_root_add_136_4_U302  ( .A1(_add_2_root_add_136_4_n129 ),.A2(_add_2_root_add_136_4_n130 ), .A3(_add_2_root_add_136_4_n131 ),.A4(_add_2_root_add_136_4_n132 ), .ZN(_add_2_root_add_136_4_n180 ) );
INV_X4 _add_2_root_add_136_4_U301  ( .A(_add_2_root_add_136_4_n126 ), .ZN(_add_2_root_add_136_4_n184 ) );
NAND2_X2 _add_2_root_add_136_4_U300  ( .A1(_add_2_root_add_136_4_n122 ),.A2(_add_2_root_add_136_4_n123 ), .ZN(_add_2_root_add_136_4_n182 ) );
NAND2_X2 _add_2_root_add_136_4_U299  ( .A1(_add_2_root_add_136_4_n112 ),.A2(_add_2_root_add_136_4_n116 ), .ZN(_add_2_root_add_136_4_n152 ) );
INV_X4 _add_2_root_add_136_4_U298  ( .A(_add_2_root_add_136_4_n171 ), .ZN(_add_2_root_add_136_4_n100 ) );
INV_X4 _add_2_root_add_136_4_U297  ( .A(_add_2_root_add_136_4_n170 ), .ZN(_add_2_root_add_136_4_n177 ) );
INV_X4 _add_2_root_add_136_4_U296  ( .A(_add_2_root_add_136_4_n105 ), .ZN(_add_2_root_add_136_4_n175 ) );
NAND2_X2 _add_2_root_add_136_4_U295  ( .A1(_add_2_root_add_136_4_n150 ),.A2(_add_2_root_add_136_4_n175 ), .ZN(_add_2_root_add_136_4_n174 ) );
NAND2_X2 _add_2_root_add_136_4_U294  ( .A1(_add_2_root_add_136_4_n107 ),.A2(_add_2_root_add_136_4_n106 ), .ZN(_add_2_root_add_136_4_n169 ) );
INV_X4 _add_2_root_add_136_4_U293  ( .A(_add_2_root_add_136_4_n167 ), .ZN(_add_2_root_add_136_4_n166 ) );
NAND2_X2 _add_2_root_add_136_4_U292  ( .A1(_add_2_root_add_136_4_n161 ),.A2(_add_2_root_add_136_4_n162 ), .ZN(_add_2_root_add_136_4_n157 ) );
NAND2_X2 _add_2_root_add_136_4_U291  ( .A1(Kt[29]), .A2(SHA1_result[29]),.ZN(_add_2_root_add_136_4_n95 ) );
INV_X4 _add_2_root_add_136_4_U290  ( .A(Kt[29]), .ZN(_add_2_root_add_136_4_n159 ) );
INV_X4 _add_2_root_add_136_4_U289  ( .A(SHA1_result[29]), .ZN(_add_2_root_add_136_4_n160 ) );
NAND2_X2 _add_2_root_add_136_4_U288  ( .A1(_add_2_root_add_136_4_n159 ),.A2(_add_2_root_add_136_4_n160 ), .ZN(_add_2_root_add_136_4_n145 ) );
NAND2_X2 _add_2_root_add_136_4_U287  ( .A1(_add_2_root_add_136_4_n95 ), .A2(_add_2_root_add_136_4_n145 ), .ZN(_add_2_root_add_136_4_n158 ) );
XNOR2_X2 _add_2_root_add_136_4_U286  ( .A(_add_2_root_add_136_4_n157 ), .B(_add_2_root_add_136_4_n158 ), .ZN(N125) );
XNOR2_X2 _add_2_root_add_136_4_U285  ( .A(_add_2_root_add_136_4_n87 ), .B(_add_2_root_add_136_4_n154 ), .ZN(N98) );
NAND2_X2 _add_2_root_add_136_4_U284  ( .A1(_add_2_root_add_136_4_n145 ),.A2(_add_2_root_add_136_4_n150 ), .ZN(_add_2_root_add_136_4_n149 ) );
NAND2_X2 _add_2_root_add_136_4_U283  ( .A1(_add_2_root_add_136_4_n104 ),.A2(_add_2_root_add_136_4_n145 ), .ZN(_add_2_root_add_136_4_n140 ) );
NAND2_X2 _add_2_root_add_136_4_U282  ( .A1(_add_2_root_add_136_4_n5 ), .A2(_add_2_root_add_136_4_n145 ), .ZN(_add_2_root_add_136_4_n141 ) );
INV_X4 _add_2_root_add_136_4_U281  ( .A(_add_2_root_add_136_4_n95 ), .ZN(_add_2_root_add_136_4_n146 ) );
INV_X4 _add_2_root_add_136_4_U280  ( .A(_add_2_root_add_136_4_n145 ), .ZN(_add_2_root_add_136_4_n101 ) );
INV_X4 _add_2_root_add_136_4_U279  ( .A(_add_2_root_add_136_4_n107 ), .ZN(_add_2_root_add_136_4_n144 ) );
NAND2_X2 _add_2_root_add_136_4_U278  ( .A1(_add_2_root_add_136_4_n144 ),.A2(_add_2_root_add_136_4_n145 ), .ZN(_add_2_root_add_136_4_n143 ) );
NAND4_X2 _add_2_root_add_136_4_U277  ( .A1(_add_2_root_add_136_4_n140 ),.A2(_add_2_root_add_136_4_n141 ), .A3(_add_2_root_add_136_4_n142 ),.A4(_add_2_root_add_136_4_n143 ), .ZN(_add_2_root_add_136_4_n139 ) );
INV_X4 _add_2_root_add_136_4_U276  ( .A(Kt[30]), .ZN(_add_2_root_add_136_4_n136 ) );
INV_X4 _add_2_root_add_136_4_U275  ( .A(SHA1_result[30]), .ZN(_add_2_root_add_136_4_n137 ) );
NAND2_X2 _add_2_root_add_136_4_U274  ( .A1(_add_2_root_add_136_4_n136 ),.A2(_add_2_root_add_136_4_n137 ), .ZN(_add_2_root_add_136_4_n93 ) );
INV_X4 _add_2_root_add_136_4_U273  ( .A(_add_2_root_add_136_4_n93 ), .ZN(_add_2_root_add_136_4_n102 ) );
NAND2_X2 _add_2_root_add_136_4_U272  ( .A1(Kt[30]), .A2(SHA1_result[30]),.ZN(_add_2_root_add_136_4_n94 ) );
INV_X4 _add_2_root_add_136_4_U271  ( .A(_add_2_root_add_136_4_n94 ), .ZN(_add_2_root_add_136_4_n135 ) );
XNOR2_X2 _add_2_root_add_136_4_U270  ( .A(_add_2_root_add_136_4_n133 ), .B(_add_2_root_add_136_4_n134 ), .ZN(N126) );
NAND4_X2 _add_2_root_add_136_4_U269  ( .A1(_add_2_root_add_136_4_n129 ),.A2(_add_2_root_add_136_4_n130 ), .A3(_add_2_root_add_136_4_n131 ),.A4(_add_2_root_add_136_4_n132 ), .ZN(_add_2_root_add_136_4_n119 ) );
NAND2_X2 _add_2_root_add_136_4_U268  ( .A1(_add_2_root_add_136_4_n122 ),.A2(_add_2_root_add_136_4_n123 ), .ZN(_add_2_root_add_136_4_n121 ) );
INV_X4 _add_2_root_add_136_4_U267  ( .A(_add_2_root_add_136_4_n116 ), .ZN(_add_2_root_add_136_4_n114 ) );
INV_X4 _add_2_root_add_136_4_U266  ( .A(_add_2_root_add_136_4_n106 ), .ZN(_add_2_root_add_136_4_n115 ) );
NAND4_X2 _add_2_root_add_136_4_U265  ( .A1(_add_2_root_add_136_4_n107 ),.A2(_add_2_root_add_136_4_n111 ), .A3(_add_2_root_add_136_4_n112 ),.A4(_add_2_root_add_136_4_n113 ), .ZN(_add_2_root_add_136_4_n110 ) );
NAND2_X2 _add_2_root_add_136_4_U264  ( .A1(_add_2_root_add_136_4_n94 ), .A2(_add_2_root_add_136_4_n95 ), .ZN(_add_2_root_add_136_4_n92 ) );
NAND2_X2 _add_2_root_add_136_4_U263  ( .A1(_add_2_root_add_136_4_n92 ), .A2(_add_2_root_add_136_4_n93 ), .ZN(_add_2_root_add_136_4_n91 ) );
INV_X4 _add_2_root_add_136_4_U262  ( .A(Kt[31]), .ZN(_add_2_root_add_136_4_n90 ) );
XNOR2_X2 _add_2_root_add_136_4_U261  ( .A(_add_2_root_add_136_4_n90 ), .B(SHA1_result[31]), .ZN(_add_2_root_add_136_4_n89 ) );
XNOR2_X2 _add_2_root_add_136_4_U260  ( .A(_add_2_root_add_136_4_n88 ), .B(_add_2_root_add_136_4_n89 ), .ZN(N127) );
XNOR2_X2 _add_2_root_add_136_4_U259  ( .A(_add_2_root_add_136_4_n81 ), .B(_add_2_root_add_136_4_n82 ), .ZN(N99) );
INV_X4 _add_2_root_add_136_4_U258  ( .A(_add_2_root_add_136_4_n68 ), .ZN(_add_2_root_add_136_4_n75 ) );
XNOR2_X2 _add_2_root_add_136_4_U257  ( .A(_add_2_root_add_136_4_n53 ), .B(_add_2_root_add_136_4_n80 ), .ZN(N100) );
INV_X4 _add_2_root_add_136_4_U256  ( .A(_add_2_root_add_136_4_n69 ), .ZN(_add_2_root_add_136_4_n72 ) );
XNOR2_X2 _add_2_root_add_136_4_U255  ( .A(_add_2_root_add_136_4_n77 ), .B(_add_2_root_add_136_4_n78 ), .ZN(N101) );
XNOR2_X2 _add_2_root_add_136_4_U254  ( .A(_add_2_root_add_136_4_n70 ), .B(_add_2_root_add_136_4_n71 ), .ZN(N102) );
NAND2_X2 _add_2_root_add_136_4_U253  ( .A1(_add_2_root_add_136_4_n68 ), .A2(_add_2_root_add_136_4_n69 ), .ZN(_add_2_root_add_136_4_n67 ) );
INV_X4 _add_2_root_add_136_4_U252  ( .A(_add_2_root_add_136_4_n62 ), .ZN(_add_2_root_add_136_4_n60 ) );
XNOR2_X2 _add_2_root_add_136_4_U251  ( .A(_add_2_root_add_136_4_n58 ), .B(_add_2_root_add_136_4_n59 ), .ZN(N103) );
XNOR2_X2 _add_2_root_add_136_4_U250  ( .A(_add_2_root_add_136_4_n55 ), .B(_add_2_root_add_136_4_n56 ), .ZN(N104) );
XNOR2_X2 _add_2_root_add_136_4_U249  ( .A(_add_2_root_add_136_4_n44 ), .B(_add_2_root_add_136_4_n45 ), .ZN(N105) );
NAND2_X2 _add_2_root_add_136_4_U248  ( .A1(_add_2_root_add_136_4_n245 ),.A2(_add_2_root_add_136_4_n246 ), .ZN(_add_2_root_add_136_4_n225 ) );
OR2_X2 _add_2_root_add_136_4_U247  ( .A1(SHA1_result[16]), .A2(Kt[16]), .ZN(_add_2_root_add_136_4_n43 ) );
OR2_X2 _add_2_root_add_136_4_U246  ( .A1(SHA1_result[15]), .A2(Kt[15]), .ZN(_add_2_root_add_136_4_n42 ) );
AND2_X2 _add_2_root_add_136_4_U245  ( .A1(SHA1_result[8]), .A2(Kt[8]), .ZN(_add_2_root_add_136_4_n407 ) );
NOR2_X2 _add_2_root_add_136_4_U244  ( .A1(SHA1_result[9]), .A2(Kt[9]), .ZN(_add_2_root_add_136_4_n410 ) );
NOR2_X2 _add_2_root_add_136_4_U243  ( .A1(_add_2_root_add_136_4_n409 ), .A2(_add_2_root_add_136_4_n410 ), .ZN(_add_2_root_add_136_4_n408 ) );
AND2_X2 _add_2_root_add_136_4_U242  ( .A1(Kt[2]), .A2(SHA1_result[2]), .ZN(_add_2_root_add_136_4_n40 ) );
NOR2_X2 _add_2_root_add_136_4_U241  ( .A1(_add_2_root_add_136_4_n336 ), .A2(_add_2_root_add_136_4_n337 ), .ZN(_add_2_root_add_136_4_n335 ) );
AND3_X4 _add_2_root_add_136_4_U240  ( .A1(SHA1_result[17]), .A2(Kt[17]),.A3(SHA1_result[18]), .ZN(_add_2_root_add_136_4_n39 ) );
OR2_X2 _add_2_root_add_136_4_U239  ( .A1(_add_2_root_add_136_4_n335 ), .A2(_add_2_root_add_136_4_n39 ), .ZN(_add_2_root_add_136_4_n264 ) );
NOR2_X2 _add_2_root_add_136_4_U238  ( .A1(_add_2_root_add_136_4_n406 ), .A2(_add_2_root_add_136_4_n22 ), .ZN(_add_2_root_add_136_4_n405 ) );
NAND3_X2 _add_2_root_add_136_4_U237  ( .A1(SHA1_result[9]), .A2(_add_2_root_add_136_4_n41 ), .A3(Kt[9]), .ZN(_add_2_root_add_136_4_n404 ) );
NAND3_X2 _add_2_root_add_136_4_U236  ( .A1(_add_2_root_add_136_4_n403 ),.A2(_add_2_root_add_136_4_n404 ), .A3(_add_2_root_add_136_4_n405 ),.ZN(_add_2_root_add_136_4_n363 ) );
NAND3_X2 _add_2_root_add_136_4_U235  ( .A1(SHA1_result[20]), .A2(Kt[20]),.A3(_add_2_root_add_136_4_n289 ), .ZN(_add_2_root_add_136_4_n288 ) );
NAND3_X2 _add_2_root_add_136_4_U234  ( .A1(_add_2_root_add_136_4_n286 ),.A2(_add_2_root_add_136_4_n287 ), .A3(_add_2_root_add_136_4_n288 ),.ZN(_add_2_root_add_136_4_n165 ) );
NOR2_X2 _add_2_root_add_136_4_U233  ( .A1(SHA1_result[5]), .A2(Kt[5]), .ZN(_add_2_root_add_136_4_n431 ) );
NOR2_X2 _add_2_root_add_136_4_U232  ( .A1(SHA1_result[8]), .A2(Kt[8]), .ZN(_add_2_root_add_136_4_n413 ) );
NOR2_X2 _add_2_root_add_136_4_U231  ( .A1(SHA1_result[6]), .A2(Kt[6]), .ZN(_add_2_root_add_136_4_n432 ) );
NOR2_X2 _add_2_root_add_136_4_U230  ( .A1(SHA1_result[10]), .A2(Kt[10]),.ZN(_add_2_root_add_136_4_n412 ) );
NOR2_X2 _add_2_root_add_136_4_U229  ( .A1(SHA1_result[12]), .A2(Kt[12]),.ZN(_add_2_root_add_136_4_n378 ) );
NOR2_X2 _add_2_root_add_136_4_U228  ( .A1(SHA1_result[14]), .A2(Kt[14]),.ZN(_add_2_root_add_136_4_n377 ) );
NOR2_X2 _add_2_root_add_136_4_U227  ( .A1(_add_2_root_add_136_4_n377 ), .A2(_add_2_root_add_136_4_n378 ), .ZN(_add_2_root_add_136_4_n376 ) );
NAND3_X2 _add_2_root_add_136_4_U226  ( .A1(Kt[16]), .A2(SHA1_result[16]),.A3(SHA1_result[18]), .ZN(_add_2_root_add_136_4_n337 ) );
NAND3_X2 _add_2_root_add_136_4_U225  ( .A1(SHA1_result[2]), .A2(Kt[2]), .A3(_add_2_root_add_136_4_n353 ), .ZN(_add_2_root_add_136_4_n244 ) );
NAND3_X2 _add_2_root_add_136_4_U224  ( .A1(SHA1_result[16]), .A2(Kt[16]),.A3(_add_2_root_add_136_4_n342 ), .ZN(_add_2_root_add_136_4_n339 ) );
NOR2_X2 _add_2_root_add_136_4_U223  ( .A1(SHA1_result[15]), .A2(Kt[15]),.ZN(_add_2_root_add_136_4_n369 ) );
NOR2_X2 _add_2_root_add_136_4_U222  ( .A1(SHA1_result[21]), .A2(Kt[21]),.ZN(_add_2_root_add_136_4_n292 ) );
NOR2_X2 _add_2_root_add_136_4_U221  ( .A1(SHA1_result[17]), .A2(Kt[17]),.ZN(_add_2_root_add_136_4_n336 ) );
NOR2_X2 _add_2_root_add_136_4_U220  ( .A1(SHA1_result[17]), .A2(Kt[17]),.ZN(_add_2_root_add_136_4_n333 ) );
NOR2_X2 _add_2_root_add_136_4_U219  ( .A1(SHA1_result[16]), .A2(Kt[16]),.ZN(_add_2_root_add_136_4_n334 ) );
NAND3_X2 _add_2_root_add_136_4_U218  ( .A1(SHA1_result[6]), .A2(Kt[6]), .A3(_add_2_root_add_136_4_n374 ), .ZN(_add_2_root_add_136_4_n234 ) );
OR2_X4 _add_2_root_add_136_4_U217  ( .A1(SHA1_result[0]), .A2(Kt[0]), .ZN(_add_2_root_add_136_4_n38 ) );
AND2_X2 _add_2_root_add_136_4_U216  ( .A1(_add_2_root_add_136_4_n327 ), .A2(_add_2_root_add_136_4_n38 ), .ZN(N96) );
NOR2_X2 _add_2_root_add_136_4_U215  ( .A1(SHA1_result[21]), .A2(Kt[21]),.ZN(_add_2_root_add_136_4_n290 ) );
NOR2_X2 _add_2_root_add_136_4_U214  ( .A1(SHA1_result[1]), .A2(Kt[1]), .ZN(_add_2_root_add_136_4_n155 ) );
NOR2_X2 _add_2_root_add_136_4_U213  ( .A1(SHA1_result[4]), .A2(Kt[4]), .ZN(_add_2_root_add_136_4_n76 ) );
NOR2_X2 _add_2_root_add_136_4_U212  ( .A1(SHA1_result[9]), .A2(Kt[9]), .ZN(_add_2_root_add_136_4_n47 ) );
NOR2_X2 _add_2_root_add_136_4_U211  ( .A1(SHA1_result[13]), .A2(Kt[13]),.ZN(_add_2_root_add_136_4_n385 ) );
NOR2_X2 _add_2_root_add_136_4_U210  ( .A1(SHA1_result[25]), .A2(Kt[25]),.ZN(_add_2_root_add_136_4_n199 ) );
NOR2_X2 _add_2_root_add_136_4_U209  ( .A1(SHA1_result[7]), .A2(Kt[7]), .ZN(_add_2_root_add_136_4_n61 ) );
NOR2_X2 _add_2_root_add_136_4_U208  ( .A1(SHA1_result[2]), .A2(Kt[2]), .ZN(_add_2_root_add_136_4_n86 ) );
NOR2_X2 _add_2_root_add_136_4_U207  ( .A1(SHA1_result[24]), .A2(Kt[24]),.ZN(_add_2_root_add_136_4_n208 ) );
NOR2_X2 _add_2_root_add_136_4_U206  ( .A1(SHA1_result[6]), .A2(Kt[6]), .ZN(_add_2_root_add_136_4_n65 ) );
NOR2_X2 _add_2_root_add_136_4_U205  ( .A1(SHA1_result[14]), .A2(Kt[14]),.ZN(_add_2_root_add_136_4_n368 ) );
NOR2_X2 _add_2_root_add_136_4_U204  ( .A1(SHA1_result[20]), .A2(Kt[20]),.ZN(_add_2_root_add_136_4_n294 ) );
NOR2_X2 _add_2_root_add_136_4_U203  ( .A1(SHA1_result[12]), .A2(Kt[12]),.ZN(_add_2_root_add_136_4_n384 ) );
NOR2_X2 _add_2_root_add_136_4_U202  ( .A1(SHA1_result[5]), .A2(Kt[5]), .ZN(_add_2_root_add_136_4_n64 ) );
OR2_X2 _add_2_root_add_136_4_U201  ( .A1(Kt[3]), .A2(SHA1_result[3]), .ZN(_add_2_root_add_136_4_n353 ) );
OR2_X2 _add_2_root_add_136_4_U200  ( .A1(_add_2_root_add_136_4_n384 ), .A2(_add_2_root_add_136_4_n24 ), .ZN(_add_2_root_add_136_4_n37 ) );
OR2_X2 _add_2_root_add_136_4_U199  ( .A1(_add_2_root_add_136_4_n368 ), .A2(_add_2_root_add_136_4_n370 ), .ZN(_add_2_root_add_136_4_n36 ) );
NAND2_X2 _add_2_root_add_136_4_U198  ( .A1(_add_2_root_add_136_4_n279 ),.A2(_add_2_root_add_136_4_n164 ), .ZN(_add_2_root_add_136_4_n105 ) );
OR2_X2 _add_2_root_add_136_4_U197  ( .A1(_add_2_root_add_136_4_n49 ), .A2(_add_2_root_add_136_4_n47 ), .ZN(_add_2_root_add_136_4_n35 ) );
NAND3_X2 _add_2_root_add_136_4_U196  ( .A1(_add_2_root_add_136_4_n108 ),.A2(_add_2_root_add_136_4_n106 ), .A3(_add_2_root_add_136_4_n107 ),.ZN(_add_2_root_add_136_4_n98 ) );
NOR3_X2 _add_2_root_add_136_4_U195  ( .A1(_add_2_root_add_136_4_n100 ), .A2(_add_2_root_add_136_4_n101 ), .A3(_add_2_root_add_136_4_n102 ), .ZN(_add_2_root_add_136_4_n99 ) );
NAND3_X2 _add_2_root_add_136_4_U194  ( .A1(_add_2_root_add_136_4_n98 ), .A2(_add_2_root_add_136_4_n16 ), .A3(_add_2_root_add_136_4_n99 ), .ZN(_add_2_root_add_136_4_n97 ) );
NOR2_X2 _add_2_root_add_136_4_U193  ( .A1(_add_2_root_add_136_4_n173 ), .A2(_add_2_root_add_136_4_n174 ), .ZN(_add_2_root_add_136_4_n168 ) );
NOR2_X2 _add_2_root_add_136_4_U192  ( .A1(_add_2_root_add_136_4_n168 ), .A2(_add_2_root_add_136_4_n169 ), .ZN(_add_2_root_add_136_4_n161 ) );
AND3_X2 _add_2_root_add_136_4_U191  ( .A1(_add_2_root_add_136_4_n352 ), .A2(_add_2_root_add_136_4_n353 ), .A3(_add_2_root_add_136_4_n354 ), .ZN(_add_2_root_add_136_4_n34 ) );
OR2_X4 _add_2_root_add_136_4_U190  ( .A1(_add_2_root_add_136_4_n96 ), .A2(_add_2_root_add_136_4_n97 ), .ZN(_add_2_root_add_136_4_n33 ) );
AND2_X2 _add_2_root_add_136_4_U189  ( .A1(_add_2_root_add_136_4_n33 ), .A2(_add_2_root_add_136_4_n91 ), .ZN(_add_2_root_add_136_4_n88 ) );
NOR2_X2 _add_2_root_add_136_4_U188  ( .A1(_add_2_root_add_136_4_n416 ), .A2(_add_2_root_add_136_4_n417 ), .ZN(_add_2_root_add_136_4_n414 ) );
NOR2_X2 _add_2_root_add_136_4_U187  ( .A1(_add_2_root_add_136_4_n402 ), .A2(_add_2_root_add_136_4_n22 ), .ZN(_add_2_root_add_136_4_n415 ) );
NOR2_X2 _add_2_root_add_136_4_U186  ( .A1(_add_2_root_add_136_4_n218 ), .A2(_add_2_root_add_136_4_n8 ), .ZN(_add_2_root_add_136_4_n216 ) );
NOR2_X2 _add_2_root_add_136_4_U185  ( .A1(_add_2_root_add_136_4_n199 ), .A2(_add_2_root_add_136_4_n15 ), .ZN(_add_2_root_add_136_4_n217 ) );
NOR2_X2 _add_2_root_add_136_4_U184  ( .A1(_add_2_root_add_136_4_n326 ), .A2(_add_2_root_add_136_4_n155 ), .ZN(_add_2_root_add_136_4_n325 ) );
OR2_X4 _add_2_root_add_136_4_U183  ( .A1(_add_2_root_add_136_4_n212 ), .A2(_add_2_root_add_136_4_n13 ), .ZN(_add_2_root_add_136_4_n32 ) );
XNOR2_X2 _add_2_root_add_136_4_U182  ( .A(_add_2_root_add_136_4_n32 ), .B(_add_2_root_add_136_4_n209 ), .ZN(N122) );
NAND3_X2 _add_2_root_add_136_4_U181  ( .A1(_add_2_root_add_136_4_n373 ),.A2(_add_2_root_add_136_4_n374 ), .A3(_add_2_root_add_136_4_n375 ),.ZN(_add_2_root_add_136_4_n236 ) );
NAND3_X2 _add_2_root_add_136_4_U180  ( .A1(_add_2_root_add_136_4_n434 ),.A2(_add_2_root_add_136_4_n354 ), .A3(_add_2_root_add_136_4_n435 ),.ZN(_add_2_root_add_136_4_n433 ) );
NAND3_X2 _add_2_root_add_136_4_U179  ( .A1(_add_2_root_add_136_4_n244 ),.A2(_add_2_root_add_136_4_n433 ), .A3(_add_2_root_add_136_4_n241 ),.ZN(_add_2_root_add_136_4_n394 ) );
OR2_X2 _add_2_root_add_136_4_U178  ( .A1(_add_2_root_add_136_4_n419 ), .A2(_add_2_root_add_136_4_n420 ), .ZN(_add_2_root_add_136_4_n31 ) );
NOR2_X2 _add_2_root_add_136_4_U177  ( .A1(_add_2_root_add_136_4_n421 ), .A2(_add_2_root_add_136_4_n9 ), .ZN(_add_2_root_add_136_4_n416 ) );
NOR2_X2 _add_2_root_add_136_4_U176  ( .A1(_add_2_root_add_136_4_n383 ), .A2(_add_2_root_add_136_4_n14 ), .ZN(_add_2_root_add_136_4_n381 ) );
OR2_X4 _add_2_root_add_136_4_U175  ( .A1(_add_2_root_add_136_4_n155 ), .A2(_add_2_root_add_136_4_n436 ), .ZN(_add_2_root_add_136_4_n30 ) );
AND2_X2 _add_2_root_add_136_4_U174  ( .A1(_add_2_root_add_136_4_n156 ), .A2(_add_2_root_add_136_4_n30 ), .ZN(_add_2_root_add_136_4_n87 ) );
NOR2_X2 _add_2_root_add_136_4_U173  ( .A1(_add_2_root_add_136_4_n105 ), .A2(_add_2_root_add_136_4_n112 ), .ZN(_add_2_root_add_136_4_n222 ) );
NOR3_X2 _add_2_root_add_136_4_U172  ( .A1(_add_2_root_add_136_4_n220 ), .A2(_add_2_root_add_136_4_n221 ), .A3(_add_2_root_add_136_4_n222 ), .ZN(_add_2_root_add_136_4_n219 ) );
NOR2_X2 _add_2_root_add_136_4_U171  ( .A1(_add_2_root_add_136_4_n208 ), .A2(_add_2_root_add_136_4_n219 ), .ZN(_add_2_root_add_136_4_n218 ) );
NOR3_X2 _add_2_root_add_136_4_U170  ( .A1(_add_2_root_add_136_4_n180 ), .A2(_add_2_root_add_136_4_n181 ), .A3(_add_2_root_add_136_4_n182 ), .ZN(_add_2_root_add_136_4_n179 ) );
NOR2_X2 _add_2_root_add_136_4_U169  ( .A1(_add_2_root_add_136_4_n179 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n178 ) );
NOR2_X2 _add_2_root_add_136_4_U168  ( .A1(_add_2_root_add_136_4_n178 ), .A2(_add_2_root_add_136_4_n152 ), .ZN(_add_2_root_add_136_4_n173 ) );
NOR2_X2 _add_2_root_add_136_4_U167  ( .A1(_add_2_root_add_136_4_n86 ), .A2(_add_2_root_add_136_4_n87 ), .ZN(_add_2_root_add_136_4_n85 ) );
NOR2_X2 _add_2_root_add_136_4_U166  ( .A1(_add_2_root_add_136_4_n85 ), .A2(_add_2_root_add_136_4_n40 ), .ZN(_add_2_root_add_136_4_n81 ) );
NOR2_X2 _add_2_root_add_136_4_U165  ( .A1(_add_2_root_add_136_4_n83 ), .A2(_add_2_root_add_136_4_n84 ), .ZN(_add_2_root_add_136_4_n82 ) );
NOR3_X2 _add_2_root_add_136_4_U164  ( .A1(_add_2_root_add_136_4_n317 ), .A2(_add_2_root_add_136_4_n318 ), .A3(_add_2_root_add_136_4_n319 ), .ZN(_add_2_root_add_136_4_n316 ) );
NOR2_X2 _add_2_root_add_136_4_U163  ( .A1(_add_2_root_add_136_4_n316 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n315 ) );
NOR2_X2 _add_2_root_add_136_4_U162  ( .A1(_add_2_root_add_136_4_n315 ), .A2(_add_2_root_add_136_4_n296 ), .ZN(_add_2_root_add_136_4_n314 ) );
NOR2_X2 _add_2_root_add_136_4_U161  ( .A1(_add_2_root_add_136_4_n294 ), .A2(_add_2_root_add_136_4_n314 ), .ZN(_add_2_root_add_136_4_n313 ) );
AND3_X4 _add_2_root_add_136_4_U160  ( .A1(_add_2_root_add_136_4_n163 ), .A2(_add_2_root_add_136_4_n164 ), .A3(_add_2_root_add_136_4_n165 ), .ZN(_add_2_root_add_136_4_n29 ) );
AND2_X2 _add_2_root_add_136_4_U159  ( .A1(_add_2_root_add_136_4_n150 ), .A2(_add_2_root_add_136_4_n29 ), .ZN(_add_2_root_add_136_4_n104 ) );
OR2_X2 _add_2_root_add_136_4_U158  ( .A1(_add_2_root_add_136_4_n105 ), .A2(_add_2_root_add_136_4_n116 ), .ZN(_add_2_root_add_136_4_n28 ) );
NAND3_X2 _add_2_root_add_136_4_U157  ( .A1(_add_2_root_add_136_4_n207 ),.A2(_add_2_root_add_136_4_n197 ), .A3(_add_2_root_add_136_4_n198 ),.ZN(_add_2_root_add_136_4_n196 ) );
NAND3_X2 _add_2_root_add_136_4_U156  ( .A1(_add_2_root_add_136_4_n194 ),.A2(_add_2_root_add_136_4_n195 ), .A3(_add_2_root_add_136_4_n196 ),.ZN(_add_2_root_add_136_4_n172 ) );
NOR2_X2 _add_2_root_add_136_4_U155  ( .A1(_add_2_root_add_136_4_n53 ), .A2(_add_2_root_add_136_4_n54 ), .ZN(_add_2_root_add_136_4_n425 ) );
NOR3_X2 _add_2_root_add_136_4_U154  ( .A1(_add_2_root_add_136_4_n425 ), .A2(_add_2_root_add_136_4_n2 ), .A3(_add_2_root_add_136_4_n52 ), .ZN(_add_2_root_add_136_4_n421 ) );
NOR2_X2 _add_2_root_add_136_4_U153  ( .A1(_add_2_root_add_136_4_n101 ), .A2(_add_2_root_add_136_4_n106 ), .ZN(_add_2_root_add_136_4_n147 ) );
NAND3_X2 _add_2_root_add_136_4_U152  ( .A1(_add_2_root_add_136_4_n105 ),.A2(_add_2_root_add_136_4_n106 ), .A3(_add_2_root_add_136_4_n107 ),.ZN(_add_2_root_add_136_4_n103 ) );
NOR2_X2 _add_2_root_add_136_4_U151  ( .A1(_add_2_root_add_136_4_n105 ), .A2(_add_2_root_add_136_4_n116 ), .ZN(_add_2_root_add_136_4_n258 ) );
NAND3_X2 _add_2_root_add_136_4_U150  ( .A1(_add_2_root_add_136_4_n184 ),.A2(_add_2_root_add_136_4_n125 ), .A3(_add_2_root_add_136_4_n124 ),.ZN(_add_2_root_add_136_4_n120 ) );
NOR3_X2 _add_2_root_add_136_4_U149  ( .A1(_add_2_root_add_136_4_n119 ), .A2(_add_2_root_add_136_4_n120 ), .A3(_add_2_root_add_136_4_n121 ), .ZN(_add_2_root_add_136_4_n117 ) );
NOR2_X2 _add_2_root_add_136_4_U148  ( .A1(_add_2_root_add_136_4_n84 ), .A2(_add_2_root_add_136_4_n86 ), .ZN(_add_2_root_add_136_4_n435 ) );
NAND3_X2 _add_2_root_add_136_4_U147  ( .A1(_add_2_root_add_136_4_n206 ),.A2(_add_2_root_add_136_4_n197 ), .A3(_add_2_root_add_136_4_n207 ),.ZN(_add_2_root_add_136_4_n176 ) );
NOR3_X2 _add_2_root_add_136_4_U146  ( .A1(_add_2_root_add_136_4_n390 ), .A2(_add_2_root_add_136_4_n11 ), .A3(_add_2_root_add_136_4_n391 ), .ZN(_add_2_root_add_136_4_n383 ) );
NOR3_X2 _add_2_root_add_136_4_U145  ( .A1(_add_2_root_add_136_4_n215 ), .A2(_add_2_root_add_136_4_n199 ), .A3(_add_2_root_add_136_4_n208 ), .ZN(_add_2_root_add_136_4_n212 ) );
NOR3_X2 _add_2_root_add_136_4_U144  ( .A1(_add_2_root_add_136_4_n383 ), .A2(_add_2_root_add_136_4_n385 ), .A3(_add_2_root_add_136_4_n384 ), .ZN(_add_2_root_add_136_4_n389 ) );
NAND3_X2 _add_2_root_add_136_4_U143  ( .A1(_add_2_root_add_136_4_n237 ),.A2(_add_2_root_add_136_4_n362 ), .A3(_add_2_root_add_136_4_n363 ),.ZN(_add_2_root_add_136_4_n129 ) );
NOR2_X2 _add_2_root_add_136_4_U142  ( .A1(_add_2_root_add_136_4_n151 ), .A2(_add_2_root_add_136_4_n152 ), .ZN(_add_2_root_add_136_4_n148 ) );
NOR3_X2 _add_2_root_add_136_4_U141  ( .A1(_add_2_root_add_136_4_n148 ), .A2(_add_2_root_add_136_4_n105 ), .A3(_add_2_root_add_136_4_n149 ), .ZN(_add_2_root_add_136_4_n138 ) );
NOR2_X2 _add_2_root_add_136_4_U140  ( .A1(_add_2_root_add_136_4_n294 ), .A2(_add_2_root_add_136_4_n292 ), .ZN(_add_2_root_add_136_4_n305 ) );
NOR2_X2 _add_2_root_add_136_4_U139  ( .A1(_add_2_root_add_136_4_n53 ), .A2(_add_2_root_add_136_4_n76 ), .ZN(_add_2_root_add_136_4_n66 ) );
NOR3_X2 _add_2_root_add_136_4_U138  ( .A1(_add_2_root_add_136_4_n105 ), .A2(_add_2_root_add_136_4_n262 ), .A3(_add_2_root_add_136_4_n263 ), .ZN(_add_2_root_add_136_4_n257 ) );
NOR3_X2 _add_2_root_add_136_4_U137  ( .A1(_add_2_root_add_136_4_n333 ), .A2(_add_2_root_add_136_4_n338 ), .A3(_add_2_root_add_136_4_n334 ), .ZN(_add_2_root_add_136_4_n324 ) );
OR2_X4 _add_2_root_add_136_4_U136  ( .A1(_add_2_root_add_136_4_n293 ), .A2(_add_2_root_add_136_4_n294 ), .ZN(_add_2_root_add_136_4_n26 ) );
OR2_X2 _add_2_root_add_136_4_U135  ( .A1(_add_2_root_add_136_4_n26 ), .A2(_add_2_root_add_136_4_n292 ), .ZN(_add_2_root_add_136_4_n280 ) );
NAND3_X2 _add_2_root_add_136_4_U134  ( .A1(_add_2_root_add_136_4_n170 ),.A2(_add_2_root_add_136_4_n171 ), .A3(_add_2_root_add_136_4_n172 ),.ZN(_add_2_root_add_136_4_n107 ) );
NOR3_X2 _add_2_root_add_136_4_U133  ( .A1(_add_2_root_add_136_4_n61 ), .A2(_add_2_root_add_136_4_n64 ), .A3(_add_2_root_add_136_4_n65 ), .ZN(_add_2_root_add_136_4_n427 ) );
NAND3_X2 _add_2_root_add_136_4_U132  ( .A1(_add_2_root_add_136_4_n62 ), .A2(_add_2_root_add_136_4_n426 ), .A3(_add_2_root_add_136_4_n234 ), .ZN(_add_2_root_add_136_4_n52 ) );
NOR2_X2 _add_2_root_add_136_4_U131  ( .A1(_add_2_root_add_136_4_n146 ), .A2(_add_2_root_add_136_4_n147 ), .ZN(_add_2_root_add_136_4_n142 ) );
NOR2_X2 _add_2_root_add_136_4_U130  ( .A1(_add_2_root_add_136_4_n431 ), .A2(_add_2_root_add_136_4_n432 ), .ZN(_add_2_root_add_136_4_n430 ) );
NAND3_X2 _add_2_root_add_136_4_U129  ( .A1(_add_2_root_add_136_4_n4 ), .A2(_add_2_root_add_136_4_n374 ), .A3(_add_2_root_add_136_4_n430 ), .ZN(_add_2_root_add_136_4_n54 ) );
XNOR2_X2 _add_2_root_add_136_4_U128  ( .A(_add_2_root_add_136_4_n25 ), .B(_add_2_root_add_136_4_n281 ), .ZN(N119) );
NOR2_X2 _add_2_root_add_136_4_U127  ( .A1(_add_2_root_add_136_4_n381 ), .A2(_add_2_root_add_136_4_n382 ), .ZN(_add_2_root_add_136_4_n379 ) );
NOR2_X2 _add_2_root_add_136_4_U126  ( .A1(_add_2_root_add_136_4_n369 ), .A2(_add_2_root_add_136_4_n252 ), .ZN(_add_2_root_add_136_4_n380 ) );
NOR2_X2 _add_2_root_add_136_4_U125  ( .A1(_add_2_root_add_136_4_n313 ), .A2(_add_2_root_add_136_4_n7 ), .ZN(_add_2_root_add_136_4_n310 ) );
NOR2_X2 _add_2_root_add_136_4_U124  ( .A1(_add_2_root_add_136_4_n290 ), .A2(_add_2_root_add_136_4_n312 ), .ZN(_add_2_root_add_136_4_n311 ) );
NOR3_X2 _add_2_root_add_136_4_U123  ( .A1(_add_2_root_add_136_4_n176 ), .A2(_add_2_root_add_136_4_n100 ), .A3(_add_2_root_add_136_4_n177 ), .ZN(_add_2_root_add_136_4_n150 ) );
NAND3_X2 _add_2_root_add_136_4_U122  ( .A1(_add_2_root_add_136_4_n301 ),.A2(_add_2_root_add_136_4_n302 ), .A3(_add_2_root_add_136_4_n303 ),.ZN(_add_2_root_add_136_4_n297 ) );
NOR2_X2 _add_2_root_add_136_4_U121  ( .A1(_add_2_root_add_136_4_n398 ), .A2(_add_2_root_add_136_4_n389 ), .ZN(_add_2_root_add_136_4_n386 ) );
NOR2_X2 _add_2_root_add_136_4_U120  ( .A1(_add_2_root_add_136_4_n368 ), .A2(_add_2_root_add_136_4_n388 ), .ZN(_add_2_root_add_136_4_n387 ) );
NOR2_X2 _add_2_root_add_136_4_U119  ( .A1(_add_2_root_add_136_4_n138 ), .A2(_add_2_root_add_136_4_n139 ), .ZN(_add_2_root_add_136_4_n133 ) );
NOR2_X2 _add_2_root_add_136_4_U118  ( .A1(_add_2_root_add_136_4_n102 ), .A2(_add_2_root_add_136_4_n135 ), .ZN(_add_2_root_add_136_4_n134 ) );
NOR2_X2 _add_2_root_add_136_4_U117  ( .A1(_add_2_root_add_136_4_n208 ), .A2(_add_2_root_add_136_4_n8 ), .ZN(_add_2_root_add_136_4_n254 ) );
NOR2_X2 _add_2_root_add_136_4_U116  ( .A1(_add_2_root_add_136_4_n5 ), .A2(_add_2_root_add_136_4_n104 ), .ZN(_add_2_root_add_136_4_n162 ) );
NOR2_X2 _add_2_root_add_136_4_U115  ( .A1(_add_2_root_add_136_4_n360 ), .A2(_add_2_root_add_136_4_n384 ), .ZN(_add_2_root_add_136_4_n399 ) );
NOR2_X2 _add_2_root_add_136_4_U114  ( .A1(_add_2_root_add_136_4_n63 ), .A2(_add_2_root_add_136_4_n6 ), .ZN(_add_2_root_add_136_4_n58 ) );
NOR2_X2 _add_2_root_add_136_4_U113  ( .A1(_add_2_root_add_136_4_n60 ), .A2(_add_2_root_add_136_4_n61 ), .ZN(_add_2_root_add_136_4_n59 ) );
NAND3_X2 _add_2_root_add_136_4_U112  ( .A1(_add_2_root_add_136_4_n204 ),.A2(_add_2_root_add_136_4_n195 ), .A3(_add_2_root_add_136_4_n205 ),.ZN(_add_2_root_add_136_4_n200 ) );
NOR2_X2 _add_2_root_add_136_4_U111  ( .A1(_add_2_root_add_136_4_n323 ), .A2(_add_2_root_add_136_4_n296 ), .ZN(_add_2_root_add_136_4_n321 ) );
NOR2_X2 _add_2_root_add_136_4_U110  ( .A1(_add_2_root_add_136_4_n294 ), .A2(_add_2_root_add_136_4_n7 ), .ZN(_add_2_root_add_136_4_n322 ) );
NOR2_X2 _add_2_root_add_136_4_U109  ( .A1(_add_2_root_add_136_4_n1 ), .A2(_add_2_root_add_136_4_n62 ), .ZN(_add_2_root_add_136_4_n361 ) );
NOR2_X2 _add_2_root_add_136_4_U108  ( .A1(_add_2_root_add_136_4_n412 ), .A2(_add_2_root_add_136_4_n413 ), .ZN(_add_2_root_add_136_4_n411 ) );
NAND3_X2 _add_2_root_add_136_4_U107  ( .A1(_add_2_root_add_136_4_n362 ),.A2(_add_2_root_add_136_4_n3 ), .A3(_add_2_root_add_136_4_n411 ), .ZN(_add_2_root_add_136_4_n233 ) );
NOR2_X2 _add_2_root_add_136_4_U106  ( .A1(_add_2_root_add_136_4_n53 ), .A2(_add_2_root_add_136_4_n54 ), .ZN(_add_2_root_add_136_4_n57 ) );
NOR2_X2 _add_2_root_add_136_4_U105  ( .A1(_add_2_root_add_136_4_n57 ), .A2(_add_2_root_add_136_4_n52 ), .ZN(_add_2_root_add_136_4_n55 ) );
NOR2_X2 _add_2_root_add_136_4_U104  ( .A1(_add_2_root_add_136_4_n49 ), .A2(_add_2_root_add_136_4_n2 ), .ZN(_add_2_root_add_136_4_n56 ) );
NOR2_X2 _add_2_root_add_136_4_U103  ( .A1(_add_2_root_add_136_4_n49 ), .A2(_add_2_root_add_136_4_n50 ), .ZN(_add_2_root_add_136_4_n48 ) );
NOR2_X2 _add_2_root_add_136_4_U102  ( .A1(_add_2_root_add_136_4_n2 ), .A2(_add_2_root_add_136_4_n48 ), .ZN(_add_2_root_add_136_4_n44 ) );
NOR2_X2 _add_2_root_add_136_4_U101  ( .A1(_add_2_root_add_136_4_n46 ), .A2(_add_2_root_add_136_4_n47 ), .ZN(_add_2_root_add_136_4_n45 ) );
NOR2_X2 _add_2_root_add_136_4_U100  ( .A1(_add_2_root_add_136_4_n75 ), .A2(_add_2_root_add_136_4_n76 ), .ZN(_add_2_root_add_136_4_n80 ) );
NAND2_X2 _add_2_root_add_136_4_U99  ( .A1(_add_2_root_add_136_4_n324 ), .A2(_add_2_root_add_136_4_n265 ), .ZN(_add_2_root_add_136_4_n118 ) );
NOR2_X2 _add_2_root_add_136_4_U98  ( .A1(_add_2_root_add_136_4_n398 ), .A2(_add_2_root_add_136_4_n385 ), .ZN(_add_2_root_add_136_4_n397 ) );
XOR2_X2 _add_2_root_add_136_4_U97  ( .A(_add_2_root_add_136_4_n396 ), .B(_add_2_root_add_136_4_n397 ), .Z(N109) );
NOR2_X2 _add_2_root_add_136_4_U96  ( .A1(_add_2_root_add_136_4_n53 ), .A2(_add_2_root_add_136_4_n76 ), .ZN(_add_2_root_add_136_4_n79 ) );
NOR2_X2 _add_2_root_add_136_4_U95  ( .A1(_add_2_root_add_136_4_n79 ), .A2(_add_2_root_add_136_4_n75 ), .ZN(_add_2_root_add_136_4_n77 ) );
NOR2_X2 _add_2_root_add_136_4_U94  ( .A1(_add_2_root_add_136_4_n72 ), .A2(_add_2_root_add_136_4_n64 ), .ZN(_add_2_root_add_136_4_n78 ) );
NOR2_X2 _add_2_root_add_136_4_U93  ( .A1(_add_2_root_add_136_4_n421 ), .A2(_add_2_root_add_136_4_n35 ), .ZN(_add_2_root_add_136_4_n424 ) );
NOR2_X2 _add_2_root_add_136_4_U92  ( .A1(_add_2_root_add_136_4_n46 ), .A2(_add_2_root_add_136_4_n424 ), .ZN(_add_2_root_add_136_4_n423 ) );
NOR2_X2 _add_2_root_add_136_4_U91  ( .A1(_add_2_root_add_136_4_n406 ), .A2(_add_2_root_add_136_4_n419 ), .ZN(_add_2_root_add_136_4_n422 ) );
NOR2_X2 _add_2_root_add_136_4_U90  ( .A1(_add_2_root_add_136_4_n40 ), .A2(_add_2_root_add_136_4_n86 ), .ZN(_add_2_root_add_136_4_n154 ) );
NOR2_X2 _add_2_root_add_136_4_U89  ( .A1(_add_2_root_add_136_4_n64 ), .A2(_add_2_root_add_136_4_n74 ), .ZN(_add_2_root_add_136_4_n73 ) );
NOR2_X2 _add_2_root_add_136_4_U88  ( .A1(_add_2_root_add_136_4_n72 ), .A2(_add_2_root_add_136_4_n73 ), .ZN(_add_2_root_add_136_4_n70 ) );
NOR2_X2 _add_2_root_add_136_4_U87  ( .A1(_add_2_root_add_136_4_n6 ), .A2(_add_2_root_add_136_4_n65 ), .ZN(_add_2_root_add_136_4_n71 ) );
NOR2_X2 _add_2_root_add_136_4_U86  ( .A1(_add_2_root_add_136_4_n5 ), .A2(_add_2_root_add_136_4_n104 ), .ZN(_add_2_root_add_136_4_n113 ) );
AND3_X2 _add_2_root_add_136_4_U85  ( .A1(_add_2_root_add_136_4_n400 ), .A2(_add_2_root_add_136_4_n392 ), .A3(_add_2_root_add_136_4_n18 ), .ZN(_add_2_root_add_136_4_n24 ) );
NOR3_X2 _add_2_root_add_136_4_U84  ( .A1(_add_2_root_add_136_4_n230 ), .A2(_add_2_root_add_136_4_n231 ), .A3(_add_2_root_add_136_4_n232 ), .ZN(_add_2_root_add_136_4_n229 ) );
NAND3_X2 _add_2_root_add_136_4_U83  ( .A1(_add_2_root_add_136_4_n227 ), .A2(_add_2_root_add_136_4_n228 ), .A3(_add_2_root_add_136_4_n229 ), .ZN(_add_2_root_add_136_4_n226 ) );
NOR3_X2 _add_2_root_add_136_4_U82  ( .A1(_add_2_root_add_136_4_n270 ), .A2(_add_2_root_add_136_4_n271 ), .A3(_add_2_root_add_136_4_n272 ), .ZN(_add_2_root_add_136_4_n269 ) );
NAND3_X2 _add_2_root_add_136_4_U81  ( .A1(_add_2_root_add_136_4_n238 ), .A2(_add_2_root_add_136_4_n237 ), .A3(_add_2_root_add_136_4_n372 ), .ZN(_add_2_root_add_136_4_n278 ) );
NOR2_X2 _add_2_root_add_136_4_U80  ( .A1(_add_2_root_add_136_4_n54 ), .A2(_add_2_root_add_136_4_n1 ), .ZN(_add_2_root_add_136_4_n240 ) );
NOR2_X2 _add_2_root_add_136_4_U79  ( .A1(_add_2_root_add_136_4_n66 ), .A2(_add_2_root_add_136_4_n75 ), .ZN(_add_2_root_add_136_4_n74 ) );
NOR2_X2 _add_2_root_add_136_4_U78  ( .A1(_add_2_root_add_136_4_n153 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n295 ) );
NOR2_X2 _add_2_root_add_136_4_U77  ( .A1(_add_2_root_add_136_4_n295 ), .A2(_add_2_root_add_136_4_n296 ), .ZN(_add_2_root_add_136_4_n291 ) );
NOR2_X2 _add_2_root_add_136_4_U76  ( .A1(_add_2_root_add_136_4_n291 ), .A2(_add_2_root_add_136_4_n280 ), .ZN(_add_2_root_add_136_4_n284 ) );
NOR2_X2 _add_2_root_add_136_4_U75  ( .A1(_add_2_root_add_136_4_n105 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n266 ) );
NOR2_X2 _add_2_root_add_136_4_U74  ( .A1(_add_2_root_add_136_4_n114 ), .A2(_add_2_root_add_136_4_n115 ), .ZN(_add_2_root_add_136_4_n111 ) );
NOR2_X2 _add_2_root_add_136_4_U73  ( .A1(_add_2_root_add_136_4_n117 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n109 ) );
NOR2_X2 _add_2_root_add_136_4_U72  ( .A1(_add_2_root_add_136_4_n109 ), .A2(_add_2_root_add_136_4_n110 ), .ZN(_add_2_root_add_136_4_n96 ) );
NOR2_X2 _add_2_root_add_136_4_U71  ( .A1(_add_2_root_add_136_4_n53 ), .A2(_add_2_root_add_136_4_n54 ), .ZN(_add_2_root_add_136_4_n51 ) );
NOR2_X2 _add_2_root_add_136_4_U70  ( .A1(_add_2_root_add_136_4_n51 ), .A2(_add_2_root_add_136_4_n52 ), .ZN(_add_2_root_add_136_4_n50 ) );
NOR2_X2 _add_2_root_add_136_4_U69  ( .A1(_add_2_root_add_136_4_n273 ), .A2(_add_2_root_add_136_4_n274 ), .ZN(_add_2_root_add_136_4_n271 ) );
NOR2_X2 _add_2_root_add_136_4_U68  ( .A1(_add_2_root_add_136_4_n105 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n224 ) );
OR2_X4 _add_2_root_add_136_4_U67  ( .A1(_add_2_root_add_136_4_n225 ), .A2(_add_2_root_add_136_4_n226 ), .ZN(_add_2_root_add_136_4_n23 ) );
AND2_X2 _add_2_root_add_136_4_U66  ( .A1(_add_2_root_add_136_4_n23 ), .A2(_add_2_root_add_136_4_n224 ), .ZN(_add_2_root_add_136_4_n220 ) );
NOR2_X2 _add_2_root_add_136_4_U65  ( .A1(_add_2_root_add_136_4_n126 ), .A2(_add_2_root_add_136_4_n128 ), .ZN(_add_2_root_add_136_4_n277 ) );
INV_X4 _add_2_root_add_136_4_U64  ( .A(_add_2_root_add_136_4_n233 ), .ZN(_add_2_root_add_136_4_n185 ) );
NOR2_X2 _add_2_root_add_136_4_U63  ( .A1(_add_2_root_add_136_4_n248 ), .A2(_add_2_root_add_136_4_n249 ), .ZN(_add_2_root_add_136_4_n247 ) );
NOR3_X2 _add_2_root_add_136_4_U62  ( .A1(_add_2_root_add_136_4_n251 ), .A2(_add_2_root_add_136_4_n252 ), .A3(_add_2_root_add_136_4_n253 ), .ZN(_add_2_root_add_136_4_n245 ) );
NOR2_X2 _add_2_root_add_136_4_U61  ( .A1(_add_2_root_add_136_4_n128 ), .A2(_add_2_root_add_136_4_n247 ), .ZN(_add_2_root_add_136_4_n246 ) );
NOR2_X2 _add_2_root_add_136_4_U60  ( .A1(_add_2_root_add_136_4_n127 ), .A2(_add_2_root_add_136_4_n128 ), .ZN(_add_2_root_add_136_4_n320 ) );
NAND3_X2 _add_2_root_add_136_4_U59  ( .A1(_add_2_root_add_136_4_n184 ), .A2(_add_2_root_add_136_4_n125 ), .A3(_add_2_root_add_136_4_n320 ), .ZN(_add_2_root_add_136_4_n318 ) );
NOR2_X2 _add_2_root_add_136_4_U58  ( .A1(_add_2_root_add_136_4_n127 ), .A2(_add_2_root_add_136_4_n128 ), .ZN(_add_2_root_add_136_4_n183 ) );
NAND3_X2 _add_2_root_add_136_4_U57  ( .A1(_add_2_root_add_136_4_n184 ), .A2(_add_2_root_add_136_4_n125 ), .A3(_add_2_root_add_136_4_n183 ), .ZN(_add_2_root_add_136_4_n181 ) );
NOR2_X2 _add_2_root_add_136_4_U56  ( .A1(_add_2_root_add_136_4_n127 ), .A2(_add_2_root_add_136_4_n128 ), .ZN(_add_2_root_add_136_4_n124 ) );
NOR3_X2 _add_2_root_add_136_4_U55  ( .A1(_add_2_root_add_136_4_n126 ), .A2(_add_2_root_add_136_4_n127 ), .A3(_add_2_root_add_136_4_n128 ), .ZN(_add_2_root_add_136_4_n348 ) );
NAND3_X2 _add_2_root_add_136_4_U54  ( .A1(_add_2_root_add_136_4_n348 ), .A2(_add_2_root_add_136_4_n349 ), .A3(_add_2_root_add_136_4_n125 ), .ZN(_add_2_root_add_136_4_n306 ) );
NOR3_X2 _add_2_root_add_136_4_U53  ( .A1(_add_2_root_add_136_4_n257 ), .A2(_add_2_root_add_136_4_n258 ), .A3(_add_2_root_add_136_4_n259 ), .ZN(_add_2_root_add_136_4_n256 ) );
NOR2_X2 _add_2_root_add_136_4_U52  ( .A1(_add_2_root_add_136_4_n351 ), .A2(_add_2_root_add_136_4_n54 ), .ZN(_add_2_root_add_136_4_n350 ) );
AND2_X2 _add_2_root_add_136_4_U51  ( .A1(Kt[11]), .A2(SHA1_result[11]), .ZN(_add_2_root_add_136_4_n22 ) );
NOR2_X1 _add_2_root_add_136_4_U50  ( .A1(SHA1_result[11]), .A2(Kt[11]), .ZN(_add_2_root_add_136_4_n402 ) );
OR2_X4 _add_2_root_add_136_4_U49  ( .A1(_add_2_root_add_136_4_n64 ), .A2(_add_2_root_add_136_4_n65 ), .ZN(_add_2_root_add_136_4_n21 ) );
NOR2_X2 _add_2_root_add_136_4_U48  ( .A1(_add_2_root_add_136_4_n66 ), .A2(_add_2_root_add_136_4_n67 ), .ZN(_add_2_root_add_136_4_n20 ) );
NOR2_X2 _add_2_root_add_136_4_U47  ( .A1(_add_2_root_add_136_4_n20 ), .A2(_add_2_root_add_136_4_n21 ), .ZN(_add_2_root_add_136_4_n63 ) );
NAND3_X1 _add_2_root_add_136_4_U46  ( .A1(_add_2_root_add_136_4_n342 ), .A2(_add_2_root_add_136_4_n43 ), .A3(_add_2_root_add_136_4_n306 ), .ZN(_add_2_root_add_136_4_n341 ) );
NOR2_X1 _add_2_root_add_136_4_U45  ( .A1(_add_2_root_add_136_4_n241 ), .A2(_add_2_root_add_136_4_n233 ), .ZN(_add_2_root_add_136_4_n239 ) );
OR2_X2 _add_2_root_add_136_4_U44  ( .A1(_add_2_root_add_136_4_n284 ), .A2(_add_2_root_add_136_4_n285 ), .ZN(_add_2_root_add_136_4_n25 ) );
NOR3_X1 _add_2_root_add_136_4_U43  ( .A1(_add_2_root_add_136_4_n233 ), .A2(_add_2_root_add_136_4_n1 ), .A3(_add_2_root_add_136_4_n234 ), .ZN(_add_2_root_add_136_4_n232 ) );
NOR3_X1 _add_2_root_add_136_4_U42  ( .A1(_add_2_root_add_136_4_n233 ), .A2(_add_2_root_add_136_4_n1 ), .A3(_add_2_root_add_136_4_n62 ), .ZN(_add_2_root_add_136_4_n231 ) );
NAND3_X2 _add_2_root_add_136_4_U41  ( .A1(_add_2_root_add_136_4_n339 ), .A2(_add_2_root_add_136_4_n340 ), .A3(_add_2_root_add_136_4_n341 ), .ZN(_add_2_root_add_136_4_n19 ) );
XNOR2_X2 _add_2_root_add_136_4_U40  ( .A(_add_2_root_add_136_4_n19 ), .B(_add_2_root_add_136_4_n338 ), .ZN(N114) );
NOR2_X1 _add_2_root_add_136_4_U39  ( .A1(_add_2_root_add_136_4_n241 ), .A2(_add_2_root_add_136_4_n233 ), .ZN(_add_2_root_add_136_4_n364 ) );
NOR2_X1 _add_2_root_add_136_4_U38  ( .A1(_add_2_root_add_136_4_n233 ), .A2(_add_2_root_add_136_4_n244 ), .ZN(_add_2_root_add_136_4_n358 ) );
NOR3_X1 _add_2_root_add_136_4_U37  ( .A1(_add_2_root_add_136_4_n233 ), .A2(_add_2_root_add_136_4_n1 ), .A3(_add_2_root_add_136_4_n234 ), .ZN(_add_2_root_add_136_4_n126 ) );
NOR3_X1 _add_2_root_add_136_4_U36  ( .A1(_add_2_root_add_136_4_n235 ), .A2(_add_2_root_add_136_4_n233 ), .A3(_add_2_root_add_136_4_n236 ), .ZN(_add_2_root_add_136_4_n230 ) );
NAND2_X1 _add_2_root_add_136_4_U35  ( .A1(_add_2_root_add_136_4_n34 ), .A2(_add_2_root_add_136_4_n185 ), .ZN(_add_2_root_add_136_4_n274 ) );
NOR2_X1 _add_2_root_add_136_4_U34  ( .A1(_add_2_root_add_136_4_n233 ), .A2(_add_2_root_add_136_4_n236 ), .ZN(_add_2_root_add_136_4_n372 ) );
OR2_X1 _add_2_root_add_136_4_U33  ( .A1(SHA1_result[10]), .A2(Kt[10]), .ZN(_add_2_root_add_136_4_n41 ) );
NOR2_X1 _add_2_root_add_136_4_U32  ( .A1(SHA1_result[10]), .A2(Kt[10]), .ZN(_add_2_root_add_136_4_n409 ) );
NOR2_X1 _add_2_root_add_136_4_U31  ( .A1(SHA1_result[10]), .A2(Kt[10]), .ZN(_add_2_root_add_136_4_n419 ) );
NOR2_X1 _add_2_root_add_136_4_U30  ( .A1(SHA1_result[8]), .A2(Kt[8]), .ZN(_add_2_root_add_136_4_n49 ) );
NOR2_X1 _add_2_root_add_136_4_U29  ( .A1(_add_2_root_add_136_4_n395 ), .A2(_add_2_root_add_136_4_n233 ), .ZN(_add_2_root_add_136_4_n390 ) );
NAND2_X1 _add_2_root_add_136_4_U28  ( .A1(_add_2_root_add_136_4_n129 ), .A2(_add_2_root_add_136_4_n132 ), .ZN(_add_2_root_add_136_4_n270 ) );
NOR2_X1 _add_2_root_add_136_4_U27  ( .A1(_add_2_root_add_136_4_n233 ), .A2(_add_2_root_add_136_4_n244 ), .ZN(_add_2_root_add_136_4_n243 ) );
NOR2_X1 _add_2_root_add_136_4_U26  ( .A1(_add_2_root_add_136_4_n153 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n151 ) );
NOR2_X1 _add_2_root_add_136_4_U25  ( .A1(_add_2_root_add_136_4_n54 ), .A2(_add_2_root_add_136_4_n1 ), .ZN(_add_2_root_add_136_4_n365 ) );
NOR2_X1 _add_2_root_add_136_4_U24  ( .A1(_add_2_root_add_136_4_n54 ), .A2(_add_2_root_add_136_4_n1 ), .ZN(_add_2_root_add_136_4_n359 ) );
NOR2_X1 _add_2_root_add_136_4_U23  ( .A1(_add_2_root_add_136_4_n153 ), .A2(_add_2_root_add_136_4_n118 ), .ZN(_add_2_root_add_136_4_n323 ) );
INV_X2 _add_2_root_add_136_4_U22  ( .A(_add_2_root_add_136_4_n129 ), .ZN(_add_2_root_add_136_4_n251 ) );
NAND3_X1 _add_2_root_add_136_4_U21  ( .A1(_add_2_root_add_136_4_n304 ), .A2(_add_2_root_add_136_4_n305 ), .A3(_add_2_root_add_136_4_n306 ), .ZN(_add_2_root_add_136_4_n303 ) );
OR2_X4 _add_2_root_add_136_4_U20  ( .A1(_add_2_root_add_136_4_n53 ), .A2(_add_2_root_add_136_4_n401 ), .ZN(_add_2_root_add_136_4_n18 ) );
OR2_X4 _add_2_root_add_136_4_U19  ( .A1(SHA1_result[13]), .A2(Kt[13]), .ZN(_add_2_root_add_136_4_n17 ) );
OR3_X4 _add_2_root_add_136_4_U18  ( .A1(_add_2_root_add_136_4_n103 ), .A2(_add_2_root_add_136_4_n5 ), .A3(_add_2_root_add_136_4_n104 ), .ZN(_add_2_root_add_136_4_n16 ) );
AND2_X4 _add_2_root_add_136_4_U17  ( .A1(Kt[25]), .A2(SHA1_result[25]), .ZN(_add_2_root_add_136_4_n15 ) );
OR3_X4 _add_2_root_add_136_4_U16  ( .A1(_add_2_root_add_136_4_n384 ), .A2(_add_2_root_add_136_4_n368 ), .A3(_add_2_root_add_136_4_n385 ), .ZN(_add_2_root_add_136_4_n14 ) );
AND2_X4 _add_2_root_add_136_4_U15  ( .A1(_add_2_root_add_136_4_n198 ), .A2(_add_2_root_add_136_4_n207 ), .ZN(_add_2_root_add_136_4_n13 ) );
XOR2_X2 _add_2_root_add_136_4_U14  ( .A(_add_2_root_add_136_4_n186 ), .B(_add_2_root_add_136_4_n10 ), .Z(N124) );
AND3_X4 _add_2_root_add_136_4_U13  ( .A1(_add_2_root_add_136_4_n242 ), .A2(_add_2_root_add_136_4_n185 ), .A3(_add_2_root_add_136_4_n394 ), .ZN(_add_2_root_add_136_4_n11 ) );
AND2_X4 _add_2_root_add_136_4_U12  ( .A1(_add_2_root_add_136_4_n106 ), .A2(_add_2_root_add_136_4_n171 ), .ZN(_add_2_root_add_136_4_n10 ) );
OR3_X4 _add_2_root_add_136_4_U11  ( .A1(_add_2_root_add_136_4_n419 ), .A2(_add_2_root_add_136_4_n49 ), .A3(_add_2_root_add_136_4_n47 ), .ZN(_add_2_root_add_136_4_n9 ) );
AND2_X4 _add_2_root_add_136_4_U10  ( .A1(Kt[24]), .A2(SHA1_result[24]), .ZN(_add_2_root_add_136_4_n8 ) );
AND2_X4 _add_2_root_add_136_4_U9  ( .A1(Kt[20]), .A2(SHA1_result[20]), .ZN(_add_2_root_add_136_4_n7 ) );
AND2_X4 _add_2_root_add_136_4_U8  ( .A1(Kt[6]), .A2(SHA1_result[6]), .ZN(_add_2_root_add_136_4_n6 ) );
AND2_X4 _add_2_root_add_136_4_U7  ( .A1(_add_2_root_add_136_4_n166 ), .A2(_add_2_root_add_136_4_n150 ), .ZN(_add_2_root_add_136_4_n5 ) );
OR2_X4 _add_2_root_add_136_4_U6  ( .A1(SHA1_result[4]), .A2(Kt[4]), .ZN(_add_2_root_add_136_4_n4 ) );
OR2_X4 _add_2_root_add_136_4_U5  ( .A1(SHA1_result[9]), .A2(Kt[9]), .ZN(_add_2_root_add_136_4_n3 ) );
AND2_X4 _add_2_root_add_136_4_U4  ( .A1(Kt[8]), .A2(SHA1_result[8]), .ZN(_add_2_root_add_136_4_n2 ) );
NAND3_X2 _add_2_root_add_136_4_U3  ( .A1(_add_2_root_add_136_4_n17 ), .A2(_add_2_root_add_136_4_n42 ), .A3(_add_2_root_add_136_4_n376 ), .ZN(_add_2_root_add_136_4_n1 ) );
NOR3_X2 _add_2_root_add_136_4_U2  ( .A1(_add_2_root_add_136_4_n355 ), .A2(_add_2_root_add_136_4_n356 ), .A3(_add_2_root_add_136_4_n357 ), .ZN(_add_2_root_add_136_4_n349 ) );
NAND2_X2 _add_514_U409  ( .A1(H2[7]), .A2(next_C[7]), .ZN(_add_514_n50 ) );
NAND2_X2 _add_514_U408  ( .A1(H2[6]), .A2(next_C[6]), .ZN(_add_514_n53 ) );
NAND2_X2 _add_514_U407  ( .A1(_add_514_n50 ), .A2(_add_514_n53 ), .ZN(_add_514_n332 ) );
NAND2_X2 _add_514_U406  ( .A1(_add_514_n377 ), .A2(_add_514_n332 ), .ZN(_add_514_n375 ) );
NAND2_X2 _add_514_U405  ( .A1(H2[8]), .A2(next_C[8]), .ZN(_add_514_n44 ) );
NAND2_X2 _add_514_U404  ( .A1(H2[4]), .A2(next_C[4]), .ZN(_add_514_n280 ) );
NAND2_X2 _add_514_U403  ( .A1(H2[5]), .A2(next_C[5]), .ZN(_add_514_n58 ) );
NAND2_X2 _add_514_U402  ( .A1(_add_514_n280 ), .A2(_add_514_n58 ), .ZN(_add_514_n353 ) );
INV_X4 _add_514_U401  ( .A(next_C[0]), .ZN(_add_514_n373 ) );
INV_X4 _add_514_U400  ( .A(H2[0]), .ZN(_add_514_n374 ) );
INV_X4 _add_514_U399  ( .A(_add_514_n69 ), .ZN(_add_514_n371 ) );
INV_X4 _add_514_U398  ( .A(_add_514_n117 ), .ZN(_add_514_n372 ) );
NAND2_X2 _add_514_U397  ( .A1(H2[1]), .A2(next_C[1]), .ZN(_add_514_n369 ) );
XNOR2_X2 _add_514_U396  ( .A(_add_514_n360 ), .B(_add_514_n361 ), .ZN(N926));
XNOR2_X2 _add_514_U395  ( .A(_add_514_n354 ), .B(_add_514_n355 ), .ZN(N927));
INV_X4 _add_514_U394  ( .A(_add_514_n332 ), .ZN(_add_514_n351 ) );
NAND2_X2 _add_514_U393  ( .A1(_add_514_n333 ), .A2(_add_514_n353 ), .ZN(_add_514_n352 ) );
NAND2_X2 _add_514_U392  ( .A1(_add_514_n351 ), .A2(_add_514_n352 ), .ZN(_add_514_n350 ) );
INV_X4 _add_514_U391  ( .A(_add_514_n285 ), .ZN(_add_514_n345 ) );
INV_X4 _add_514_U390  ( .A(_add_514_n284 ), .ZN(_add_514_n346 ) );
NAND2_X2 _add_514_U389  ( .A1(H2[8]), .A2(next_C[8]), .ZN(_add_514_n342 ) );
NAND2_X2 _add_514_U388  ( .A1(next_C[9]), .A2(H2[9]), .ZN(_add_514_n341 ) );
INV_X4 _add_514_U387  ( .A(_add_514_n138 ), .ZN(_add_514_n209 ) );
NAND2_X2 _add_514_U386  ( .A1(H2[12]), .A2(next_C[12]), .ZN(_add_514_n299 ));
INV_X4 _add_514_U385  ( .A(_add_514_n299 ), .ZN(_add_514_n312 ) );
INV_X4 _add_514_U384  ( .A(_add_514_n325 ), .ZN(_add_514_n270 ) );
XNOR2_X2 _add_514_U383  ( .A(_add_514_n335 ), .B(_add_514_n336 ), .ZN(N928));
NAND2_X2 _add_514_U382  ( .A1(_add_514_n280 ), .A2(_add_514_n58 ), .ZN(_add_514_n334 ) );
NAND2_X2 _add_514_U381  ( .A1(_add_514_n332 ), .A2(_add_514_n2 ), .ZN(_add_514_n331 ) );
NAND2_X2 _add_514_U380  ( .A1(_add_514_n345 ), .A2(_add_514_n325 ), .ZN(_add_514_n324 ) );
NAND2_X2 _add_514_U379  ( .A1(H2[13]), .A2(next_C[13]), .ZN(_add_514_n309 ));
INV_X4 _add_514_U378  ( .A(_add_514_n309 ), .ZN(_add_514_n318 ) );
XNOR2_X2 _add_514_U377  ( .A(_add_514_n320 ), .B(_add_514_n321 ), .ZN(N929));
INV_X4 _add_514_U376  ( .A(_add_514_n310 ), .ZN(_add_514_n316 ) );
XNOR2_X2 _add_514_U375  ( .A(_add_514_n314 ), .B(_add_514_n315 ), .ZN(N930));
NAND2_X2 _add_514_U374  ( .A1(H2[15]), .A2(next_C[15]), .ZN(_add_514_n296 ));
NAND2_X2 _add_514_U373  ( .A1(_add_514_n296 ), .A2(_add_514_n271 ), .ZN(_add_514_n306 ) );
NAND2_X2 _add_514_U372  ( .A1(H2[16]), .A2(next_C[16]), .ZN(_add_514_n264 ));
NAND2_X2 _add_514_U371  ( .A1(_add_514_n264 ), .A2(_add_514_n266 ), .ZN(_add_514_n267 ) );
INV_X4 _add_514_U370  ( .A(_add_514_n271 ), .ZN(_add_514_n275 ) );
INV_X4 _add_514_U369  ( .A(_add_514_n272 ), .ZN(_add_514_n301 ) );
INV_X4 _add_514_U368  ( .A(_add_514_n269 ), .ZN(_add_514_n302 ) );
NAND2_X2 _add_514_U367  ( .A1(_add_514_n292 ), .A2(_add_514_n293 ), .ZN(_add_514_n147 ) );
NAND2_X2 _add_514_U366  ( .A1(H2[2]), .A2(next_C[2]), .ZN(_add_514_n289 ) );
NAND2_X2 _add_514_U365  ( .A1(H2[0]), .A2(next_C[0]), .ZN(_add_514_n149 ) );
NAND2_X2 _add_514_U364  ( .A1(H2[1]), .A2(next_C[1]), .ZN(_add_514_n148 ) );
NAND2_X2 _add_514_U363  ( .A1(_add_514_n56 ), .A2(_add_514_n50 ), .ZN(_add_514_n282 ) );
NAND2_X2 _add_514_U362  ( .A1(_add_514_n281 ), .A2(_add_514_n282 ), .ZN(_add_514_n276 ) );
NAND2_X2 _add_514_U361  ( .A1(_add_514_n58 ), .A2(_add_514_n53 ), .ZN(_add_514_n278 ) );
INV_X4 _add_514_U360  ( .A(_add_514_n50 ), .ZN(_add_514_n279 ) );
INV_X4 _add_514_U359  ( .A(_add_514_n280 ), .ZN(_add_514_n64 ) );
NAND2_X2 _add_514_U358  ( .A1(_add_514_n273 ), .A2(_add_514_n274 ), .ZN(_add_514_n150 ) );
INV_X4 _add_514_U357  ( .A(_add_514_n150 ), .ZN(_add_514_n207 ) );
XNOR2_X2 _add_514_U356  ( .A(_add_514_n267 ), .B(_add_514_n247 ), .ZN(N932));
INV_X4 _add_514_U355  ( .A(_add_514_n248 ), .ZN(_add_514_n266 ) );
NAND2_X2 _add_514_U354  ( .A1(_add_514_n247 ), .A2(_add_514_n266 ), .ZN(_add_514_n265 ) );
NAND2_X2 _add_514_U353  ( .A1(_add_514_n264 ), .A2(_add_514_n265 ), .ZN(_add_514_n261 ) );
INV_X4 _add_514_U352  ( .A(_add_514_n259 ), .ZN(_add_514_n250 ) );
NAND2_X2 _add_514_U351  ( .A1(H2[17]), .A2(next_C[17]), .ZN(_add_514_n258 ));
INV_X4 _add_514_U350  ( .A(_add_514_n258 ), .ZN(_add_514_n263 ) );
INV_X4 _add_514_U349  ( .A(_add_514_n247 ), .ZN(_add_514_n260 ) );
NAND2_X2 _add_514_U348  ( .A1(_add_514_n257 ), .A2(_add_514_n258 ), .ZN(_add_514_n254 ) );
NAND2_X2 _add_514_U347  ( .A1(H2[18]), .A2(next_C[18]), .ZN(_add_514_n253 ));
NAND2_X2 _add_514_U346  ( .A1(_add_514_n253 ), .A2(_add_514_n251 ), .ZN(_add_514_n255 ) );
NAND2_X2 _add_514_U345  ( .A1(_add_514_n254 ), .A2(_add_514_n251 ), .ZN(_add_514_n252 ) );
NAND2_X2 _add_514_U344  ( .A1(_add_514_n252 ), .A2(_add_514_n253 ), .ZN(_add_514_n211 ) );
INV_X4 _add_514_U343  ( .A(_add_514_n211 ), .ZN(_add_514_n245 ) );
INV_X4 _add_514_U342  ( .A(_add_514_n251 ), .ZN(_add_514_n249 ) );
NAND2_X2 _add_514_U341  ( .A1(_add_514_n235 ), .A2(_add_514_n247 ), .ZN(_add_514_n246 ) );
NAND2_X2 _add_514_U340  ( .A1(_add_514_n245 ), .A2(_add_514_n246 ), .ZN(_add_514_n243 ) );
NAND2_X2 _add_514_U339  ( .A1(H2[19]), .A2(next_C[19]), .ZN(_add_514_n129 ));
NAND2_X2 _add_514_U338  ( .A1(_add_514_n212 ), .A2(_add_514_n129 ), .ZN(_add_514_n244 ) );
XNOR2_X2 _add_514_U337  ( .A(_add_514_n243 ), .B(_add_514_n244 ), .ZN(N935));
NAND2_X2 _add_514_U336  ( .A1(H2[1]), .A2(next_C[1]), .ZN(_add_514_n116 ) );
INV_X4 _add_514_U335  ( .A(_add_514_n116 ), .ZN(_add_514_n241 ) );
XNOR2_X2 _add_514_U334  ( .A(_add_514_n242 ), .B(_add_514_n240 ), .ZN(N917));
INV_X4 _add_514_U333  ( .A(_add_514_n210 ), .ZN(_add_514_n137 ) );
NAND2_X2 _add_514_U332  ( .A1(_add_514_n137 ), .A2(_add_514_n138 ), .ZN(_add_514_n237 ) );
INV_X4 _add_514_U331  ( .A(_add_514_n136 ), .ZN(_add_514_n238 ) );
INV_X4 _add_514_U330  ( .A(_add_514_n151 ), .ZN(_add_514_n239 ) );
NAND4_X2 _add_514_U329  ( .A1(_add_514_n206 ), .A2(_add_514_n237 ), .A3(_add_514_n238 ), .A4(_add_514_n239 ), .ZN(_add_514_n236 ) );
NAND2_X2 _add_514_U328  ( .A1(_add_514_n235 ), .A2(_add_514_n212 ), .ZN(_add_514_n131 ) );
NAND2_X2 _add_514_U327  ( .A1(_add_514_n211 ), .A2(_add_514_n212 ), .ZN(_add_514_n152 ) );
NAND2_X2 _add_514_U326  ( .A1(_add_514_n152 ), .A2(_add_514_n129 ), .ZN(_add_514_n233 ) );
XNOR2_X2 _add_514_U325  ( .A(_add_514_n221 ), .B(_add_514_n231 ), .ZN(N936));
NAND2_X2 _add_514_U324  ( .A1(H2[21]), .A2(next_C[21]), .ZN(_add_514_n220 ));
NAND2_X2 _add_514_U323  ( .A1(_add_514_n220 ), .A2(_add_514_n222 ), .ZN(_add_514_n229 ) );
INV_X4 _add_514_U322  ( .A(_add_514_n222 ), .ZN(_add_514_n228 ) );
NAND2_X2 _add_514_U321  ( .A1(_add_514_n219 ), .A2(_add_514_n220 ), .ZN(_add_514_n227 ) );
NAND2_X2 _add_514_U320  ( .A1(H2[22]), .A2(next_C[22]), .ZN(_add_514_n197 ));
NAND2_X2 _add_514_U319  ( .A1(_add_514_n218 ), .A2(_add_514_n197 ), .ZN(_add_514_n225 ) );
INV_X4 _add_514_U318  ( .A(_add_514_n224 ), .ZN(_add_514_n223 ) );
NAND2_X2 _add_514_U317  ( .A1(_add_514_n219 ), .A2(_add_514_n220 ), .ZN(_add_514_n217 ) );
NAND2_X2 _add_514_U316  ( .A1(_add_514_n217 ), .A2(_add_514_n218 ), .ZN(_add_514_n196 ) );
NAND2_X2 _add_514_U315  ( .A1(_add_514_n196 ), .A2(_add_514_n197 ), .ZN(_add_514_n216 ) );
NAND2_X2 _add_514_U314  ( .A1(H2[23]), .A2(next_C[23]), .ZN(_add_514_n128 ));
NAND2_X2 _add_514_U313  ( .A1(_add_514_n125 ), .A2(_add_514_n128 ), .ZN(_add_514_n214 ) );
INV_X4 _add_514_U312  ( .A(_add_514_n213 ), .ZN(_add_514_n201 ) );
NAND2_X2 _add_514_U311  ( .A1(_add_514_n201 ), .A2(_add_514_n125 ), .ZN(_add_514_n99 ) );
INV_X4 _add_514_U310  ( .A(_add_514_n99 ), .ZN(_add_514_n203 ) );
NAND3_X2 _add_514_U309  ( .A1(_add_514_n211 ), .A2(_add_514_n212 ), .A3(_add_514_n203 ), .ZN(_add_514_n190 ) );
INV_X4 _add_514_U308  ( .A(_add_514_n131 ), .ZN(_add_514_n204 ) );
INV_X4 _add_514_U307  ( .A(_add_514_n129 ), .ZN(_add_514_n200 ) );
NAND2_X2 _add_514_U306  ( .A1(_add_514_n200 ), .A2(_add_514_n201 ), .ZN(_add_514_n199 ) );
NAND2_X2 _add_514_U305  ( .A1(_add_514_n199 ), .A2(_add_514_n128 ), .ZN(_add_514_n198 ) );
NAND2_X2 _add_514_U304  ( .A1(_add_514_n198 ), .A2(_add_514_n125 ), .ZN(_add_514_n186 ) );
NAND2_X2 _add_514_U303  ( .A1(_add_514_n196 ), .A2(_add_514_n197 ), .ZN(_add_514_n126 ) );
NAND2_X2 _add_514_U302  ( .A1(_add_514_n126 ), .A2(_add_514_n125 ), .ZN(_add_514_n187 ) );
NAND2_X2 _add_514_U301  ( .A1(H2[24]), .A2(next_C[24]), .ZN(_add_514_n193 ));
INV_X4 _add_514_U300  ( .A(_add_514_n193 ), .ZN(_add_514_n195 ) );
XNOR2_X2 _add_514_U299  ( .A(_add_514_n166 ), .B(_add_514_n194 ), .ZN(N940));
NAND2_X2 _add_514_U298  ( .A1(_add_514_n10 ), .A2(_add_514_n193 ), .ZN(_add_514_n191 ) );
NAND2_X2 _add_514_U297  ( .A1(H2[25]), .A2(next_C[25]), .ZN(_add_514_n174 ));
NAND2_X2 _add_514_U296  ( .A1(_add_514_n174 ), .A2(_add_514_n175 ), .ZN(_add_514_n192 ) );
XNOR2_X2 _add_514_U295  ( .A(_add_514_n191 ), .B(_add_514_n192 ), .ZN(N941));
INV_X4 _add_514_U294  ( .A(_add_514_n190 ), .ZN(_add_514_n183 ) );
INV_X4 _add_514_U293  ( .A(_add_514_n189 ), .ZN(_add_514_n188 ) );
NAND2_X2 _add_514_U292  ( .A1(_add_514_n186 ), .A2(_add_514_n187 ), .ZN(_add_514_n185 ) );
NAND2_X2 _add_514_U291  ( .A1(_add_514_n175 ), .A2(_add_514_n176 ), .ZN(_add_514_n182 ) );
NAND2_X2 _add_514_U290  ( .A1(_add_514_n173 ), .A2(_add_514_n174 ), .ZN(_add_514_n180 ) );
NAND2_X2 _add_514_U289  ( .A1(H2[26]), .A2(next_C[26]), .ZN(_add_514_n163 ));
NAND2_X2 _add_514_U288  ( .A1(_add_514_n172 ), .A2(_add_514_n163 ), .ZN(_add_514_n178 ) );
INV_X4 _add_514_U287  ( .A(_add_514_n177 ), .ZN(_add_514_n176 ) );
NAND2_X2 _add_514_U286  ( .A1(_add_514_n173 ), .A2(_add_514_n174 ), .ZN(_add_514_n171 ) );
NAND2_X2 _add_514_U285  ( .A1(_add_514_n171 ), .A2(_add_514_n172 ), .ZN(_add_514_n164 ) );
NAND2_X2 _add_514_U284  ( .A1(_add_514_n164 ), .A2(_add_514_n163 ), .ZN(_add_514_n170 ) );
NAND2_X2 _add_514_U283  ( .A1(H2[27]), .A2(next_C[27]), .ZN(_add_514_n162 ));
NAND2_X2 _add_514_U282  ( .A1(_add_514_n154 ), .A2(_add_514_n162 ), .ZN(_add_514_n168 ) );
INV_X4 _add_514_U281  ( .A(_add_514_n167 ), .ZN(_add_514_n155 ) );
INV_X4 _add_514_U280  ( .A(_add_514_n166 ), .ZN(_add_514_n165 ) );
NAND2_X2 _add_514_U279  ( .A1(_add_514_n7 ), .A2(_add_514_n154 ), .ZN(_add_514_n161 ) );
NAND2_X2 _add_514_U278  ( .A1(_add_514_n160 ), .A2(_add_514_n161 ), .ZN(_add_514_n156 ) );
INV_X4 _add_514_U277  ( .A(H2[28]), .ZN(_add_514_n158 ) );
INV_X4 _add_514_U276  ( .A(next_C[28]), .ZN(_add_514_n159 ) );
NAND2_X2 _add_514_U275  ( .A1(_add_514_n158 ), .A2(_add_514_n159 ), .ZN(_add_514_n153 ) );
NAND2_X2 _add_514_U274  ( .A1(H2[28]), .A2(next_C[28]), .ZN(_add_514_n114 ));
NAND2_X2 _add_514_U273  ( .A1(_add_514_n153 ), .A2(_add_514_n114 ), .ZN(_add_514_n157 ) );
XNOR2_X2 _add_514_U272  ( .A(_add_514_n156 ), .B(_add_514_n157 ), .ZN(N944));
INV_X4 _add_514_U271  ( .A(_add_514_n114 ), .ZN(_add_514_n94 ) );
INV_X4 _add_514_U270  ( .A(_add_514_n110 ), .ZN(_add_514_n85 ) );
NAND4_X2 _add_514_U269  ( .A1(_add_514_n148 ), .A2(_add_514_n71 ), .A3(_add_514_n149 ), .A4(_add_514_n143 ), .ZN(_add_514_n144 ) );
NAND2_X2 _add_514_U268  ( .A1(_add_514_n144 ), .A2(_add_514_n145 ), .ZN(_add_514_n139 ) );
NAND2_X2 _add_514_U267  ( .A1(_add_514_n71 ), .A2(_add_514_n143 ), .ZN(_add_514_n142 ) );
NAND2_X2 _add_514_U266  ( .A1(_add_514_n137 ), .A2(_add_514_n138 ), .ZN(_add_514_n135 ) );
NAND2_X2 _add_514_U265  ( .A1(_add_514_n135 ), .A2(_add_514_n238 ), .ZN(_add_514_n134 ) );
INV_X4 _add_514_U264  ( .A(_add_514_n128 ), .ZN(_add_514_n127 ) );
NAND2_X2 _add_514_U263  ( .A1(_add_514_n127 ), .A2(_add_514_n4 ), .ZN(_add_514_n113 ) );
INV_X4 _add_514_U262  ( .A(_add_514_n113 ), .ZN(_add_514_n87 ) );
NAND2_X2 _add_514_U261  ( .A1(H2[29]), .A2(next_C[29]), .ZN(_add_514_n96 ));
INV_X4 _add_514_U260  ( .A(H2[29]), .ZN(_add_514_n120 ) );
INV_X4 _add_514_U259  ( .A(next_C[29]), .ZN(_add_514_n121 ) );
NAND2_X2 _add_514_U258  ( .A1(_add_514_n120 ), .A2(_add_514_n121 ), .ZN(_add_514_n109 ) );
NAND2_X2 _add_514_U257  ( .A1(_add_514_n96 ), .A2(_add_514_n109 ), .ZN(_add_514_n119 ) );
XNOR2_X2 _add_514_U256  ( .A(_add_514_n118 ), .B(_add_514_n119 ), .ZN(N945));
NAND2_X2 _add_514_U255  ( .A1(H2[2]), .A2(next_C[2]), .ZN(_add_514_n74 ) );
NAND2_X2 _add_514_U254  ( .A1(_add_514_n1 ), .A2(_add_514_n74 ), .ZN(_add_514_n115 ) );
NAND2_X2 _add_514_U253  ( .A1(_add_514_n25 ), .A2(_add_514_n116 ), .ZN(_add_514_n77 ) );
XNOR2_X2 _add_514_U252  ( .A(_add_514_n115 ), .B(_add_514_n77 ), .ZN(N918));
INV_X4 _add_514_U251  ( .A(_add_514_n109 ), .ZN(_add_514_n101 ) );
NAND2_X2 _add_514_U250  ( .A1(_add_514_n27 ), .A2(_add_514_n109 ), .ZN(_add_514_n105 ) );
INV_X4 _add_514_U249  ( .A(_add_514_n97 ), .ZN(_add_514_n108 ) );
NAND4_X2 _add_514_U248  ( .A1(_add_514_n203 ), .A2(_add_514_n108 ), .A3(_add_514_n109 ), .A4(_add_514_n4 ), .ZN(_add_514_n107 ) );
NAND4_X2 _add_514_U247  ( .A1(_add_514_n104 ), .A2(_add_514_n105 ), .A3(_add_514_n106 ), .A4(_add_514_n107 ), .ZN(_add_514_n102 ) );
NAND2_X2 _add_514_U246  ( .A1(H2[30]), .A2(next_C[30]), .ZN(_add_514_n95 ));
NAND2_X2 _add_514_U245  ( .A1(_add_514_n95 ), .A2(_add_514_n91 ), .ZN(_add_514_n103 ) );
XNOR2_X2 _add_514_U244  ( .A(_add_514_n102 ), .B(_add_514_n103 ), .ZN(N946));
INV_X4 _add_514_U243  ( .A(_add_514_n91 ), .ZN(_add_514_n100 ) );
NAND2_X2 _add_514_U242  ( .A1(_add_514_n86 ), .A2(_add_514_n4 ), .ZN(_add_514_n98 ) );
NAND2_X2 _add_514_U241  ( .A1(_add_514_n94 ), .A2(_add_514_n86 ), .ZN(_add_514_n93 ) );
NAND2_X2 _add_514_U240  ( .A1(_add_514_n92 ), .A2(_add_514_n93 ), .ZN(_add_514_n90 ) );
NAND2_X2 _add_514_U239  ( .A1(_add_514_n90 ), .A2(_add_514_n91 ), .ZN(_add_514_n88 ) );
NAND2_X2 _add_514_U238  ( .A1(_add_514_n27 ), .A2(_add_514_n86 ), .ZN(_add_514_n89 ) );
NAND2_X2 _add_514_U237  ( .A1(_add_514_n88 ), .A2(_add_514_n89 ), .ZN(_add_514_n81 ) );
NAND2_X2 _add_514_U236  ( .A1(_add_514_n87 ), .A2(_add_514_n86 ), .ZN(_add_514_n83 ) );
NAND2_X2 _add_514_U235  ( .A1(_add_514_n85 ), .A2(_add_514_n86 ), .ZN(_add_514_n84 ) );
NAND2_X2 _add_514_U234  ( .A1(_add_514_n83 ), .A2(_add_514_n84 ), .ZN(_add_514_n82 ) );
NOR2_X2 _add_514_U233  ( .A1(_add_514_n81 ), .A2(_add_514_n82 ), .ZN(_add_514_n80 ) );
NAND2_X2 _add_514_U232  ( .A1(_add_514_n15 ), .A2(_add_514_n80 ), .ZN(_add_514_n78 ) );
XNOR2_X2 _add_514_U231  ( .A(_add_514_n78 ), .B(_add_514_n79 ), .ZN(N947) );
INV_X4 _add_514_U230  ( .A(_add_514_n77 ), .ZN(_add_514_n76 ) );
INV_X4 _add_514_U229  ( .A(_add_514_n74 ), .ZN(_add_514_n73 ) );
INV_X4 _add_514_U228  ( .A(_add_514_n71 ), .ZN(_add_514_n70 ) );
XNOR2_X2 _add_514_U227  ( .A(_add_514_n67 ), .B(_add_514_n68 ), .ZN(N919) );
XNOR2_X2 _add_514_U226  ( .A(_add_514_n46 ), .B(_add_514_n66 ), .ZN(N920) );
INV_X4 _add_514_U225  ( .A(_add_514_n58 ), .ZN(_add_514_n62 ) );
XNOR2_X2 _add_514_U224  ( .A(_add_514_n60 ), .B(_add_514_n61 ), .ZN(N921) );
NAND2_X2 _add_514_U223  ( .A1(_add_514_n53 ), .A2(_add_514_n55 ), .ZN(_add_514_n57 ) );
NAND2_X2 _add_514_U222  ( .A1(_add_514_n16 ), .A2(_add_514_n58 ), .ZN(_add_514_n54 ) );
XNOR2_X2 _add_514_U221  ( .A(_add_514_n57 ), .B(_add_514_n54 ), .ZN(N922) );
INV_X4 _add_514_U220  ( .A(_add_514_n56 ), .ZN(_add_514_n55 ) );
NAND2_X2 _add_514_U219  ( .A1(_add_514_n54 ), .A2(_add_514_n55 ), .ZN(_add_514_n52 ) );
NAND2_X2 _add_514_U218  ( .A1(_add_514_n52 ), .A2(_add_514_n53 ), .ZN(_add_514_n48 ) );
NAND2_X2 _add_514_U217  ( .A1(_add_514_n50 ), .A2(_add_514_n2 ), .ZN(_add_514_n49 ) );
XNOR2_X2 _add_514_U216  ( .A(_add_514_n48 ), .B(_add_514_n49 ), .ZN(N923) );
INV_X4 _add_514_U215  ( .A(_add_514_n44 ), .ZN(_add_514_n43 ) );
XNOR2_X2 _add_514_U214  ( .A(_add_514_n40 ), .B(_add_514_n41 ), .ZN(N924) );
XNOR2_X2 _add_514_U213  ( .A(_add_514_n37 ), .B(_add_514_n38 ), .ZN(N925) );
NAND2_X1 _add_514_U212  ( .A1(H2[3]), .A2(n13081), .ZN(_add_514_n71 ) );
NOR2_X1 _add_514_U211  ( .A1(n13081), .A2(H2[3]), .ZN(_add_514_n69 ) );
NAND2_X2 _add_514_U210  ( .A1(_add_514_n71 ), .A2(_add_514_n143 ), .ZN(_add_514_n368 ) );
NAND2_X2 _add_514_U209  ( .A1(_add_514_n150 ), .A2(_add_514_n239 ), .ZN(_add_514_n132 ) );
NAND3_X1 _add_514_U208  ( .A1(next_C[2]), .A2(_add_514_n371 ), .A3(H2[2]),.ZN(_add_514_n143 ) );
NAND3_X1 _add_514_U207  ( .A1(H2[2]), .A2(_add_514_n371 ), .A3(next_C[2]),.ZN(_add_514_n290 ) );
OR2_X2 _add_514_U206  ( .A1(H2[27]), .A2(next_C[27]), .ZN(_add_514_n154 ) );
OR2_X2 _add_514_U205  ( .A1(H2[25]), .A2(next_C[25]), .ZN(_add_514_n175 ) );
AND2_X2 _add_514_U204  ( .A1(H2[11]), .A2(next_C[11]), .ZN(_add_514_n35 ) );
NOR2_X1 _add_514_U203  ( .A1(next_C[10]), .A2(H2[10]), .ZN(_add_514_n343 ));
AND2_X2 _add_514_U202  ( .A1(H2[9]), .A2(next_C[9]), .ZN(_add_514_n34 ) );
NOR2_X1 _add_514_U201  ( .A1(next_C[5]), .A2(H2[5]), .ZN(_add_514_n365 ) );
NOR2_X1 _add_514_U200  ( .A1(next_C[6]), .A2(H2[6]), .ZN(_add_514_n366 ) );
AND2_X2 _add_514_U199  ( .A1(H2[20]), .A2(next_C[20]), .ZN(_add_514_n33 ) );
NAND3_X1 _add_514_U198  ( .A1(H2[13]), .A2(next_C[13]), .A3(_add_514_n271 ),.ZN(_add_514_n298 ) );
NAND3_X1 _add_514_U197  ( .A1(next_C[20]), .A2(H2[20]), .A3(_add_514_n222 ),.ZN(_add_514_n219 ) );
NAND3_X1 _add_514_U196  ( .A1(next_C[24]), .A2(H2[24]), .A3(_add_514_n175 ),.ZN(_add_514_n173 ) );
NOR2_X1 _add_514_U195  ( .A1(next_C[10]), .A2(H2[10]), .ZN(_add_514_n340 ));
NOR2_X1 _add_514_U194  ( .A1(next_C[10]), .A2(H2[10]), .ZN(_add_514_n348 ));
NAND3_X1 _add_514_U193  ( .A1(next_C[16]), .A2(H2[16]), .A3(_add_514_n259 ),.ZN(_add_514_n257 ) );
NOR2_X1 _add_514_U192  ( .A1(next_C[4]), .A2(H2[4]), .ZN(_add_514_n65 ) );
NOR2_X1 _add_514_U191  ( .A1(next_C[8]), .A2(H2[8]), .ZN(_add_514_n327 ) );
NOR2_X1 _add_514_U190  ( .A1(next_C[10]), .A2(H2[10]), .ZN(_add_514_n357 ));
NOR2_X1 _add_514_U189  ( .A1(next_C[10]), .A2(H2[10]), .ZN(_add_514_n283 ));
NOR2_X1 _add_514_U188  ( .A1(next_C[11]), .A2(H2[11]), .ZN(_add_514_n285 ));
NOR2_X1 _add_514_U187  ( .A1(next_C[11]), .A2(H2[11]), .ZN(_add_514_n305 ));
NOR2_X1 _add_514_U186  ( .A1(next_C[9]), .A2(H2[9]), .ZN(_add_514_n284 ) );
NOR2_X1 _add_514_U185  ( .A1(next_C[6]), .A2(H2[6]), .ZN(_add_514_n56 ) );
NOR2_X1 _add_514_U184  ( .A1(next_C[9]), .A2(H2[9]), .ZN(_add_514_n39 ) );
OR2_X2 _add_514_U183  ( .A1(H2[26]), .A2(next_C[26]), .ZN(_add_514_n172 ) );
NOR2_X1 _add_514_U182  ( .A1(next_C[5]), .A2(H2[5]), .ZN(_add_514_n59 ) );
NOR2_X1 _add_514_U181  ( .A1(next_C[24]), .A2(H2[24]), .ZN(_add_514_n177 ));
NOR2_X1 _add_514_U180  ( .A1(next_C[7]), .A2(H2[7]), .ZN(_add_514_n51 ) );
NOR2_X1 _add_514_U179  ( .A1(next_C[1]), .A2(H2[1]), .ZN(_add_514_n117 ) );
NOR2_X1 _add_514_U178  ( .A1(next_C[16]), .A2(H2[16]), .ZN(_add_514_n248 ));
NOR2_X1 _add_514_U177  ( .A1(next_C[20]), .A2(H2[20]), .ZN(_add_514_n224 ));
NOR2_X1 _add_514_U176  ( .A1(next_C[8]), .A2(H2[8]), .ZN(_add_514_n42 ) );
AND2_X2 _add_514_U175  ( .A1(H2[10]), .A2(next_C[10]), .ZN(_add_514_n32 ) );
NAND3_X1 _add_514_U174  ( .A1(next_C[14]), .A2(H2[14]), .A3(_add_514_n271 ),.ZN(_add_514_n297 ) );
NAND3_X2 _add_514_U173  ( .A1(_add_514_n296 ), .A2(_add_514_n5 ), .A3(_add_514_n297 ), .ZN(_add_514_n136 ) );
AND4_X2 _add_514_U172  ( .A1(_add_514_n289 ), .A2(_add_514_n149 ), .A3(_add_514_n71 ), .A4(_add_514_n148 ), .ZN(_add_514_n31 ) );
NOR2_X1 _add_514_U171  ( .A1(next_C[14]), .A2(H2[14]), .ZN(_add_514_n294 ));
NOR2_X2 _add_514_U170  ( .A1(_add_514_n275 ), .A2(_add_514_n269 ), .ZN(_add_514_n293 ) );
NOR2_X2 _add_514_U169  ( .A1(_add_514_n270 ), .A2(_add_514_n294 ), .ZN(_add_514_n292 ) );
NOR2_X1 _add_514_U168  ( .A1(next_C[2]), .A2(H2[2]), .ZN(_add_514_n75 ) );
NOR2_X1 _add_514_U167  ( .A1(next_C[13]), .A2(H2[13]), .ZN(_add_514_n269 ));
NOR2_X1 _add_514_U166  ( .A1(next_C[14]), .A2(H2[14]), .ZN(_add_514_n272 ));
NOR2_X2 _add_514_U165  ( .A1(_add_514_n75 ), .A2(_add_514_n76 ), .ZN(_add_514_n72 ) );
AND2_X4 _add_514_U164  ( .A1(_add_514_n162 ), .A2(_add_514_n163 ), .ZN(_add_514_n30 ) );
NOR2_X2 _add_514_U163  ( .A1(_add_514_n241 ), .A2(_add_514_n117 ), .ZN(_add_514_n240 ) );
AND2_X2 _add_514_U162  ( .A1(_add_514_n96 ), .A2(_add_514_n95 ), .ZN(_add_514_n92 ) );
OR2_X4 _add_514_U161  ( .A1(_add_514_n101 ), .A2(_add_514_n110 ), .ZN(_add_514_n29 ) );
AND2_X2 _add_514_U160  ( .A1(_add_514_n96 ), .A2(_add_514_n29 ), .ZN(_add_514_n106 ) );
NAND3_X2 _add_514_U159  ( .A1(_add_514_n371 ), .A2(_add_514_n372 ), .A3(_add_514_n1 ), .ZN(_add_514_n291 ) );
OR2_X4 _add_514_U158  ( .A1(_add_514_n179 ), .A2(_add_514_n180 ), .ZN(_add_514_n28 ) );
XNOR2_X2 _add_514_U157  ( .A(_add_514_n28 ), .B(_add_514_n178 ), .ZN(N942));
NOR3_X2 _add_514_U156  ( .A1(_add_514_n278 ), .A2(_add_514_n279 ), .A3(_add_514_n64 ), .ZN(_add_514_n277 ) );
AND3_X2 _add_514_U155  ( .A1(_add_514_n4 ), .A2(_add_514_n125 ), .A3(_add_514_n126 ), .ZN(_add_514_n27 ) );
NOR2_X2 _add_514_U154  ( .A1(_add_514_n101 ), .A2(_add_514_n113 ), .ZN(_add_514_n112 ) );
NOR2_X2 _add_514_U153  ( .A1(_add_514_n101 ), .A2(_add_514_n114 ), .ZN(_add_514_n111 ) );
NOR2_X2 _add_514_U152  ( .A1(_add_514_n111 ), .A2(_add_514_n112 ), .ZN(_add_514_n104 ) );
NOR2_X2 _add_514_U151  ( .A1(_add_514_n275 ), .A2(_add_514_n269 ), .ZN(_add_514_n304 ) );
NOR2_X2 _add_514_U150  ( .A1(_add_514_n270 ), .A2(_add_514_n305 ), .ZN(_add_514_n303 ) );
NAND3_X2 _add_514_U149  ( .A1(_add_514_n303 ), .A2(_add_514_n301 ), .A3(_add_514_n304 ), .ZN(_add_514_n210 ) );
NOR2_X2 _add_514_U148  ( .A1(_add_514_n209 ), .A2(_add_514_n210 ), .ZN(_add_514_n295 ) );
NOR3_X2 _add_514_U147  ( .A1(_add_514_n295 ), .A2(_add_514_n151 ), .A3(_add_514_n136 ), .ZN(_add_514_n268 ) );
NAND3_X2 _add_514_U146  ( .A1(_add_514_n268 ), .A2(_add_514_n206 ), .A3(_add_514_n150 ), .ZN(_add_514_n247 ) );
NOR2_X2 _add_514_U145  ( .A1(_add_514_n327 ), .A2(_add_514_n348 ), .ZN(_add_514_n347 ) );
NAND3_X2 _add_514_U144  ( .A1(_add_514_n345 ), .A2(_add_514_n346 ), .A3(_add_514_n347 ), .ZN(_add_514_n146 ) );
NOR2_X2 _add_514_U143  ( .A1(_add_514_n272 ), .A2(_add_514_n309 ), .ZN(_add_514_n308 ) );
NAND3_X2 _add_514_U142  ( .A1(_add_514_n175 ), .A2(_add_514_n172 ), .A3(_add_514_n176 ), .ZN(_add_514_n167 ) );
NAND3_X2 _add_514_U141  ( .A1(_add_514_n222 ), .A2(_add_514_n218 ), .A3(_add_514_n223 ), .ZN(_add_514_n213 ) );
NOR3_X2 _add_514_U140  ( .A1(_add_514_n283 ), .A2(_add_514_n284 ), .A3(_add_514_n285 ), .ZN(_add_514_n281 ) );
NOR3_X2 _add_514_U139  ( .A1(_add_514_n183 ), .A2(_add_514_n184 ), .A3(_add_514_n185 ), .ZN(_add_514_n181 ) );
NOR2_X2 _add_514_U138  ( .A1(_add_514_n181 ), .A2(_add_514_n182 ), .ZN(_add_514_n179 ) );
NOR3_X2 _add_514_U137  ( .A1(_add_514_n260 ), .A2(_add_514_n250 ), .A3(_add_514_n248 ), .ZN(_add_514_n256 ) );
NOR3_X2 _add_514_U136  ( .A1(_add_514_n327 ), .A2(_add_514_n283 ), .A3(_add_514_n284 ), .ZN(_add_514_n326 ) );
NOR3_X2 _add_514_U135  ( .A1(_add_514_n248 ), .A2(_add_514_n249 ), .A3(_add_514_n250 ), .ZN(_add_514_n235 ) );
NOR2_X2 _add_514_U134  ( .A1(_add_514_n250 ), .A2(_add_514_n263 ), .ZN(_add_514_n262 ) );
XOR2_X2 _add_514_U133  ( .A(_add_514_n261 ), .B(_add_514_n262 ), .Z(N933) );
NOR2_X2 _add_514_U132  ( .A1(_add_514_n62 ), .A2(_add_514_n59 ), .ZN(_add_514_n61 ) );
NOR2_X2 _add_514_U131  ( .A1(_add_514_n34 ), .A2(_add_514_n39 ), .ZN(_add_514_n38 ) );
OR2_X4 _add_514_U130  ( .A1(_add_514_n256 ), .A2(_add_514_n254 ), .ZN(_add_514_n26 ) );
XNOR2_X2 _add_514_U129  ( .A(_add_514_n26 ), .B(_add_514_n255 ), .ZN(N934));
NOR2_X2 _add_514_U128  ( .A1(_add_514_n45 ), .A2(_add_514_n8 ), .ZN(_add_514_n40 ) );
NOR2_X2 _add_514_U127  ( .A1(_add_514_n42 ), .A2(_add_514_n43 ), .ZN(_add_514_n41 ) );
NOR2_X2 _add_514_U126  ( .A1(_add_514_n224 ), .A2(_add_514_n33 ), .ZN(_add_514_n231 ) );
NOR2_X2 _add_514_U125  ( .A1(_add_514_n177 ), .A2(_add_514_n195 ), .ZN(_add_514_n194 ) );
NOR2_X2 _add_514_U124  ( .A1(_add_514_n69 ), .A2(_add_514_n70 ), .ZN(_add_514_n68 ) );
NOR2_X2 _add_514_U123  ( .A1(_add_514_n72 ), .A2(_add_514_n73 ), .ZN(_add_514_n67 ) );
NOR2_X2 _add_514_U122  ( .A1(_add_514_n64 ), .A2(_add_514_n65 ), .ZN(_add_514_n66 ) );
NAND3_X2 _add_514_U121  ( .A1(_add_514_n154 ), .A2(_add_514_n153 ), .A3(_add_514_n7 ), .ZN(_add_514_n110 ) );
NOR2_X2 _add_514_U120  ( .A1(_add_514_n51 ), .A2(_add_514_n42 ), .ZN(_add_514_n377 ) );
OR2_X2 _add_514_U119  ( .A1(_add_514_n117 ), .A2(_add_514_n242 ), .ZN(_add_514_n25 ) );
NOR2_X2 _add_514_U118  ( .A1(_add_514_n365 ), .A2(_add_514_n366 ), .ZN(_add_514_n364 ) );
NAND3_X2 _add_514_U117  ( .A1(_add_514_n9 ), .A2(_add_514_n2 ), .A3(_add_514_n364 ), .ZN(_add_514_n47 ) );
NOR2_X2 _add_514_U116  ( .A1(_add_514_n100 ), .A2(_add_514_n101 ), .ZN(_add_514_n86 ) );
NOR2_X2 _add_514_U115  ( .A1(_add_514_n59 ), .A2(_add_514_n56 ), .ZN(_add_514_n333 ) );
NAND3_X2 _add_514_U114  ( .A1(_add_514_n301 ), .A2(_add_514_n271 ), .A3(_add_514_n302 ), .ZN(_add_514_n300 ) );
NOR2_X2 _add_514_U113  ( .A1(_add_514_n299 ), .A2(_add_514_n300 ), .ZN(_add_514_n151 ) );
NOR2_X2 _add_514_U112  ( .A1(_add_514_n94 ), .A2(_add_514_n85 ), .ZN(_add_514_n122 ) );
NAND3_X2 _add_514_U111  ( .A1(_add_514_n122 ), .A2(_add_514_n123 ), .A3(_add_514_n124 ), .ZN(_add_514_n118 ) );
NOR2_X2 _add_514_U110  ( .A1(_add_514_n209 ), .A2(_add_514_n305 ), .ZN(_add_514_n338 ) );
NOR2_X2 _add_514_U109  ( .A1(_add_514_n337 ), .A2(_add_514_n338 ), .ZN(_add_514_n335 ) );
NOR2_X2 _add_514_U108  ( .A1(_add_514_n312 ), .A2(_add_514_n270 ), .ZN(_add_514_n336 ) );
NOR2_X2 _add_514_U107  ( .A1(_add_514_n357 ), .A2(_add_514_n358 ), .ZN(_add_514_n356 ) );
NOR2_X2 _add_514_U106  ( .A1(_add_514_n356 ), .A2(_add_514_n32 ), .ZN(_add_514_n354 ) );
NOR2_X2 _add_514_U105  ( .A1(_add_514_n305 ), .A2(_add_514_n35 ), .ZN(_add_514_n355 ) );
NOR2_X2 _add_514_U104  ( .A1(_add_514_n34 ), .A2(_add_514_n359 ), .ZN(_add_514_n360 ) );
NOR2_X2 _add_514_U103  ( .A1(_add_514_n32 ), .A2(_add_514_n357 ), .ZN(_add_514_n361 ) );
OR2_X4 _add_514_U102  ( .A1(_add_514_n230 ), .A2(_add_514_n33 ), .ZN(_add_514_n24 ) );
XNOR2_X2 _add_514_U101  ( .A(_add_514_n24 ), .B(_add_514_n229 ), .ZN(N937));
OR2_X4 _add_514_U100  ( .A1(_add_514_n226 ), .A2(_add_514_n227 ), .ZN(_add_514_n23 ) );
XNOR2_X2 _add_514_U99  ( .A(_add_514_n23 ), .B(_add_514_n225 ), .ZN(N938) );
NOR2_X2 _add_514_U98  ( .A1(_add_514_n317 ), .A2(_add_514_n318 ), .ZN(_add_514_n314 ) );
NOR2_X2 _add_514_U97  ( .A1(_add_514_n316 ), .A2(_add_514_n272 ), .ZN(_add_514_n315 ) );
NOR2_X2 _add_514_U96  ( .A1(_add_514_n236 ), .A2(_add_514_n207 ), .ZN(_add_514_n234 ) );
NOR2_X2 _add_514_U95  ( .A1(_add_514_n234 ), .A2(_add_514_n131 ), .ZN(_add_514_n232 ) );
NOR2_X2 _add_514_U94  ( .A1(_add_514_n232 ), .A2(_add_514_n233 ), .ZN(_add_514_n221 ) );
NOR2_X2 _add_514_U93  ( .A1(_add_514_n34 ), .A2(_add_514_n359 ), .ZN(_add_514_n358 ) );
NOR2_X2 _add_514_U92  ( .A1(_add_514_n209 ), .A2(_add_514_n210 ), .ZN(_add_514_n208 ) );
NOR3_X2 _add_514_U91  ( .A1(_add_514_n208 ), .A2(_add_514_n151 ), .A3(_add_514_n136 ), .ZN(_add_514_n205 ) );
NAND3_X2 _add_514_U90  ( .A1(_add_514_n205 ), .A2(_add_514_n206 ), .A3(_add_514_n150 ), .ZN(_add_514_n189 ) );
OR2_X2 _add_514_U89  ( .A1(_add_514_n270 ), .A2(_add_514_n269 ), .ZN(_add_514_n22 ) );
NAND3_X2 _add_514_U88  ( .A1(_add_514_n155 ), .A2(_add_514_n154 ), .A3(_add_514_n165 ), .ZN(_add_514_n160 ) );
OR2_X4 _add_514_U87  ( .A1(_add_514_n130 ), .A2(_add_514_n131 ), .ZN(_add_514_n21 ) );
AND3_X2 _add_514_U86  ( .A1(_add_514_n152 ), .A2(_add_514_n21 ), .A3(_add_514_n129 ), .ZN(_add_514_n97 ) );
NOR2_X2 _add_514_U85  ( .A1(_add_514_n224 ), .A2(_add_514_n221 ), .ZN(_add_514_n230 ) );
NOR2_X2 _add_514_U84  ( .A1(_add_514_n32 ), .A2(_add_514_n35 ), .ZN(_add_514_n339 ) );
NAND3_X2 _add_514_U83  ( .A1(_add_514_n3 ), .A2(_add_514_n6 ), .A3(_add_514_n339 ), .ZN(_add_514_n138 ) );
NOR2_X2 _add_514_U82  ( .A1(_add_514_n312 ), .A2(_add_514_n313 ), .ZN(_add_514_n319 ) );
NOR2_X2 _add_514_U81  ( .A1(_add_514_n269 ), .A2(_add_514_n319 ), .ZN(_add_514_n317 ) );
OR3_X4 _add_514_U80  ( .A1(_add_514_n307 ), .A2(_add_514_n316 ), .A3(_add_514_n308 ), .ZN(_add_514_n20 ) );
XNOR2_X2 _add_514_U79  ( .A(_add_514_n20 ), .B(_add_514_n306 ), .ZN(N931) );
NOR2_X2 _add_514_U78  ( .A1(_add_514_n47 ), .A2(_add_514_n31 ), .ZN(_add_514_n288 ) );
NOR2_X2 _add_514_U77  ( .A1(_add_514_n146 ), .A2(_add_514_n147 ), .ZN(_add_514_n286 ) );
NAND3_X2 _add_514_U76  ( .A1(_add_514_n71 ), .A2(_add_514_n290 ), .A3(_add_514_n291 ), .ZN(_add_514_n287 ) );
NAND3_X2 _add_514_U75  ( .A1(_add_514_n286 ), .A2(_add_514_n287 ), .A3(_add_514_n288 ), .ZN(_add_514_n206 ) );
OR3_X2 _add_514_U74  ( .A1(_add_514_n275 ), .A2(_add_514_n51 ), .A3(_add_514_n42 ), .ZN(_add_514_n19 ) );
NOR3_X2 _add_514_U73  ( .A1(_add_514_n146 ), .A2(_add_514_n147 ), .A3(_add_514_n47 ), .ZN(_add_514_n145 ) );
NOR3_X2 _add_514_U72  ( .A1(_add_514_n221 ), .A2(_add_514_n228 ), .A3(_add_514_n224 ), .ZN(_add_514_n226 ) );
NAND3_X2 _add_514_U71  ( .A1(_add_514_n353 ), .A2(_add_514_n377 ), .A3(_add_514_n333 ), .ZN(_add_514_n376 ) );
NOR3_X2 _add_514_U70  ( .A1(_add_514_n46 ), .A2(_add_514_n47 ), .A3(_add_514_n42 ), .ZN(_add_514_n363 ) );
NAND3_X2 _add_514_U69  ( .A1(_add_514_n375 ), .A2(_add_514_n44 ), .A3(_add_514_n376 ), .ZN(_add_514_n362 ) );
NOR2_X2 _add_514_U68  ( .A1(_add_514_n362 ), .A2(_add_514_n363 ), .ZN(_add_514_n37 ) );
NOR2_X2 _add_514_U67  ( .A1(_add_514_n46 ), .A2(_add_514_n65 ), .ZN(_add_514_n63 ) );
NOR2_X2 _add_514_U66  ( .A1(_add_514_n63 ), .A2(_add_514_n64 ), .ZN(_add_514_n60 ) );
OR2_X4 _add_514_U65  ( .A1(_add_514_n215 ), .A2(_add_514_n216 ), .ZN(_add_514_n18 ) );
XNOR2_X2 _add_514_U64  ( .A(_add_514_n18 ), .B(_add_514_n214 ), .ZN(N939) );
OR2_X4 _add_514_U63  ( .A1(_add_514_n169 ), .A2(_add_514_n170 ), .ZN(_add_514_n17 ) );
XNOR2_X2 _add_514_U62  ( .A(_add_514_n17 ), .B(_add_514_n168 ), .ZN(N943) );
NOR2_X2 _add_514_U61  ( .A1(_add_514_n312 ), .A2(_add_514_n313 ), .ZN(_add_514_n320 ) );
NOR2_X2 _add_514_U60  ( .A1(_add_514_n318 ), .A2(_add_514_n269 ), .ZN(_add_514_n321 ) );
NOR2_X2 _add_514_U59  ( .A1(_add_514_n37 ), .A2(_add_514_n39 ), .ZN(_add_514_n359 ) );
OR2_X2 _add_514_U58  ( .A1(_add_514_n59 ), .A2(_add_514_n60 ), .ZN(_add_514_n16 ) );
NOR2_X2 _add_514_U57  ( .A1(_add_514_n312 ), .A2(_add_514_n313 ), .ZN(_add_514_n311 ) );
NOR3_X2 _add_514_U56  ( .A1(_add_514_n311 ), .A2(_add_514_n272 ), .A3(_add_514_n269 ), .ZN(_add_514_n307 ) );
NOR2_X2 _add_514_U55  ( .A1(_add_514_n373 ), .A2(_add_514_n374 ), .ZN(_add_514_n370 ) );
NOR3_X2 _add_514_U54  ( .A1(_add_514_n139 ), .A2(_add_514_n69 ), .A3(_add_514_n140 ), .ZN(_add_514_n133 ) );
NOR3_X2 _add_514_U53  ( .A1(_add_514_n132 ), .A2(_add_514_n133 ), .A3(_add_514_n134 ), .ZN(_add_514_n130 ) );
NOR2_X2 _add_514_U52  ( .A1(_add_514_n75 ), .A2(_add_514_n117 ), .ZN(_add_514_n141 ) );
NOR2_X2 _add_514_U51  ( .A1(_add_514_n141 ), .A2(_add_514_n142 ), .ZN(_add_514_n140 ) );
NOR3_X2 _add_514_U50  ( .A1(_add_514_n19 ), .A2(_add_514_n272 ), .A3(_add_514_n22 ), .ZN(_add_514_n274 ) );
NOR3_X2 _add_514_U49  ( .A1(_add_514_n276 ), .A2(_add_514_n277 ), .A3(_add_514_n11 ), .ZN(_add_514_n273 ) );
NOR2_X2 _add_514_U48  ( .A1(_add_514_n328 ), .A2(_add_514_n329 ), .ZN(_add_514_n322 ) );
NOR2_X2 _add_514_U47  ( .A1(_add_514_n326 ), .A2(_add_514_n138 ), .ZN(_add_514_n323 ) );
NOR3_X2 _add_514_U46  ( .A1(_add_514_n322 ), .A2(_add_514_n323 ), .A3(_add_514_n324 ), .ZN(_add_514_n313 ) );
NOR3_X2 _add_514_U45  ( .A1(_add_514_n75 ), .A2(_add_514_n369 ), .A3(_add_514_n69 ), .ZN(_add_514_n367 ) );
NOR3_X2 _add_514_U44  ( .A1(_add_514_n12 ), .A2(_add_514_n367 ), .A3(_add_514_n368 ), .ZN(_add_514_n46 ) );
NAND3_X2 _add_514_U43  ( .A1(_add_514_n333 ), .A2(_add_514_n334 ), .A3(_add_514_n2 ), .ZN(_add_514_n330 ) );
NAND3_X2 _add_514_U42  ( .A1(_add_514_n330 ), .A2(_add_514_n331 ), .A3(_add_514_n209 ), .ZN(_add_514_n328 ) );
NOR2_X2 _add_514_U41  ( .A1(_add_514_n46 ), .A2(_add_514_n47 ), .ZN(_add_514_n45 ) );
NOR2_X2 _add_514_U40  ( .A1(_add_514_n87 ), .A2(_add_514_n27 ), .ZN(_add_514_n124 ) );
NOR3_X2 _add_514_U39  ( .A1(_add_514_n188 ), .A2(_add_514_n99 ), .A3(_add_514_n131 ), .ZN(_add_514_n184 ) );
NAND3_X2 _add_514_U38  ( .A1(_add_514_n203 ), .A2(_add_514_n189 ), .A3(_add_514_n204 ), .ZN(_add_514_n202 ) );
NAND3_X2 _add_514_U37  ( .A1(_add_514_n4 ), .A2(_add_514_n203 ), .A3(_add_514_n108 ), .ZN(_add_514_n123 ) );
NOR2_X2 _add_514_U36  ( .A1(_add_514_n46 ), .A2(_add_514_n47 ), .ZN(_add_514_n349 ) );
NOR2_X2 _add_514_U35  ( .A1(_add_514_n349 ), .A2(_add_514_n8 ), .ZN(_add_514_n344 ) );
NOR2_X2 _add_514_U34  ( .A1(_add_514_n344 ), .A2(_add_514_n146 ), .ZN(_add_514_n337 ) );
NOR2_X2 _add_514_U33  ( .A1(_add_514_n166 ), .A2(_add_514_n167 ), .ZN(_add_514_n169 ) );
NOR2_X2 _add_514_U32  ( .A1(_add_514_n221 ), .A2(_add_514_n213 ), .ZN(_add_514_n215 ) );
NOR2_X2 _add_514_U31  ( .A1(_add_514_n46 ), .A2(_add_514_n47 ), .ZN(_add_514_n329 ) );
OR3_X2 _add_514_U30  ( .A1(_add_514_n97 ), .A2(_add_514_n98 ), .A3(_add_514_n99 ), .ZN(_add_514_n15 ) );
AND2_X4 _add_514_U29  ( .A1(_add_514_n190 ), .A2(_add_514_n202 ), .ZN(_add_514_n14 ) );
AND3_X2 _add_514_U28  ( .A1(_add_514_n14 ), .A2(_add_514_n186 ), .A3(_add_514_n187 ), .ZN(_add_514_n166 ) );
OR2_X4 _add_514_U27  ( .A1(next_C[0]), .A2(H2[0]), .ZN(_add_514_n36 ) );
OR2_X1 _add_514_U26  ( .A1(H2[17]), .A2(next_C[17]), .ZN(_add_514_n259 ) );
OR2_X1 _add_514_U25  ( .A1(H2[22]), .A2(next_C[22]), .ZN(_add_514_n218 ) );
OR2_X1 _add_514_U24  ( .A1(H2[30]), .A2(next_C[30]), .ZN(_add_514_n91 ) );
OR2_X1 _add_514_U23  ( .A1(H2[18]), .A2(next_C[18]), .ZN(_add_514_n251 ) );
OR2_X1 _add_514_U22  ( .A1(H2[19]), .A2(next_C[19]), .ZN(_add_514_n212 ) );
OR2_X1 _add_514_U21  ( .A1(H2[21]), .A2(next_C[21]), .ZN(_add_514_n222 ) );
OR2_X1 _add_514_U20  ( .A1(H2[23]), .A2(next_C[23]), .ZN(_add_514_n125 ) );
OR2_X1 _add_514_U19  ( .A1(H2[12]), .A2(next_C[12]), .ZN(_add_514_n325 ) );
OR2_X1 _add_514_U18  ( .A1(H2[15]), .A2(next_C[15]), .ZN(_add_514_n271 ) );
AND2_X4 _add_514_U17  ( .A1(_add_514_n242 ), .A2(_add_514_n36 ), .ZN(N916));
NAND2_X1 _add_514_U16  ( .A1(H2[14]), .A2(next_C[14]), .ZN(_add_514_n310 ));
NAND2_X1 _add_514_U15  ( .A1(H2[0]), .A2(next_C[0]), .ZN(_add_514_n242 ) );
AND4_X4 _add_514_U14  ( .A1(_add_514_n370 ), .A2(_add_514_n371 ), .A3(_add_514_n372 ), .A4(_add_514_n1 ), .ZN(_add_514_n12 ) );
AND3_X4 _add_514_U13  ( .A1(_add_514_n50 ), .A2(_add_514_n53 ), .A3(_add_514_n59 ), .ZN(_add_514_n11 ) );
OR2_X4 _add_514_U12  ( .A1(_add_514_n166 ), .A2(_add_514_n177 ), .ZN(_add_514_n10 ) );
OR2_X4 _add_514_U11  ( .A1(next_C[4]), .A2(H2[4]), .ZN(_add_514_n9 ) );
AND2_X4 _add_514_U10  ( .A1(_add_514_n350 ), .A2(_add_514_n2 ), .ZN(_add_514_n8 ) );
NAND2_X2 _add_514_U9  ( .A1(_add_514_n164 ), .A2(_add_514_n30 ), .ZN(_add_514_n7 ) );
OR2_X4 _add_514_U8  ( .A1(_add_514_n340 ), .A2(_add_514_n341 ), .ZN(_add_514_n6 ) );
OR2_X4 _add_514_U7  ( .A1(_add_514_n272 ), .A2(_add_514_n298 ), .ZN(_add_514_n5 ) );
AND3_X4 _add_514_U6  ( .A1(_add_514_n153 ), .A2(_add_514_n154 ), .A3(_add_514_n155 ), .ZN(_add_514_n4 ) );
OR3_X4 _add_514_U5  ( .A1(_add_514_n342 ), .A2(_add_514_n39 ), .A3(_add_514_n343 ), .ZN(_add_514_n3 ) );
OR2_X4 _add_514_U4  ( .A1(next_C[7]), .A2(H2[7]), .ZN(_add_514_n2 ) );
OR2_X4 _add_514_U3  ( .A1(next_C[2]), .A2(H2[2]), .ZN(_add_514_n1 ) );
XNOR2_X1 _add_514_U2  ( .A(H2[31]), .B(next_C[31]), .ZN(_add_514_n79 ) );
NAND2_X2 _add_513_U409  ( .A1(H1[0]), .A2(SHA1_result_128), .ZN(_add_513_n199 ) );
INV_X4 _add_513_U408  ( .A(H1[0]), .ZN(_add_513_n376 ) );
INV_X4 _add_513_U407  ( .A(SHA1_result_128), .ZN(_add_513_n377 ) );
NAND2_X2 _add_513_U406  ( .A1(_add_513_n376 ), .A2(_add_513_n377 ), .ZN(_add_513_n368 ) );
INV_X4 _add_513_U405  ( .A(_add_513_n29 ), .ZN(_add_513_n361 ) );
NAND2_X2 _add_513_U404  ( .A1(SHA1_result_134), .A2(H1[6]), .ZN(_add_513_n375 ) );
NAND2_X2 _add_513_U403  ( .A1(H1[4]), .A2(SHA1_result_132), .ZN(_add_513_n51 ) );
NAND2_X2 _add_513_U402  ( .A1(H1[5]), .A2(SHA1_result_133), .ZN(_add_513_n46 ) );
NAND2_X2 _add_513_U401  ( .A1(_add_513_n51 ), .A2(_add_513_n46 ), .ZN(_add_513_n283 ) );
NAND2_X2 _add_513_U400  ( .A1(_add_513_n283 ), .A2(_add_513_n374 ), .ZN(_add_513_n373 ) );
NAND2_X2 _add_513_U399  ( .A1(_add_513_n372 ), .A2(_add_513_n373 ), .ZN(_add_513_n34 ) );
NAND2_X2 _add_513_U398  ( .A1(_add_513_n32 ), .A2(_add_513_n34 ), .ZN(_add_513_n362 ) );
NAND2_X2 _add_513_U397  ( .A1(H1[8]), .A2(SHA1_result_136), .ZN(_add_513_n31 ) );
INV_X4 _add_513_U396  ( .A(_add_513_n53 ), .ZN(_add_513_n370 ) );
NAND2_X2 _add_513_U395  ( .A1(H1[1]), .A2(SHA1_result_129), .ZN(_add_513_n367 ) );
NAND2_X2 _add_513_U394  ( .A1(SHA1_result_130), .A2(H1[2]), .ZN(_add_513_n366 ) );
NAND2_X2 _add_513_U393  ( .A1(H1[3]), .A2(SHA1_result_131), .ZN(_add_513_n195 ) );
NAND2_X2 _add_513_U392  ( .A1(_add_513_n361 ), .A2(_add_513_n27 ), .ZN(_add_513_n360 ) );
NAND2_X2 _add_513_U391  ( .A1(H1[9]), .A2(n14443), .ZN(_add_513_n28 ) );
NAND2_X2 _add_513_U390  ( .A1(_add_513_n360 ), .A2(_add_513_n28 ), .ZN(_add_513_n358 ) );
NAND2_X2 _add_513_U389  ( .A1(H1[10]), .A2(n14440), .ZN(_add_513_n315 ) );
NAND2_X2 _add_513_U388  ( .A1(_add_513_n347 ), .A2(_add_513_n315 ), .ZN(_add_513_n359 ) );
XNOR2_X2 _add_513_U387  ( .A(_add_513_n358 ), .B(_add_513_n359 ), .ZN(N894));
INV_X4 _add_513_U386  ( .A(_add_513_n27 ), .ZN(_add_513_n357 ) );
NAND2_X2 _add_513_U385  ( .A1(_add_513_n357 ), .A2(_add_513_n28 ), .ZN(_add_513_n356 ) );
NAND2_X2 _add_513_U384  ( .A1(_add_513_n355 ), .A2(_add_513_n356 ), .ZN(_add_513_n354 ) );
NAND2_X2 _add_513_U383  ( .A1(_add_513_n354 ), .A2(_add_513_n315 ), .ZN(_add_513_n352 ) );
NAND2_X2 _add_513_U382  ( .A1(H1[11]), .A2(n14437), .ZN(_add_513_n313 ) );
NAND2_X2 _add_513_U381  ( .A1(_add_513_n313 ), .A2(_add_513_n202 ), .ZN(_add_513_n353 ) );
XNOR2_X2 _add_513_U380  ( .A(_add_513_n352 ), .B(_add_513_n353 ), .ZN(N895));
INV_X4 _add_513_U379  ( .A(_add_513_n54 ), .ZN(_add_513_n35 ) );
INV_X4 _add_513_U378  ( .A(_add_513_n350 ), .ZN(_add_513_n347 ) );
INV_X4 _add_513_U377  ( .A(_add_513_n32 ), .ZN(_add_513_n349 ) );
INV_X4 _add_513_U376  ( .A(_add_513_n315 ), .ZN(_add_513_n210 ) );
INV_X4 _add_513_U375  ( .A(_add_513_n313 ), .ZN(_add_513_n211 ) );
NAND2_X2 _add_513_U374  ( .A1(H1[9]), .A2(n14443), .ZN(_add_513_n345 ) );
NAND2_X2 _add_513_U373  ( .A1(_add_513_n31 ), .A2(_add_513_n345 ), .ZN(_add_513_n344 ) );
NAND2_X2 _add_513_U372  ( .A1(_add_513_n312 ), .A2(_add_513_n344 ), .ZN(_add_513_n343 ) );
NAND2_X2 _add_513_U371  ( .A1(_add_513_n342 ), .A2(_add_513_n343 ), .ZN(_add_513_n341 ) );
NAND2_X2 _add_513_U370  ( .A1(_add_513_n341 ), .A2(_add_513_n202 ), .ZN(_add_513_n336 ) );
INV_X4 _add_513_U369  ( .A(_add_513_n336 ), .ZN(_add_513_n338 ) );
NAND2_X2 _add_513_U368  ( .A1(H1[12]), .A2(n14434), .ZN(_add_513_n323 ) );
NAND2_X2 _add_513_U367  ( .A1(_add_513_n306 ), .A2(_add_513_n323 ), .ZN(_add_513_n339 ) );
INV_X4 _add_513_U366  ( .A(_add_513_n323 ), .ZN(_add_513_n288 ) );
NAND2_X2 _add_513_U365  ( .A1(_add_513_n194 ), .A2(_add_513_n336 ), .ZN(_add_513_n335 ) );
NAND2_X2 _add_513_U364  ( .A1(_add_513_n335 ), .A2(_add_513_n306 ), .ZN(_add_513_n334 ) );
NAND2_X2 _add_513_U363  ( .A1(H1[13]), .A2(n14431), .ZN(_add_513_n326 ) );
INV_X4 _add_513_U362  ( .A(_add_513_n326 ), .ZN(_add_513_n329 ) );
XNOR2_X2 _add_513_U361  ( .A(_add_513_n331 ), .B(_add_513_n332 ), .ZN(N897));
NAND2_X2 _add_513_U360  ( .A1(H1[14]), .A2(n14428), .ZN(_add_513_n292 ) );
NAND2_X2 _add_513_U359  ( .A1(_add_513_n292 ), .A2(_add_513_n294 ), .ZN(_add_513_n327 ) );
NAND2_X2 _add_513_U358  ( .A1(_add_513_n326 ), .A2(_add_513_n292 ), .ZN(_add_513_n325 ) );
NAND2_X2 _add_513_U357  ( .A1(_add_513_n325 ), .A2(_add_513_n294 ), .ZN(_add_513_n318 ) );
INV_X4 _add_513_U356  ( .A(_add_513_n294 ), .ZN(_add_513_n310 ) );
INV_X4 _add_513_U355  ( .A(_add_513_n324 ), .ZN(_add_513_n322 ) );
NAND2_X2 _add_513_U354  ( .A1(_add_513_n322 ), .A2(_add_513_n323 ), .ZN(_add_513_n321 ) );
NAND2_X2 _add_513_U353  ( .A1(_add_513_n320 ), .A2(_add_513_n321 ), .ZN(_add_513_n319 ) );
NAND2_X2 _add_513_U352  ( .A1(_add_513_n318 ), .A2(_add_513_n319 ), .ZN(_add_513_n316 ) );
NAND2_X2 _add_513_U351  ( .A1(H1[15]), .A2(n14425), .ZN(_add_513_n291 ) );
NAND2_X2 _add_513_U350  ( .A1(_add_513_n291 ), .A2(_add_513_n290 ), .ZN(_add_513_n317 ) );
XNOR2_X2 _add_513_U349  ( .A(_add_513_n316 ), .B(_add_513_n317 ), .ZN(N899));
NAND2_X2 _add_513_U348  ( .A1(H1[16]), .A2(n14422), .ZN(_add_513_n273 ) );
NAND2_X2 _add_513_U347  ( .A1(_add_513_n273 ), .A2(_add_513_n275 ), .ZN(_add_513_n276 ) );
NAND2_X2 _add_513_U346  ( .A1(H1[9]), .A2(n14443), .ZN(_add_513_n314 ) );
NAND4_X2 _add_513_U345  ( .A1(_add_513_n313 ), .A2(_add_513_n314 ), .A3(_add_513_n31 ), .A4(_add_513_n315 ), .ZN(_add_513_n303 ) );
INV_X4 _add_513_U344  ( .A(_add_513_n311 ), .ZN(_add_513_n307 ) );
INV_X4 _add_513_U343  ( .A(_add_513_n290 ), .ZN(_add_513_n309 ) );
INV_X4 _add_513_U342  ( .A(_add_513_n195 ), .ZN(_add_513_n59 ) );
NAND2_X2 _add_513_U341  ( .A1(H1[1]), .A2(SHA1_result_129), .ZN(_add_513_n298 ) );
INV_X4 _add_513_U340  ( .A(_add_513_n197 ), .ZN(_add_513_n299 ) );
NAND4_X2 _add_513_U339  ( .A1(_add_513_n199 ), .A2(_add_513_n298 ), .A3(_add_513_n195 ), .A4(_add_513_n299 ), .ZN(_add_513_n296 ) );
NAND4_X2 _add_513_U338  ( .A1(_add_513_n20 ), .A2(_add_513_n295 ), .A3(_add_513_n296 ), .A4(_add_513_n297 ), .ZN(_add_513_n278 ) );
INV_X4 _add_513_U337  ( .A(_add_513_n193 ), .ZN(_add_513_n286 ) );
INV_X4 _add_513_U336  ( .A(_add_513_n194 ), .ZN(_add_513_n287 ) );
NAND2_X2 _add_513_U335  ( .A1(_add_513_n289 ), .A2(_add_513_n290 ), .ZN(_add_513_n185 ) );
NAND2_X2 _add_513_U334  ( .A1(_add_513_n288 ), .A2(_add_513_n286 ), .ZN(_add_513_n189 ) );
NAND4_X2 _add_513_U333  ( .A1(_add_513_n282 ), .A2(_add_513_n283 ), .A3(_add_513_n287 ), .A4(_add_513_n284 ), .ZN(_add_513_n183 ) );
NAND2_X2 _add_513_U332  ( .A1(_add_513_n184 ), .A2(_add_513_n183 ), .ZN(_add_513_n281 ) );
XNOR2_X2 _add_513_U331  ( .A(_add_513_n276 ), .B(_add_513_n69 ), .ZN(N900));
INV_X4 _add_513_U330  ( .A(_add_513_n267 ), .ZN(_add_513_n275 ) );
NAND2_X2 _add_513_U329  ( .A1(_add_513_n69 ), .A2(_add_513_n275 ), .ZN(_add_513_n274 ) );
NAND2_X2 _add_513_U328  ( .A1(_add_513_n273 ), .A2(_add_513_n274 ), .ZN(_add_513_n270 ) );
INV_X4 _add_513_U327  ( .A(_add_513_n266 ), .ZN(_add_513_n272 ) );
NAND2_X2 _add_513_U326  ( .A1(H1[17]), .A2(n14419), .ZN(_add_513_n269 ) );
NAND2_X2 _add_513_U325  ( .A1(_add_513_n272 ), .A2(_add_513_n269 ), .ZN(_add_513_n271 ) );
XNOR2_X2 _add_513_U324  ( .A(_add_513_n270 ), .B(_add_513_n271 ), .ZN(N901));
NAND2_X2 _add_513_U323  ( .A1(_add_513_n268 ), .A2(_add_513_n269 ), .ZN(_add_513_n261 ) );
INV_X4 _add_513_U322  ( .A(_add_513_n261 ), .ZN(_add_513_n264 ) );
NAND2_X2 _add_513_U321  ( .A1(_add_513_n257 ), .A2(_add_513_n69 ), .ZN(_add_513_n265 ) );
NAND2_X2 _add_513_U320  ( .A1(_add_513_n264 ), .A2(_add_513_n265 ), .ZN(_add_513_n262 ) );
NAND2_X2 _add_513_U319  ( .A1(H1[18]), .A2(n14416), .ZN(_add_513_n260 ) );
NAND2_X2 _add_513_U318  ( .A1(_add_513_n258 ), .A2(_add_513_n260 ), .ZN(_add_513_n263 ) );
XNOR2_X2 _add_513_U317  ( .A(_add_513_n262 ), .B(_add_513_n263 ), .ZN(N902));
NAND2_X2 _add_513_U316  ( .A1(_add_513_n261 ), .A2(_add_513_n258 ), .ZN(_add_513_n259 ) );
NAND2_X2 _add_513_U315  ( .A1(_add_513_n259 ), .A2(_add_513_n260 ), .ZN(_add_513_n248 ) );
INV_X4 _add_513_U314  ( .A(_add_513_n248 ), .ZN(_add_513_n255 ) );
NAND2_X2 _add_513_U313  ( .A1(_add_513_n6 ), .A2(_add_513_n69 ), .ZN(_add_513_n256 ) );
NAND2_X2 _add_513_U312  ( .A1(_add_513_n255 ), .A2(_add_513_n256 ), .ZN(_add_513_n251 ) );
INV_X4 _add_513_U311  ( .A(H1[19]), .ZN(_add_513_n253 ) );
INV_X4 _add_513_U310  ( .A(n14413), .ZN(_add_513_n254 ) );
NAND2_X2 _add_513_U309  ( .A1(_add_513_n253 ), .A2(_add_513_n254 ), .ZN(_add_513_n247 ) );
NAND2_X2 _add_513_U308  ( .A1(H1[19]), .A2(n14413), .ZN(_add_513_n105 ) );
NAND2_X2 _add_513_U307  ( .A1(_add_513_n247 ), .A2(_add_513_n105 ), .ZN(_add_513_n252 ) );
XNOR2_X2 _add_513_U306  ( .A(_add_513_n251 ), .B(_add_513_n252 ), .ZN(N903));
NAND2_X2 _add_513_U305  ( .A1(H1[1]), .A2(SHA1_result_129), .ZN(_add_513_n116 ) );
INV_X4 _add_513_U304  ( .A(_add_513_n116 ), .ZN(_add_513_n250 ) );
XNOR2_X2 _add_513_U303  ( .A(_add_513_n199 ), .B(_add_513_n249 ), .ZN(N885));
NAND2_X2 _add_513_U302  ( .A1(_add_513_n248 ), .A2(_add_513_n247 ), .ZN(_add_513_n104 ) );
NAND2_X2 _add_513_U301  ( .A1(_add_513_n6 ), .A2(_add_513_n247 ), .ZN(_add_513_n128 ) );
INV_X4 _add_513_U300  ( .A(_add_513_n128 ), .ZN(_add_513_n68 ) );
NAND2_X2 _add_513_U299  ( .A1(_add_513_n68 ), .A2(_add_513_n69 ), .ZN(_add_513_n246 ) );
INV_X4 _add_513_U298  ( .A(H1[20]), .ZN(_add_513_n244 ) );
INV_X4 _add_513_U297  ( .A(SHA1_result_148), .ZN(_add_513_n245 ) );
NAND2_X2 _add_513_U296  ( .A1(_add_513_n244 ), .A2(_add_513_n245 ), .ZN(_add_513_n234 ) );
NAND2_X2 _add_513_U295  ( .A1(H1[20]), .A2(SHA1_result_148), .ZN(_add_513_n235 ) );
NAND2_X2 _add_513_U294  ( .A1(_add_513_n234 ), .A2(_add_513_n235 ), .ZN(_add_513_n243 ) );
XNOR2_X2 _add_513_U293  ( .A(_add_513_n225 ), .B(_add_513_n243 ), .ZN(N904));
NAND2_X2 _add_513_U292  ( .A1(_add_513_n225 ), .A2(_add_513_n234 ), .ZN(_add_513_n242 ) );
NAND2_X2 _add_513_U291  ( .A1(_add_513_n235 ), .A2(_add_513_n242 ), .ZN(_add_513_n238 ) );
NAND2_X2 _add_513_U290  ( .A1(H1[21]), .A2(n14408), .ZN(_add_513_n237 ) );
INV_X4 _add_513_U289  ( .A(H1[21]), .ZN(_add_513_n240 ) );
INV_X4 _add_513_U288  ( .A(n14408), .ZN(_add_513_n241 ) );
NAND2_X2 _add_513_U287  ( .A1(_add_513_n240 ), .A2(_add_513_n241 ), .ZN(_add_513_n236 ) );
NAND2_X2 _add_513_U286  ( .A1(_add_513_n237 ), .A2(_add_513_n236 ), .ZN(_add_513_n239 ) );
XNOR2_X2 _add_513_U285  ( .A(_add_513_n238 ), .B(_add_513_n239 ), .ZN(N905));
INV_X4 _add_513_U284  ( .A(_add_513_n237 ), .ZN(_add_513_n219 ) );
INV_X4 _add_513_U283  ( .A(_add_513_n236 ), .ZN(_add_513_n232 ) );
INV_X4 _add_513_U282  ( .A(_add_513_n234 ), .ZN(_add_513_n233 ) );
NAND2_X2 _add_513_U281  ( .A1(_add_513_n224 ), .A2(_add_513_n225 ), .ZN(_add_513_n231 ) );
NAND2_X2 _add_513_U280  ( .A1(_add_513_n230 ), .A2(_add_513_n231 ), .ZN(_add_513_n226 ) );
NAND2_X2 _add_513_U279  ( .A1(H1[22]), .A2(n14405), .ZN(_add_513_n221 ) );
INV_X4 _add_513_U278  ( .A(H1[22]), .ZN(_add_513_n228 ) );
INV_X4 _add_513_U277  ( .A(n14405), .ZN(_add_513_n229 ) );
NAND2_X2 _add_513_U276  ( .A1(_add_513_n228 ), .A2(_add_513_n229 ), .ZN(_add_513_n222 ) );
NAND2_X2 _add_513_U275  ( .A1(_add_513_n221 ), .A2(_add_513_n222 ), .ZN(_add_513_n227 ) );
XNOR2_X2 _add_513_U274  ( .A(_add_513_n226 ), .B(_add_513_n227 ), .ZN(N906));
INV_X4 _add_513_U273  ( .A(_add_513_n225 ), .ZN(_add_513_n223 ) );
NAND2_X2 _add_513_U272  ( .A1(_add_513_n224 ), .A2(_add_513_n222 ), .ZN(_add_513_n180 ) );
INV_X4 _add_513_U271  ( .A(_add_513_n222 ), .ZN(_add_513_n176 ) );
INV_X4 _add_513_U270  ( .A(_add_513_n221 ), .ZN(_add_513_n220 ) );
INV_X4 _add_513_U269  ( .A(H1[23]), .ZN(_add_513_n214 ) );
INV_X4 _add_513_U268  ( .A(SHA1_result_151), .ZN(_add_513_n215 ) );
NAND2_X2 _add_513_U267  ( .A1(_add_513_n214 ), .A2(_add_513_n215 ), .ZN(_add_513_n179 ) );
INV_X4 _add_513_U266  ( .A(_add_513_n179 ), .ZN(_add_513_n175 ) );
XNOR2_X2 _add_513_U265  ( .A(_add_513_n212 ), .B(_add_513_n213 ), .ZN(N907));
NAND2_X2 _add_513_U264  ( .A1(H1[9]), .A2(n14443), .ZN(_add_513_n207 ) );
NAND2_X2 _add_513_U263  ( .A1(_add_513_n31 ), .A2(_add_513_n207 ), .ZN(_add_513_n206 ) );
NAND2_X2 _add_513_U262  ( .A1(_add_513_n205 ), .A2(_add_513_n206 ), .ZN(_add_513_n204 ) );
NAND2_X2 _add_513_U261  ( .A1(_add_513_n203 ), .A2(_add_513_n204 ), .ZN(_add_513_n201 ) );
NAND2_X2 _add_513_U260  ( .A1(H1[1]), .A2(SHA1_result_129), .ZN(_add_513_n198 ) );
INV_X4 _add_513_U259  ( .A(_add_513_n36 ), .ZN(_add_513_n192 ) );
NAND4_X2 _add_513_U258  ( .A1(_add_513_n183 ), .A2(_add_513_n184 ), .A3(_add_513_n185 ), .A4(_add_513_n186 ), .ZN(_add_513_n182 ) );
INV_X4 _add_513_U257  ( .A(_add_513_n180 ), .ZN(_add_513_n178 ) );
NAND2_X2 _add_513_U256  ( .A1(_add_513_n178 ), .A2(_add_513_n179 ), .ZN(_add_513_n100 ) );
INV_X4 _add_513_U255  ( .A(_add_513_n104 ), .ZN(_add_513_n173 ) );
NAND2_X2 _add_513_U254  ( .A1(_add_513_n173 ), .A2(_add_513_n72 ), .ZN(_add_513_n172 ) );
NAND2_X2 _add_513_U253  ( .A1(_add_513_n171 ), .A2(_add_513_n172 ), .ZN(_add_513_n170 ) );
INV_X4 _add_513_U252  ( .A(H1[24]), .ZN(_add_513_n166 ) );
INV_X4 _add_513_U251  ( .A(n14400), .ZN(_add_513_n167 ) );
NAND2_X2 _add_513_U250  ( .A1(_add_513_n166 ), .A2(_add_513_n167 ), .ZN(_add_513_n148 ) );
INV_X4 _add_513_U249  ( .A(_add_513_n148 ), .ZN(_add_513_n159 ) );
NAND2_X2 _add_513_U248  ( .A1(H1[24]), .A2(n14400), .ZN(_add_513_n158 ) );
INV_X4 _add_513_U247  ( .A(_add_513_n158 ), .ZN(_add_513_n164 ) );
XNOR2_X2 _add_513_U246  ( .A(_add_513_n137 ), .B(_add_513_n165 ), .ZN(N908));
NAND2_X2 _add_513_U245  ( .A1(H1[25]), .A2(n14397), .ZN(_add_513_n157 ) );
INV_X4 _add_513_U244  ( .A(_add_513_n157 ), .ZN(_add_513_n162 ) );
XNOR2_X2 _add_513_U243  ( .A(_add_513_n160 ), .B(_add_513_n161 ), .ZN(N909));
NAND2_X2 _add_513_U242  ( .A1(_add_513_n157 ), .A2(_add_513_n158 ), .ZN(_add_513_n144 ) );
INV_X4 _add_513_U241  ( .A(_add_513_n144 ), .ZN(_add_513_n156 ) );
NAND2_X2 _add_513_U240  ( .A1(H1[26]), .A2(n14394), .ZN(_add_513_n136 ) );
INV_X4 _add_513_U239  ( .A(H1[26]), .ZN(_add_513_n152 ) );
INV_X4 _add_513_U238  ( .A(n14394), .ZN(_add_513_n153 ) );
NAND2_X2 _add_513_U237  ( .A1(_add_513_n152 ), .A2(_add_513_n153 ), .ZN(_add_513_n147 ) );
NAND2_X2 _add_513_U236  ( .A1(_add_513_n136 ), .A2(_add_513_n147 ), .ZN(_add_513_n151 ) );
INV_X4 _add_513_U235  ( .A(_add_513_n150 ), .ZN(_add_513_n149 ) );
INV_X4 _add_513_U234  ( .A(_add_513_n147 ), .ZN(_add_513_n145 ) );
NAND2_X2 _add_513_U233  ( .A1(_add_513_n143 ), .A2(_add_513_n144 ), .ZN(_add_513_n135 ) );
NAND2_X2 _add_513_U232  ( .A1(_add_513_n135 ), .A2(_add_513_n136 ), .ZN(_add_513_n142 ) );
NAND2_X2 _add_513_U231  ( .A1(H1[27]), .A2(n14391), .ZN(_add_513_n133 ) );
NAND2_X2 _add_513_U230  ( .A1(_add_513_n133 ), .A2(_add_513_n125 ), .ZN(_add_513_n140 ) );
INV_X4 _add_513_U229  ( .A(_add_513_n139 ), .ZN(_add_513_n126 ) );
NAND2_X2 _add_513_U228  ( .A1(_add_513_n126 ), .A2(_add_513_n125 ), .ZN(_add_513_n138 ) );
NAND2_X2 _add_513_U227  ( .A1(_add_513_n135 ), .A2(_add_513_n136 ), .ZN(_add_513_n134 ) );
NAND2_X2 _add_513_U226  ( .A1(_add_513_n134 ), .A2(_add_513_n125 ), .ZN(_add_513_n132 ) );
NAND2_X2 _add_513_U225  ( .A1(_add_513_n132 ), .A2(_add_513_n133 ), .ZN(_add_513_n89 ) );
NAND2_X2 _add_513_U224  ( .A1(H1[28]), .A2(n14388), .ZN(_add_513_n87 ) );
NAND2_X2 _add_513_U223  ( .A1(_add_513_n88 ), .A2(_add_513_n87 ), .ZN(_add_513_n130 ) );
INV_X4 _add_513_U222  ( .A(_add_513_n69 ), .ZN(_add_513_n129 ) );
NAND2_X2 _add_513_U221  ( .A1(_add_513_n104 ), .A2(_add_513_n105 ), .ZN(_add_513_n71 ) );
INV_X4 _add_513_U220  ( .A(_add_513_n100 ), .ZN(_add_513_n72 ) );
NAND2_X2 _add_513_U219  ( .A1(_add_513_n70 ), .A2(_add_513_n72 ), .ZN(_add_513_n124 ) );
NAND2_X2 _add_513_U218  ( .A1(_add_513_n89 ), .A2(_add_513_n88 ), .ZN(_add_513_n121 ) );
NAND2_X2 _add_513_U217  ( .A1(_add_513_n122 ), .A2(_add_513_n70 ), .ZN(_add_513_n113 ) );
NAND2_X2 _add_513_U216  ( .A1(_add_513_n121 ), .A2(_add_513_n113 ), .ZN(_add_513_n119 ) );
NAND2_X2 _add_513_U215  ( .A1(_add_513_n3 ), .A2(_add_513_n70 ), .ZN(_add_513_n112 ) );
NAND2_X2 _add_513_U214  ( .A1(_add_513_n112 ), .A2(_add_513_n87 ), .ZN(_add_513_n120 ) );
NAND2_X2 _add_513_U213  ( .A1(H1[29]), .A2(n14385), .ZN(_add_513_n81 ) );
NAND2_X2 _add_513_U212  ( .A1(_add_513_n81 ), .A2(_add_513_n108 ), .ZN(_add_513_n117 ) );
XNOR2_X2 _add_513_U211  ( .A(_add_513_n62 ), .B(_add_513_n114 ), .ZN(N886));
INV_X4 _add_513_U210  ( .A(_add_513_n113 ), .ZN(_add_513_n79 ) );
NAND2_X2 _add_513_U209  ( .A1(_add_513_n79 ), .A2(_add_513_n108 ), .ZN(_add_513_n110 ) );
INV_X4 _add_513_U208  ( .A(_add_513_n112 ), .ZN(_add_513_n90 ) );
NAND2_X2 _add_513_U207  ( .A1(_add_513_n90 ), .A2(_add_513_n108 ), .ZN(_add_513_n111 ) );
INV_X4 _add_513_U206  ( .A(_add_513_n81 ), .ZN(_add_513_n106 ) );
INV_X4 _add_513_U205  ( .A(_add_513_n108 ), .ZN(_add_513_n92 ) );
INV_X4 _add_513_U204  ( .A(_add_513_n105 ), .ZN(_add_513_n103 ) );
NAND2_X2 _add_513_U203  ( .A1(_add_513_n68 ), .A2(_add_513_n69 ), .ZN(_add_513_n102 ) );
NAND2_X2 _add_513_U202  ( .A1(_add_513_n101 ), .A2(_add_513_n102 ), .ZN(_add_513_n98 ) );
NAND2_X2 _add_513_U201  ( .A1(_add_513_n98 ), .A2(_add_513_n99 ), .ZN(_add_513_n97 ) );
NAND2_X2 _add_513_U200  ( .A1(H1[30]), .A2(n14382), .ZN(_add_513_n85 ) );
NAND2_X2 _add_513_U199  ( .A1(_add_513_n85 ), .A2(_add_513_n80 ), .ZN(_add_513_n94 ) );
XNOR2_X2 _add_513_U198  ( .A(_add_513_n93 ), .B(_add_513_n94 ), .ZN(N914) );
INV_X4 _add_513_U197  ( .A(_add_513_n80 ), .ZN(_add_513_n91 ) );
NAND2_X2 _add_513_U196  ( .A1(_add_513_n90 ), .A2(_add_513_n73 ), .ZN(_add_513_n82 ) );
INV_X4 _add_513_U195  ( .A(_add_513_n87 ), .ZN(_add_513_n86 ) );
NAND2_X2 _add_513_U194  ( .A1(_add_513_n86 ), .A2(_add_513_n73 ), .ZN(_add_513_n84 ) );
NAND4_X2 _add_513_U193  ( .A1(_add_513_n82 ), .A2(_add_513_n83 ), .A3(_add_513_n84 ), .A4(_add_513_n85 ), .ZN(_add_513_n75 ) );
NAND2_X2 _add_513_U192  ( .A1(_add_513_n106 ), .A2(_add_513_n80 ), .ZN(_add_513_n77 ) );
NAND2_X2 _add_513_U191  ( .A1(_add_513_n79 ), .A2(_add_513_n73 ), .ZN(_add_513_n78 ) );
NAND2_X2 _add_513_U190  ( .A1(_add_513_n77 ), .A2(_add_513_n78 ), .ZN(_add_513_n76 ) );
INV_X4 _add_513_U189  ( .A(_add_513_n74 ), .ZN(_add_513_n70 ) );
NAND4_X2 _add_513_U188  ( .A1(_add_513_n68 ), .A2(_add_513_n70 ), .A3(_add_513_n4 ), .A4(_add_513_n69 ), .ZN(_add_513_n67 ) );
XNOR2_X2 _add_513_U187  ( .A(H1[31]), .B(n14464), .ZN(_add_513_n64 ) );
XNOR2_X2 _add_513_U186  ( .A(_add_513_n63 ), .B(_add_513_n64 ), .ZN(N915) );
XNOR2_X2 _add_513_U185  ( .A(_add_513_n56 ), .B(_add_513_n57 ), .ZN(N887) );
NAND2_X2 _add_513_U184  ( .A1(_add_513_n53 ), .A2(_add_513_n51 ), .ZN(_add_513_n55 ) );
XNOR2_X2 _add_513_U183  ( .A(_add_513_n54 ), .B(_add_513_n55 ), .ZN(N888) );
NAND2_X2 _add_513_U182  ( .A1(_add_513_n46 ), .A2(_add_513_n48 ), .ZN(_add_513_n50 ) );
NAND2_X2 _add_513_U181  ( .A1(_add_513_n53 ), .A2(_add_513_n54 ), .ZN(_add_513_n52 ) );
NAND2_X2 _add_513_U180  ( .A1(_add_513_n51 ), .A2(_add_513_n52 ), .ZN(_add_513_n47 ) );
XNOR2_X2 _add_513_U179  ( .A(_add_513_n50 ), .B(_add_513_n47 ), .ZN(N889) );
NAND2_X2 _add_513_U178  ( .A1(H1[6]), .A2(SHA1_result_134), .ZN(_add_513_n40 ) );
NAND2_X2 _add_513_U177  ( .A1(_add_513_n40 ), .A2(_add_513_n1 ), .ZN(_add_513_n44 ) );
INV_X4 _add_513_U176  ( .A(_add_513_n49 ), .ZN(_add_513_n48 ) );
NAND2_X2 _add_513_U175  ( .A1(_add_513_n47 ), .A2(_add_513_n48 ), .ZN(_add_513_n45 ) );
NAND2_X2 _add_513_U174  ( .A1(_add_513_n45 ), .A2(_add_513_n46 ), .ZN(_add_513_n42 ) );
XNOR2_X2 _add_513_U173  ( .A(_add_513_n44 ), .B(_add_513_n42 ), .ZN(N890) );
NAND2_X2 _add_513_U172  ( .A1(_add_513_n42 ), .A2(_add_513_n1 ), .ZN(_add_513_n41 ) );
NAND2_X2 _add_513_U171  ( .A1(_add_513_n40 ), .A2(_add_513_n41 ), .ZN(_add_513_n37 ) );
NAND2_X2 _add_513_U170  ( .A1(_add_513_n31 ), .A2(_add_513_n32 ), .ZN(_add_513_n30 ) );
NAND2_X2 _add_513_U169  ( .A1(_add_513_n28 ), .A2(_add_513_n361 ), .ZN(_add_513_n26 ) );
XNOR2_X2 _add_513_U168  ( .A(_add_513_n26 ), .B(_add_513_n27 ), .ZN(N893) );
NAND2_X2 _add_513_U167  ( .A1(_add_513_n364 ), .A2(_add_513_n195 ), .ZN(_add_513_n54 ) );
NAND3_X2 _add_513_U166  ( .A1(_add_513_n70 ), .A2(_add_513_n4 ), .A3(_add_513_n71 ), .ZN(_add_513_n66 ) );
NAND3_X2 _add_513_U165  ( .A1(_add_513_n65 ), .A2(_add_513_n66 ), .A3(_add_513_n67 ), .ZN(_add_513_n63 ) );
AND2_X2 _add_513_U164  ( .A1(H1[2]), .A2(SHA1_result_130), .ZN(_add_513_n25 ) );
NOR2_X1 _add_513_U163  ( .A1(SHA1_result_133), .A2(H1[5]), .ZN(_add_513_n371 ) );
NOR2_X1 _add_513_U162  ( .A1(SHA1_result_130), .A2(H1[2]), .ZN(_add_513_n301 ) );
NOR2_X1 _add_513_U161  ( .A1(SHA1_result_129), .A2(H1[1]), .ZN(_add_513_n302 ) );
AND2_X2 _add_513_U160  ( .A1(H1[7]), .A2(SHA1_result_135), .ZN(_add_513_n24 ) );
NOR2_X2 _add_513_U159  ( .A1(n14419), .A2(H1[17]), .ZN(_add_513_n266 ) );
NAND3_X2 _add_513_U158  ( .A1(n14422), .A2(_add_513_n272 ), .A3(H1[16]),.ZN(_add_513_n268 ) );
NOR2_X1 _add_513_U157  ( .A1(n14440), .A2(H1[10]), .ZN(_add_513_n209 ) );
AND2_X4 _add_513_U156  ( .A1(_add_513_n198 ), .A2(_add_513_n199 ), .ZN(_add_513_n23 ) );
OR2_X2 _add_513_U155  ( .A1(_add_513_n200 ), .A2(_add_513_n23 ), .ZN(_add_513_n196 ) );
NOR2_X1 _add_513_U154  ( .A1(SHA1_result_131), .A2(H1[3]), .ZN(_add_513_n58 ) );
NOR2_X1 _add_513_U153  ( .A1(SHA1_result_130), .A2(H1[2]), .ZN(_add_513_n61 ) );
NOR2_X1 _add_513_U152  ( .A1(n14443), .A2(H1[9]), .ZN(_add_513_n208 ) );
NOR2_X1 _add_513_U151  ( .A1(SHA1_result_129), .A2(H1[1]), .ZN(_add_513_n115 ) );
OR2_X2 _add_513_U150  ( .A1(H1[18]), .A2(n14416), .ZN(_add_513_n258 ) );
NOR2_X2 _add_513_U149  ( .A1(_add_513_n39 ), .A2(_add_513_n375 ), .ZN(_add_513_n285 ) );
NOR2_X1 _add_513_U148  ( .A1(n14440), .A2(H1[10]), .ZN(_add_513_n350 ) );
NOR2_X2 _add_513_U147  ( .A1(n14422), .A2(H1[16]), .ZN(_add_513_n267 ) );
NAND3_X2 _add_513_U146  ( .A1(_add_513_n291 ), .A2(_add_513_n292 ), .A3(_add_513_n293 ), .ZN(_add_513_n289 ) );
NOR2_X2 _add_513_U145  ( .A1(H1[25]), .A2(n14397), .ZN(_add_513_n146 ) );
NOR2_X2 _add_513_U144  ( .A1(H1[25]), .A2(n14397), .ZN(_add_513_n150 ) );
NOR2_X2 _add_513_U143  ( .A1(_add_513_n58 ), .A2(_add_513_n366 ), .ZN(_add_513_n197 ) );
NOR2_X1 _add_513_U142  ( .A1(SHA1_result_133), .A2(H1[5]), .ZN(_add_513_n49 ) );
NOR2_X1 _add_513_U141  ( .A1(SHA1_result_134), .A2(H1[6]), .ZN(_add_513_n43 ) );
NOR2_X1 _add_513_U140  ( .A1(SHA1_result_135), .A2(H1[7]), .ZN(_add_513_n39 ) );
OR2_X2 _add_513_U139  ( .A1(H1[15]), .A2(n14425), .ZN(_add_513_n290 ) );
NOR2_X1 _add_513_U138  ( .A1(n14443), .A2(H1[9]), .ZN(_add_513_n29 ) );
OR2_X2 _add_513_U137  ( .A1(H1[14]), .A2(n14428), .ZN(_add_513_n294 ) );
NOR2_X2 _add_513_U136  ( .A1(_add_513_n146 ), .A2(_add_513_n156 ), .ZN(_add_513_n155 ) );
NOR2_X2 _add_513_U135  ( .A1(_add_513_n3 ), .A2(_add_513_n122 ), .ZN(_add_513_n171 ) );
NAND3_X2 _add_513_U134  ( .A1(_add_513_n195 ), .A2(_add_513_n196 ), .A3(_add_513_n299 ), .ZN(_add_513_n190 ) );
NOR2_X2 _add_513_U133  ( .A1(_add_513_n193 ), .A2(_add_513_n194 ), .ZN(_add_513_n191 ) );
NAND3_X2 _add_513_U132  ( .A1(_add_513_n190 ), .A2(_add_513_n191 ), .A3(_add_513_n192 ), .ZN(_add_513_n188 ) );
NAND3_X2 _add_513_U131  ( .A1(_add_513_n5 ), .A2(_add_513_n8 ), .A3(_add_513_n2 ), .ZN(_add_513_n200 ) );
NAND3_X2 _add_513_U130  ( .A1(_add_513_n285 ), .A2(_add_513_n286 ), .A3(_add_513_n287 ), .ZN(_add_513_n184 ) );
NOR2_X2 _add_513_U129  ( .A1(_add_513_n61 ), .A2(_add_513_n62 ), .ZN(_add_513_n60 ) );
NOR2_X2 _add_513_U128  ( .A1(_add_513_n60 ), .A2(_add_513_n25 ), .ZN(_add_513_n56 ) );
NOR2_X2 _add_513_U127  ( .A1(_add_513_n58 ), .A2(_add_513_n59 ), .ZN(_add_513_n57 ) );
OR2_X4 _add_513_U126  ( .A1(_add_513_n340 ), .A2(_add_513_n338 ), .ZN(_add_513_n22 ) );
XNOR2_X2 _add_513_U125  ( .A(_add_513_n22 ), .B(_add_513_n339 ), .ZN(N896));
OR2_X4 _add_513_U124  ( .A1(_add_513_n301 ), .A2(_add_513_n302 ), .ZN(_add_513_n21 ) );
NAND2_X2 _add_513_U123  ( .A1(_add_513_n21 ), .A2(_add_513_n300 ), .ZN(_add_513_n20 ) );
OR2_X4 _add_513_U122  ( .A1(_add_513_n328 ), .A2(_add_513_n329 ), .ZN(_add_513_n19 ) );
XNOR2_X2 _add_513_U121  ( .A(_add_513_n19 ), .B(_add_513_n327 ), .ZN(N898));
NOR2_X2 _add_513_U120  ( .A1(_add_513_n310 ), .A2(_add_513_n311 ), .ZN(_add_513_n320 ) );
NOR2_X2 _add_513_U119  ( .A1(_add_513_n197 ), .A2(_add_513_n59 ), .ZN(_add_513_n300 ) );
NOR2_X2 _add_513_U118  ( .A1(_add_513_n29 ), .A2(_add_513_n350 ), .ZN(_add_513_n355 ) );
OR2_X4 _add_513_U117  ( .A1(_add_513_n33 ), .A2(_add_513_n34 ), .ZN(_add_513_n18 ) );
XNOR2_X2 _add_513_U116  ( .A(_add_513_n18 ), .B(_add_513_n30 ), .ZN(N892) );
NAND3_X2 _add_513_U115  ( .A1(_add_513_n24 ), .A2(_add_513_n286 ), .A3(_add_513_n287 ), .ZN(_add_513_n186 ) );
OR2_X4 _add_513_U114  ( .A1(_add_513_n131 ), .A2(_add_513_n89 ), .ZN(_add_513_n17 ) );
XNOR2_X2 _add_513_U113  ( .A(_add_513_n17 ), .B(_add_513_n130 ), .ZN(N912));
NAND3_X2 _add_513_U112  ( .A1(_add_513_n201 ), .A2(_add_513_n202 ), .A3(_add_513_n286 ), .ZN(_add_513_n187 ) );
NAND3_X2 _add_513_U111  ( .A1(_add_513_n188 ), .A2(_add_513_n189 ), .A3(_add_513_n187 ), .ZN(_add_513_n181 ) );
NOR2_X2 _add_513_U110  ( .A1(_add_513_n181 ), .A2(_add_513_n182 ), .ZN(_add_513_n177 ) );
NOR2_X2 _add_513_U109  ( .A1(_add_513_n137 ), .A2(_add_513_n138 ), .ZN(_add_513_n131 ) );
NAND3_X2 _add_513_U108  ( .A1(_add_513_n148 ), .A2(_add_513_n147 ), .A3(_add_513_n149 ), .ZN(_add_513_n139 ) );
NOR2_X2 _add_513_U107  ( .A1(_add_513_n266 ), .A2(_add_513_n267 ), .ZN(_add_513_n257 ) );
NOR2_X2 _add_513_U106  ( .A1(_add_513_n288 ), .A2(_add_513_n324 ), .ZN(_add_513_n330 ) );
NOR2_X2 _add_513_U105  ( .A1(_add_513_n311 ), .A2(_add_513_n330 ), .ZN(_add_513_n328 ) );
NOR2_X2 _add_513_U104  ( .A1(_add_513_n39 ), .A2(_add_513_n24 ), .ZN(_add_513_n38 ) );
XOR2_X2 _add_513_U103  ( .A(_add_513_n37 ), .B(_add_513_n38 ), .Z(N891) );
NOR2_X2 _add_513_U102  ( .A1(_add_513_n92 ), .A2(_add_513_n87 ), .ZN(_add_513_n107 ) );
NAND3_X2 _add_513_U101  ( .A1(_add_513_n73 ), .A2(_add_513_n88 ), .A3(_add_513_n89 ), .ZN(_add_513_n83 ) );
NAND3_X2 _add_513_U100  ( .A1(_add_513_n32 ), .A2(_add_513_n192 ), .A3(_add_513_n54 ), .ZN(_add_513_n363 ) );
NAND3_X2 _add_513_U99  ( .A1(_add_513_n362 ), .A2(_add_513_n31 ), .A3(_add_513_n363 ), .ZN(_add_513_n27 ) );
NAND3_X2 _add_513_U98  ( .A1(_add_513_n88 ), .A2(_add_513_n108 ), .A3(_add_513_n89 ), .ZN(_add_513_n109 ) );
AND2_X4 _add_513_U97  ( .A1(_add_513_n110 ), .A2(_add_513_n111 ), .ZN(_add_513_n16 ) );
AND2_X2 _add_513_U96  ( .A1(_add_513_n16 ), .A2(_add_513_n109 ), .ZN(_add_513_n95 ) );
NOR2_X2 _add_513_U95  ( .A1(_add_513_n145 ), .A2(_add_513_n146 ), .ZN(_add_513_n143 ) );
NOR2_X2 _add_513_U94  ( .A1(_add_513_n208 ), .A2(_add_513_n209 ), .ZN(_add_513_n312 ) );
OR2_X4 _add_513_U93  ( .A1(_add_513_n115 ), .A2(_add_513_n199 ), .ZN(_add_513_n15 ) );
AND2_X2 _add_513_U92  ( .A1(_add_513_n116 ), .A2(_add_513_n15 ), .ZN(_add_513_n62 ) );
NAND3_X2 _add_513_U91  ( .A1(_add_513_n125 ), .A2(_add_513_n88 ), .A3(_add_513_n126 ), .ZN(_add_513_n74 ) );
NOR2_X2 _add_513_U90  ( .A1(_add_513_n106 ), .A2(_add_513_n107 ), .ZN(_add_513_n96 ) );
NAND3_X2 _add_513_U89  ( .A1(_add_513_n95 ), .A2(_add_513_n96 ), .A3(_add_513_n97 ), .ZN(_add_513_n93 ) );
NOR2_X2 _add_513_U88  ( .A1(_add_513_n288 ), .A2(_add_513_n324 ), .ZN(_add_513_n331 ) );
NOR2_X2 _add_513_U87  ( .A1(_add_513_n329 ), .A2(_add_513_n311 ), .ZN(_add_513_n332 ) );
OR3_X4 _add_513_U86  ( .A1(_add_513_n118 ), .A2(_add_513_n119 ), .A3(_add_513_n120 ), .ZN(_add_513_n14 ) );
XNOR2_X2 _add_513_U85  ( .A(_add_513_n14 ), .B(_add_513_n117 ), .ZN(N913) );
NOR2_X2 _add_513_U84  ( .A1(_add_513_n25 ), .A2(_add_513_n61 ), .ZN(_add_513_n114 ) );
OR2_X4 _add_513_U83  ( .A1(_add_513_n141 ), .A2(_add_513_n142 ), .ZN(_add_513_n13 ) );
XNOR2_X2 _add_513_U82  ( .A(_add_513_n13 ), .B(_add_513_n140 ), .ZN(N911) );
NOR2_X2 _add_513_U81  ( .A1(_add_513_n250 ), .A2(_add_513_n115 ), .ZN(_add_513_n249 ) );
NOR2_X2 _add_513_U80  ( .A1(_add_513_n208 ), .A2(_add_513_n209 ), .ZN(_add_513_n205 ) );
NOR2_X2 _add_513_U79  ( .A1(_add_513_n210 ), .A2(_add_513_n211 ), .ZN(_add_513_n203 ) );
NOR2_X2 _add_513_U78  ( .A1(_add_513_n210 ), .A2(_add_513_n211 ), .ZN(_add_513_n342 ) );
NOR2_X2 _add_513_U77  ( .A1(_add_513_n232 ), .A2(_add_513_n235 ), .ZN(_add_513_n218 ) );
NOR2_X2 _add_513_U76  ( .A1(_add_513_n370 ), .A2(_add_513_n371 ), .ZN(_add_513_n369 ) );
NAND3_X2 _add_513_U75  ( .A1(_add_513_n7 ), .A2(_add_513_n1 ), .A3(_add_513_n369 ), .ZN(_add_513_n36 ) );
NOR3_X2 _add_513_U74  ( .A1(_add_513_n337 ), .A2(_add_513_n338 ), .A3(_add_513_n34 ), .ZN(_add_513_n333 ) );
NOR2_X2 _add_513_U73  ( .A1(_add_513_n333 ), .A2(_add_513_n334 ), .ZN(_add_513_n324 ) );
NOR2_X2 _add_513_U72  ( .A1(_add_513_n75 ), .A2(_add_513_n76 ), .ZN(_add_513_n65 ) );
NOR3_X2 _add_513_U71  ( .A1(_add_513_n218 ), .A2(_add_513_n219 ), .A3(_add_513_n220 ), .ZN(_add_513_n174 ) );
NOR2_X2 _add_513_U70  ( .A1(_add_513_n91 ), .A2(_add_513_n92 ), .ZN(_add_513_n73 ) );
NOR2_X2 _add_513_U69  ( .A1(_add_513_n10 ), .A2(_add_513_n200 ), .ZN(_add_513_n365 ) );
NOR2_X2 _add_513_U68  ( .A1(_add_513_n365 ), .A2(_add_513_n197 ), .ZN(_add_513_n364 ) );
NOR3_X2 _add_513_U67  ( .A1(_add_513_n49 ), .A2(_add_513_n43 ), .A3(_add_513_n39 ), .ZN(_add_513_n374 ) );
NOR2_X2 _add_513_U66  ( .A1(_add_513_n24 ), .A2(_add_513_n285 ), .ZN(_add_513_n372 ) );
NAND3_X2 _add_513_U65  ( .A1(_add_513_n185 ), .A2(_add_513_n189 ), .A3(_add_513_n186 ), .ZN(_add_513_n280 ) );
NOR2_X2 _add_513_U64  ( .A1(_add_513_n39 ), .A2(_add_513_n193 ), .ZN(_add_513_n284 ) );
NOR2_X2 _add_513_U63  ( .A1(_add_513_n43 ), .A2(_add_513_n49 ), .ZN(_add_513_n282 ) );
OR2_X4 _add_513_U62  ( .A1(_add_513_n154 ), .A2(_add_513_n155 ), .ZN(_add_513_n12 ) );
XNOR2_X2 _add_513_U61  ( .A(_add_513_n12 ), .B(_add_513_n151 ), .ZN(N910) );
NOR2_X2 _add_513_U60  ( .A1(_add_513_n163 ), .A2(_add_513_n164 ), .ZN(_add_513_n160 ) );
NOR2_X2 _add_513_U59  ( .A1(_add_513_n150 ), .A2(_add_513_n162 ), .ZN(_add_513_n161 ) );
NOR2_X2 _add_513_U58  ( .A1(_add_513_n232 ), .A2(_add_513_n233 ), .ZN(_add_513_n224 ) );
NOR2_X2 _add_513_U57  ( .A1(_add_513_n219 ), .A2(_add_513_n218 ), .ZN(_add_513_n230 ) );
NOR3_X2 _add_513_U56  ( .A1(_add_513_n137 ), .A2(_add_513_n150 ), .A3(_add_513_n159 ), .ZN(_add_513_n154 ) );
NOR2_X2 _add_513_U55  ( .A1(_add_513_n280 ), .A2(_add_513_n281 ), .ZN(_add_513_n279 ) );
NAND3_X2 _add_513_U54  ( .A1(_add_513_n202 ), .A2(_add_513_n303 ), .A3(_add_513_n304 ), .ZN(_add_513_n277 ) );
NAND3_X2 _add_513_U53  ( .A1(_add_513_n277 ), .A2(_add_513_n278 ), .A3(_add_513_n279 ), .ZN(_add_513_n69 ) );
NAND3_X2 _add_513_U52  ( .A1(_add_513_n104 ), .A2(_add_513_n105 ), .A3(_add_513_n246 ), .ZN(_add_513_n225 ) );
NOR2_X2 _add_513_U51  ( .A1(_add_513_n309 ), .A2(_add_513_n310 ), .ZN(_add_513_n308 ) );
NAND3_X2 _add_513_U50  ( .A1(_add_513_n306 ), .A2(_add_513_n307 ), .A3(_add_513_n308 ), .ZN(_add_513_n193 ) );
NOR2_X2 _add_513_U49  ( .A1(_add_513_n349 ), .A2(_add_513_n29 ), .ZN(_add_513_n348 ) );
NAND3_X2 _add_513_U48  ( .A1(_add_513_n202 ), .A2(_add_513_n347 ), .A3(_add_513_n348 ), .ZN(_add_513_n194 ) );
NOR2_X2 _add_513_U47  ( .A1(_add_513_n177 ), .A2(_add_513_n11 ), .ZN(_add_513_n168 ) );
NOR2_X2 _add_513_U46  ( .A1(_add_513_n100 ), .A2(_add_513_n105 ), .ZN(_add_513_n169 ) );
NOR3_X2 _add_513_U45  ( .A1(_add_513_n168 ), .A2(_add_513_n169 ), .A3(_add_513_n170 ), .ZN(_add_513_n137 ) );
OR2_X2 _add_513_U44  ( .A1(_add_513_n128 ), .A2(_add_513_n100 ), .ZN(_add_513_n11 ) );
NOR2_X2 _add_513_U43  ( .A1(_add_513_n137 ), .A2(_add_513_n139 ), .ZN(_add_513_n141 ) );
NOR2_X2 _add_513_U42  ( .A1(_add_513_n35 ), .A2(_add_513_n36 ), .ZN(_add_513_n33 ) );
NOR2_X2 _add_513_U41  ( .A1(_add_513_n35 ), .A2(_add_513_n36 ), .ZN(_add_513_n351 ) );
NOR2_X2 _add_513_U40  ( .A1(_add_513_n351 ), .A2(_add_513_n34 ), .ZN(_add_513_n346 ) );
NOR2_X2 _add_513_U39  ( .A1(_add_513_n346 ), .A2(_add_513_n194 ), .ZN(_add_513_n340 ) );
NOR2_X2 _add_513_U38  ( .A1(_add_513_n128 ), .A2(_add_513_n129 ), .ZN(_add_513_n127 ) );
NOR2_X2 _add_513_U37  ( .A1(_add_513_n127 ), .A2(_add_513_n71 ), .ZN(_add_513_n123 ) );
NOR2_X2 _add_513_U36  ( .A1(_add_513_n123 ), .A2(_add_513_n124 ), .ZN(_add_513_n118 ) );
NOR2_X2 _add_513_U35  ( .A1(_add_513_n35 ), .A2(_add_513_n36 ), .ZN(_add_513_n337 ) );
NOR3_X2 _add_513_U34  ( .A1(_add_513_n193 ), .A2(_add_513_n194 ), .A3(_add_513_n36 ), .ZN(_add_513_n297 ) );
NOR3_X2 _add_513_U33  ( .A1(_add_513_n211 ), .A2(_add_513_n312 ), .A3(_add_513_n210 ), .ZN(_add_513_n305 ) );
NOR2_X2 _add_513_U32  ( .A1(_add_513_n305 ), .A2(_add_513_n193 ), .ZN(_add_513_n304 ) );
NOR2_X2 _add_513_U31  ( .A1(_add_513_n159 ), .A2(_add_513_n164 ), .ZN(_add_513_n165 ) );
NOR2_X2 _add_513_U30  ( .A1(_add_513_n103 ), .A2(_add_513_n173 ), .ZN(_add_513_n101 ) );
NOR3_X2 _add_513_U29  ( .A1(_add_513_n92 ), .A2(_add_513_n100 ), .A3(_add_513_n74 ), .ZN(_add_513_n99 ) );
NOR3_X2 _add_513_U28  ( .A1(_add_513_n174 ), .A2(_add_513_n175 ), .A3(_add_513_n176 ), .ZN(_add_513_n122 ) );
NOR2_X2 _add_513_U27  ( .A1(_add_513_n176 ), .A2(_add_513_n174 ), .ZN(_add_513_n217 ) );
NOR2_X2 _add_513_U26  ( .A1(_add_513_n216 ), .A2(_add_513_n217 ), .ZN(_add_513_n212 ) );
NOR2_X2 _add_513_U25  ( .A1(_add_513_n175 ), .A2(_add_513_n3 ), .ZN(_add_513_n213 ) );
NOR2_X2 _add_513_U24  ( .A1(_add_513_n223 ), .A2(_add_513_n180 ), .ZN(_add_513_n216 ) );
NOR2_X2 _add_513_U23  ( .A1(_add_513_n159 ), .A2(_add_513_n137 ), .ZN(_add_513_n163 ) );
OR2_X1 _add_513_U22  ( .A1(H1[3]), .A2(SHA1_result_131), .ZN(_add_513_n295 ));
OR2_X1 _add_513_U21  ( .A1(H1[30]), .A2(n14382), .ZN(_add_513_n80 ) );
OR2_X1 _add_513_U20  ( .A1(H1[27]), .A2(n14391), .ZN(_add_513_n125 ) );
OR2_X1 _add_513_U19  ( .A1(H1[28]), .A2(n14388), .ZN(_add_513_n88 ) );
OR2_X1 _add_513_U18  ( .A1(H1[29]), .A2(n14385), .ZN(_add_513_n108 ) );
OR2_X1 _add_513_U17  ( .A1(H1[4]), .A2(SHA1_result_132), .ZN(_add_513_n53 ));
OR2_X1 _add_513_U16  ( .A1(H1[8]), .A2(SHA1_result_136), .ZN(_add_513_n32 ));
NAND3_X1 _add_513_U15  ( .A1(n14431), .A2(H1[13]), .A3(_add_513_n294 ), .ZN(_add_513_n293 ) );
OR2_X1 _add_513_U14  ( .A1(H1[12]), .A2(n14434), .ZN(_add_513_n306 ) );
OR2_X1 _add_513_U13  ( .A1(H1[11]), .A2(n14437), .ZN(_add_513_n202 ) );
NOR2_X1 _add_513_U12  ( .A1(n14431), .A2(H1[13]), .ZN(_add_513_n311 ) );
AND2_X4 _add_513_U11  ( .A1(_add_513_n367 ), .A2(_add_513_n199 ), .ZN(_add_513_n10 ) );
AND2_X4 _add_513_U10  ( .A1(_add_513_n199 ), .A2(_add_513_n368 ), .ZN(N884));
OR2_X4 _add_513_U9  ( .A1(SHA1_result_131), .A2(H1[3]), .ZN(_add_513_n8 ) );
OR2_X4 _add_513_U8  ( .A1(SHA1_result_135), .A2(H1[7]), .ZN(_add_513_n7 ) );
AND2_X4 _add_513_U7  ( .A1(_add_513_n257 ), .A2(_add_513_n258 ), .ZN(_add_513_n6 ) );
OR2_X4 _add_513_U6  ( .A1(SHA1_result_130), .A2(H1[2]), .ZN(_add_513_n5 ) );
AND2_X4 _add_513_U5  ( .A1(_add_513_n72 ), .A2(_add_513_n73 ), .ZN(_add_513_n4 ) );
AND2_X4 _add_513_U4  ( .A1(H1[23]), .A2(SHA1_result_151), .ZN(_add_513_n3 ));
OR2_X4 _add_513_U3  ( .A1(SHA1_result_129), .A2(H1[1]), .ZN(_add_513_n2 ) );
OR2_X4 _add_513_U2  ( .A1(SHA1_result_134), .A2(H1[6]), .ZN(_add_513_n1 ) );
INV_X4 _add_516_U423  ( .A(H4[8]), .ZN(_add_516_n389 ) );
INV_X4 _add_516_U422  ( .A(SHA1_result[40]), .ZN(_add_516_n390 ) );
NAND2_X2 _add_516_U421  ( .A1(_add_516_n389 ), .A2(_add_516_n390 ), .ZN(_add_516_n260 ) );
INV_X4 _add_516_U420  ( .A(_add_516_n45 ), .ZN(_add_516_n388 ) );
NAND2_X2 _add_516_U419  ( .A1(H4[7]), .A2(SHA1_result[39]), .ZN(_add_516_n47 ) );
NAND2_X2 _add_516_U418  ( .A1(H4[4]), .A2(SHA1_result[36]), .ZN(_add_516_n386 ) );
NAND2_X2 _add_516_U417  ( .A1(H4[5]), .A2(SHA1_result[37]), .ZN(_add_516_n387 ) );
NAND2_X2 _add_516_U416  ( .A1(_add_516_n386 ), .A2(_add_516_n387 ), .ZN(_add_516_n384 ) );
NAND2_X2 _add_516_U415  ( .A1(_add_516_n260 ), .A2(_add_516_n40 ), .ZN(_add_516_n365 ) );
NAND2_X2 _add_516_U414  ( .A1(H4[8]), .A2(SHA1_result[40]), .ZN(_add_516_n304 ) );
INV_X4 _add_516_U413  ( .A(H4[3]), .ZN(_add_516_n381 ) );
INV_X4 _add_516_U412  ( .A(SHA1_result[35]), .ZN(_add_516_n382 ) );
NAND2_X2 _add_516_U411  ( .A1(_add_516_n381 ), .A2(_add_516_n382 ), .ZN(_add_516_n69 ) );
INV_X4 _add_516_U410  ( .A(_add_516_n117 ), .ZN(_add_516_n377 ) );
INV_X4 _add_516_U409  ( .A(_add_516_n69 ), .ZN(_add_516_n294 ) );
NAND2_X2 _add_516_U408  ( .A1(H4[3]), .A2(SHA1_result[35]), .ZN(_add_516_n68 ) );
NAND2_X2 _add_516_U407  ( .A1(H4[0]), .A2(SHA1_result[32]), .ZN(_add_516_n379 ) );
NAND2_X2 _add_516_U406  ( .A1(H4[1]), .A2(SHA1_result[33]), .ZN(_add_516_n380 ) );
NAND2_X2 _add_516_U405  ( .A1(_add_516_n379 ), .A2(_add_516_n380 ), .ZN(_add_516_n376 ) );
INV_X4 _add_516_U404  ( .A(_add_516_n42 ), .ZN(_add_516_n274 ) );
NAND2_X2 _add_516_U403  ( .A1(_add_516_n274 ), .A2(_add_516_n260 ), .ZN(_add_516_n363 ) );
INV_X4 _add_516_U402  ( .A(H4[9]), .ZN(_add_516_n371 ) );
INV_X4 _add_516_U401  ( .A(n14797), .ZN(_add_516_n372 ) );
NAND2_X2 _add_516_U400  ( .A1(_add_516_n371 ), .A2(_add_516_n372 ), .ZN(_add_516_n34 ) );
NAND2_X2 _add_516_U399  ( .A1(_add_516_n31 ), .A2(_add_516_n34 ), .ZN(_add_516_n370 ) );
NAND2_X2 _add_516_U398  ( .A1(H4[9]), .A2(n14797), .ZN(_add_516_n33 ) );
NAND2_X2 _add_516_U397  ( .A1(_add_516_n370 ), .A2(_add_516_n33 ), .ZN(_add_516_n366 ) );
INV_X4 _add_516_U396  ( .A(H4[10]), .ZN(_add_516_n368 ) );
INV_X4 _add_516_U395  ( .A(SHA1_result[42]), .ZN(_add_516_n369 ) );
NAND2_X2 _add_516_U394  ( .A1(_add_516_n368 ), .A2(_add_516_n369 ), .ZN(_add_516_n297 ) );
NAND2_X2 _add_516_U393  ( .A1(H4[10]), .A2(SHA1_result[42]), .ZN(_add_516_n305 ) );
NAND2_X2 _add_516_U392  ( .A1(_add_516_n297 ), .A2(_add_516_n305 ), .ZN(_add_516_n367 ) );
XNOR2_X2 _add_516_U391  ( .A(_add_516_n366 ), .B(_add_516_n367 ), .ZN(N990));
INV_X4 _add_516_U390  ( .A(_add_516_n304 ), .ZN(_add_516_n37 ) );
INV_X4 _add_516_U389  ( .A(_add_516_n365 ), .ZN(_add_516_n364 ) );
NAND2_X2 _add_516_U388  ( .A1(_add_516_n362 ), .A2(_add_516_n18 ), .ZN(_add_516_n361 ) );
NAND2_X2 _add_516_U387  ( .A1(_add_516_n34 ), .A2(_add_516_n361 ), .ZN(_add_516_n360 ) );
NAND2_X2 _add_516_U386  ( .A1(_add_516_n360 ), .A2(_add_516_n33 ), .ZN(_add_516_n359 ) );
NAND2_X2 _add_516_U385  ( .A1(_add_516_n359 ), .A2(_add_516_n297 ), .ZN(_add_516_n358 ) );
NAND2_X2 _add_516_U384  ( .A1(_add_516_n358 ), .A2(_add_516_n305 ), .ZN(_add_516_n354 ) );
NAND2_X2 _add_516_U383  ( .A1(H4[11]), .A2(n14810), .ZN(_add_516_n303 ) );
INV_X4 _add_516_U382  ( .A(H4[11]), .ZN(_add_516_n356 ) );
INV_X4 _add_516_U381  ( .A(n14810), .ZN(_add_516_n357 ) );
NAND2_X2 _add_516_U380  ( .A1(_add_516_n356 ), .A2(_add_516_n357 ), .ZN(_add_516_n272 ) );
NAND2_X2 _add_516_U379  ( .A1(_add_516_n303 ), .A2(_add_516_n272 ), .ZN(_add_516_n355 ) );
XNOR2_X2 _add_516_U378  ( .A(_add_516_n354 ), .B(_add_516_n355 ), .ZN(N991));
INV_X4 _add_516_U377  ( .A(_add_516_n297 ), .ZN(_add_516_n258 ) );
INV_X4 _add_516_U376  ( .A(_add_516_n272 ), .ZN(_add_516_n259 ) );
INV_X4 _add_516_U375  ( .A(_add_516_n260 ), .ZN(_add_516_n38 ) );
INV_X4 _add_516_U374  ( .A(_add_516_n34 ), .ZN(_add_516_n279 ) );
NAND2_X2 _add_516_U373  ( .A1(_add_516_n351 ), .A2(_add_516_n352 ), .ZN(_add_516_n330 ) );
INV_X4 _add_516_U372  ( .A(_add_516_n305 ), .ZN(_add_516_n348 ) );
INV_X4 _add_516_U371  ( .A(_add_516_n303 ), .ZN(_add_516_n349 ) );
NAND2_X2 _add_516_U370  ( .A1(_add_516_n304 ), .A2(_add_516_n33 ), .ZN(_add_516_n347 ) );
NAND2_X2 _add_516_U369  ( .A1(_add_516_n346 ), .A2(_add_516_n347 ), .ZN(_add_516_n345 ) );
NAND2_X2 _add_516_U368  ( .A1(_add_516_n344 ), .A2(_add_516_n345 ), .ZN(_add_516_n343 ) );
NAND2_X2 _add_516_U367  ( .A1(_add_516_n343 ), .A2(_add_516_n272 ), .ZN(_add_516_n331 ) );
INV_X4 _add_516_U366  ( .A(_add_516_n308 ), .ZN(_add_516_n321 ) );
INV_X4 _add_516_U365  ( .A(H4[12]), .ZN(_add_516_n340 ) );
INV_X4 _add_516_U364  ( .A(n14817), .ZN(_add_516_n341 ) );
NAND2_X2 _add_516_U363  ( .A1(_add_516_n340 ), .A2(_add_516_n341 ), .ZN(_add_516_n288 ) );
INV_X4 _add_516_U362  ( .A(_add_516_n288 ), .ZN(_add_516_n276 ) );
XNOR2_X2 _add_516_U361  ( .A(_add_516_n338 ), .B(_add_516_n339 ), .ZN(N992));
NAND2_X2 _add_516_U360  ( .A1(_add_516_n275 ), .A2(_add_516_n337 ), .ZN(_add_516_n336 ) );
INV_X4 _add_516_U359  ( .A(_add_516_n331 ), .ZN(_add_516_n333 ) );
NAND2_X2 _add_516_U358  ( .A1(_add_516_n330 ), .A2(_add_516_n331 ), .ZN(_add_516_n315 ) );
NAND2_X2 _add_516_U357  ( .A1(_add_516_n329 ), .A2(_add_516_n308 ), .ZN(_add_516_n327 ) );
NAND2_X2 _add_516_U356  ( .A1(H4[13]), .A2(SHA1_result[45]), .ZN(_add_516_n319 ) );
NAND2_X2 _add_516_U355  ( .A1(_add_516_n319 ), .A2(_add_516_n277 ), .ZN(_add_516_n328 ) );
XNOR2_X2 _add_516_U354  ( .A(_add_516_n327 ), .B(_add_516_n328 ), .ZN(N993));
NAND2_X2 _add_516_U353  ( .A1(_add_516_n326 ), .A2(_add_516_n308 ), .ZN(_add_516_n325 ) );
NAND2_X2 _add_516_U352  ( .A1(_add_516_n325 ), .A2(_add_516_n277 ), .ZN(_add_516_n324 ) );
NAND2_X2 _add_516_U351  ( .A1(_add_516_n324 ), .A2(_add_516_n319 ), .ZN(_add_516_n322 ) );
NAND2_X2 _add_516_U350  ( .A1(H4[14]), .A2(n14830), .ZN(_add_516_n320 ) );
NAND2_X2 _add_516_U349  ( .A1(_add_516_n264 ), .A2(_add_516_n320 ), .ZN(_add_516_n323 ) );
XNOR2_X2 _add_516_U348  ( .A(_add_516_n322 ), .B(_add_516_n323 ), .ZN(N994));
INV_X4 _add_516_U347  ( .A(_add_516_n320 ), .ZN(_add_516_n317 ) );
NAND4_X2 _add_516_U346  ( .A1(_add_516_n315 ), .A2(_add_516_n2 ), .A3(_add_516_n316 ), .A4(_add_516_n288 ), .ZN(_add_516_n314 ) );
NAND2_X2 _add_516_U345  ( .A1(_add_516_n313 ), .A2(_add_516_n314 ), .ZN(_add_516_n309 ) );
NAND2_X2 _add_516_U344  ( .A1(H4[15]), .A2(SHA1_result[47]), .ZN(_add_516_n261 ) );
INV_X4 _add_516_U343  ( .A(H4[15]), .ZN(_add_516_n311 ) );
INV_X4 _add_516_U342  ( .A(SHA1_result[47]), .ZN(_add_516_n312 ) );
NAND2_X2 _add_516_U341  ( .A1(_add_516_n311 ), .A2(_add_516_n312 ), .ZN(_add_516_n265 ) );
NAND2_X2 _add_516_U340  ( .A1(_add_516_n261 ), .A2(_add_516_n265 ), .ZN(_add_516_n310 ) );
XNOR2_X2 _add_516_U339  ( .A(_add_516_n309 ), .B(_add_516_n310 ), .ZN(N995));
NAND2_X2 _add_516_U338  ( .A1(H4[16]), .A2(SHA1_result[48]), .ZN(_add_516_n242 ) );
NAND2_X2 _add_516_U337  ( .A1(_add_516_n242 ), .A2(_add_516_n236 ), .ZN(_add_516_n244 ) );
INV_X4 _add_516_U336  ( .A(_add_516_n265 ), .ZN(_add_516_n286 ) );
NAND2_X2 _add_516_U335  ( .A1(_add_516_n321 ), .A2(_add_516_n1 ), .ZN(_add_516_n298 ) );
NAND4_X2 _add_516_U334  ( .A1(_add_516_n303 ), .A2(_add_516_n304 ), .A3(_add_516_n305 ), .A4(_add_516_n33 ), .ZN(_add_516_n301 ) );
NAND2_X2 _add_516_U333  ( .A1(_add_516_n258 ), .A2(_add_516_n303 ), .ZN(_add_516_n302 ) );
NAND4_X2 _add_516_U332  ( .A1(_add_516_n300 ), .A2(_add_516_n301 ), .A3(_add_516_n1 ), .A4(_add_516_n302 ), .ZN(_add_516_n299 ) );
NAND2_X2 _add_516_U331  ( .A1(_add_516_n272 ), .A2(_add_516_n297 ), .ZN(_add_516_n296 ) );
NAND2_X2 _add_516_U330  ( .A1(_add_516_n34 ), .A2(_add_516_n260 ), .ZN(_add_516_n295 ) );
NAND2_X2 _add_516_U329  ( .A1(H4[1]), .A2(SHA1_result[33]), .ZN(_add_516_n118 ) );
INV_X4 _add_516_U328  ( .A(_add_516_n118 ), .ZN(_add_516_n215 ) );
NAND4_X2 _add_516_U327  ( .A1(_add_516_n289 ), .A2(_add_516_n290 ), .A3(_add_516_n291 ), .A4(_add_516_n292 ), .ZN(_add_516_n281 ) );
NAND2_X2 _add_516_U326  ( .A1(_add_516_n272 ), .A2(_add_516_n288 ), .ZN(_add_516_n287 ) );
NAND4_X2 _add_516_U325  ( .A1(_add_516_n283 ), .A2(_add_516_n274 ), .A3(_add_516_n284 ), .A4(_add_516_n285 ), .ZN(_add_516_n282 ) );
NAND2_X2 _add_516_U324  ( .A1(_add_516_n281 ), .A2(_add_516_n282 ), .ZN(_add_516_n262 ) );
INV_X4 _add_516_U323  ( .A(_add_516_n280 ), .ZN(_add_516_n277 ) );
NAND4_X2 _add_516_U322  ( .A1(_add_516_n277 ), .A2(_add_516_n264 ), .A3(_add_516_n278 ), .A4(_add_516_n265 ), .ZN(_add_516_n269 ) );
INV_X4 _add_516_U321  ( .A(_add_516_n275 ), .ZN(_add_516_n273 ) );
NAND4_X2 _add_516_U320  ( .A1(_add_516_n271 ), .A2(_add_516_n272 ), .A3(_add_516_n273 ), .A4(_add_516_n274 ), .ZN(_add_516_n270 ) );
NAND2_X2 _add_516_U319  ( .A1(H4[14]), .A2(n14830), .ZN(_add_516_n267 ) );
NAND2_X2 _add_516_U318  ( .A1(H4[13]), .A2(SHA1_result[45]), .ZN(_add_516_n268 ) );
INV_X4 _add_516_U317  ( .A(_add_516_n266 ), .ZN(_add_516_n264 ) );
NAND2_X2 _add_516_U316  ( .A1(_add_516_n264 ), .A2(_add_516_n265 ), .ZN(_add_516_n263 ) );
INV_X4 _add_516_U315  ( .A(_add_516_n261 ), .ZN(_add_516_n247 ) );
NAND2_X2 _add_516_U314  ( .A1(_add_516_n34 ), .A2(_add_516_n260 ), .ZN(_add_516_n257 ) );
INV_X4 _add_516_U313  ( .A(_add_516_n255 ), .ZN(_add_516_n254 ) );
NAND2_X2 _add_516_U312  ( .A1(H4[6]), .A2(SHA1_result[38]), .ZN(_add_516_n251 ) );
NAND2_X2 _add_516_U311  ( .A1(H4[4]), .A2(SHA1_result[36]), .ZN(_add_516_n58 ) );
NAND2_X2 _add_516_U310  ( .A1(H4[5]), .A2(SHA1_result[37]), .ZN(_add_516_n52 ) );
NAND4_X2 _add_516_U309  ( .A1(_add_516_n251 ), .A2(_add_516_n58 ), .A3(_add_516_n52 ), .A4(_add_516_n47 ), .ZN(_add_516_n250 ) );
XNOR2_X2 _add_516_U308  ( .A(_add_516_n244 ), .B(_add_516_n128 ), .ZN(N996));
INV_X4 _add_516_U307  ( .A(_add_516_n225 ), .ZN(_add_516_n236 ) );
NAND2_X2 _add_516_U306  ( .A1(_add_516_n128 ), .A2(_add_516_n236 ), .ZN(_add_516_n243 ) );
NAND2_X2 _add_516_U305  ( .A1(_add_516_n242 ), .A2(_add_516_n243 ), .ZN(_add_516_n239 ) );
NAND2_X2 _add_516_U304  ( .A1(H4[17]), .A2(SHA1_result[49]), .ZN(_add_516_n238 ) );
INV_X4 _add_516_U303  ( .A(_add_516_n223 ), .ZN(_add_516_n241 ) );
NAND2_X2 _add_516_U302  ( .A1(_add_516_n238 ), .A2(_add_516_n241 ), .ZN(_add_516_n240 ) );
XNOR2_X2 _add_516_U301  ( .A(_add_516_n239 ), .B(_add_516_n240 ), .ZN(N997));
NAND2_X2 _add_516_U300  ( .A1(_add_516_n237 ), .A2(_add_516_n238 ), .ZN(_add_516_n229 ) );
INV_X4 _add_516_U299  ( .A(_add_516_n229 ), .ZN(_add_516_n234 ) );
NAND2_X2 _add_516_U298  ( .A1(_add_516_n234 ), .A2(_add_516_n235 ), .ZN(_add_516_n230 ) );
INV_X4 _add_516_U297  ( .A(H4[18]), .ZN(_add_516_n232 ) );
INV_X4 _add_516_U296  ( .A(SHA1_result[50]), .ZN(_add_516_n233 ) );
NAND2_X2 _add_516_U295  ( .A1(_add_516_n232 ), .A2(_add_516_n233 ), .ZN(_add_516_n226 ) );
NAND2_X2 _add_516_U294  ( .A1(H4[18]), .A2(SHA1_result[50]), .ZN(_add_516_n228 ) );
NAND2_X2 _add_516_U293  ( .A1(_add_516_n226 ), .A2(_add_516_n228 ), .ZN(_add_516_n231 ) );
XNOR2_X2 _add_516_U292  ( .A(_add_516_n230 ), .B(_add_516_n231 ), .ZN(N998));
NAND2_X2 _add_516_U291  ( .A1(_add_516_n229 ), .A2(_add_516_n226 ), .ZN(_add_516_n227 ) );
NAND2_X2 _add_516_U290  ( .A1(_add_516_n227 ), .A2(_add_516_n228 ), .ZN(_add_516_n177 ) );
INV_X4 _add_516_U289  ( .A(_add_516_n177 ), .ZN(_add_516_n221 ) );
INV_X4 _add_516_U288  ( .A(_add_516_n226 ), .ZN(_add_516_n224 ) );
NAND2_X2 _add_516_U287  ( .A1(_add_516_n213 ), .A2(_add_516_n128 ), .ZN(_add_516_n222 ) );
NAND2_X2 _add_516_U286  ( .A1(_add_516_n221 ), .A2(_add_516_n222 ), .ZN(_add_516_n217 ) );
NAND2_X2 _add_516_U285  ( .A1(H4[19]), .A2(SHA1_result[51]), .ZN(_add_516_n126 ) );
INV_X4 _add_516_U284  ( .A(H4[19]), .ZN(_add_516_n219 ) );
INV_X4 _add_516_U283  ( .A(SHA1_result[51]), .ZN(_add_516_n220 ) );
NAND2_X2 _add_516_U282  ( .A1(_add_516_n219 ), .A2(_add_516_n220 ), .ZN(_add_516_n178 ) );
NAND2_X2 _add_516_U281  ( .A1(_add_516_n126 ), .A2(_add_516_n178 ), .ZN(_add_516_n218 ) );
XNOR2_X2 _add_516_U280  ( .A(_add_516_n217 ), .B(_add_516_n218 ), .ZN(N999));
XNOR2_X2 _add_516_U279  ( .A(_add_516_n379 ), .B(_add_516_n214 ), .ZN(N981));
NAND2_X2 _add_516_U278  ( .A1(H4[20]), .A2(SHA1_result[52]), .ZN(_add_516_n208 ) );
NAND2_X2 _add_516_U277  ( .A1(_add_516_n208 ), .A2(_add_516_n210 ), .ZN(_add_516_n211 ) );
NAND2_X2 _add_516_U276  ( .A1(_add_516_n177 ), .A2(_add_516_n178 ), .ZN(_add_516_n125 ) );
NAND2_X2 _add_516_U275  ( .A1(_add_516_n8 ), .A2(_add_516_n128 ), .ZN(_add_516_n212 ) );
XNOR2_X2 _add_516_U274  ( .A(_add_516_n211 ), .B(_add_516_n190 ), .ZN(N1000));
INV_X4 _add_516_U273  ( .A(_add_516_n191 ), .ZN(_add_516_n210 ) );
NAND2_X2 _add_516_U272  ( .A1(_add_516_n190 ), .A2(_add_516_n210 ), .ZN(_add_516_n209 ) );
NAND2_X2 _add_516_U271  ( .A1(_add_516_n208 ), .A2(_add_516_n209 ), .ZN(_add_516_n204 ) );
NAND2_X2 _add_516_U270  ( .A1(H4[21]), .A2(SHA1_result[53]), .ZN(_add_516_n194 ) );
INV_X4 _add_516_U269  ( .A(H4[21]), .ZN(_add_516_n206 ) );
INV_X4 _add_516_U268  ( .A(SHA1_result[53]), .ZN(_add_516_n207 ) );
NAND2_X2 _add_516_U267  ( .A1(_add_516_n206 ), .A2(_add_516_n207 ), .ZN(_add_516_n202 ) );
NAND2_X2 _add_516_U266  ( .A1(_add_516_n194 ), .A2(_add_516_n202 ), .ZN(_add_516_n205 ) );
XNOR2_X2 _add_516_U265  ( .A(_add_516_n204 ), .B(_add_516_n205 ), .ZN(N1001));
INV_X4 _add_516_U264  ( .A(_add_516_n190 ), .ZN(_add_516_n203 ) );
INV_X4 _add_516_U263  ( .A(_add_516_n202 ), .ZN(_add_516_n193 ) );
NAND2_X2 _add_516_U262  ( .A1(_add_516_n196 ), .A2(_add_516_n194 ), .ZN(_add_516_n201 ) );
NAND2_X2 _add_516_U261  ( .A1(H4[22]), .A2(n14681), .ZN(_add_516_n195 ) );
INV_X4 _add_516_U260  ( .A(H4[22]), .ZN(_add_516_n198 ) );
INV_X4 _add_516_U259  ( .A(n14681), .ZN(_add_516_n199 ) );
NAND2_X2 _add_516_U258  ( .A1(_add_516_n198 ), .A2(_add_516_n199 ), .ZN(_add_516_n180 ) );
NAND2_X2 _add_516_U257  ( .A1(_add_516_n195 ), .A2(_add_516_n180 ), .ZN(_add_516_n197 ) );
NAND2_X2 _add_516_U256  ( .A1(_add_516_n182 ), .A2(_add_516_n180 ), .ZN(_add_516_n188 ) );
INV_X4 _add_516_U255  ( .A(_add_516_n180 ), .ZN(_add_516_n192 ) );
NAND2_X2 _add_516_U254  ( .A1(_add_516_n183 ), .A2(_add_516_n190 ), .ZN(_add_516_n189 ) );
NAND2_X2 _add_516_U253  ( .A1(_add_516_n188 ), .A2(_add_516_n189 ), .ZN(_add_516_n184 ) );
INV_X4 _add_516_U252  ( .A(H4[23]), .ZN(_add_516_n186 ) );
INV_X4 _add_516_U251  ( .A(SHA1_result[55]), .ZN(_add_516_n187 ) );
NAND2_X2 _add_516_U250  ( .A1(_add_516_n186 ), .A2(_add_516_n187 ), .ZN(_add_516_n181 ) );
NAND2_X2 _add_516_U249  ( .A1(H4[23]), .A2(SHA1_result[55]), .ZN(_add_516_n130 ) );
NAND2_X2 _add_516_U248  ( .A1(_add_516_n181 ), .A2(_add_516_n130 ), .ZN(_add_516_n185 ) );
XNOR2_X2 _add_516_U247  ( .A(_add_516_n184 ), .B(_add_516_n185 ), .ZN(N1003));
NAND2_X2 _add_516_U246  ( .A1(_add_516_n183 ), .A2(_add_516_n181 ), .ZN(_add_516_n81 ) );
INV_X4 _add_516_U245  ( .A(_add_516_n81 ), .ZN(_add_516_n124 ) );
INV_X4 _add_516_U244  ( .A(_add_516_n26 ), .ZN(_add_516_n179 ) );
NAND2_X2 _add_516_U243  ( .A1(_add_516_n11 ), .A2(_add_516_n29 ), .ZN(_add_516_n176 ) );
NAND2_X2 _add_516_U242  ( .A1(_add_516_n169 ), .A2(_add_516_n175 ), .ZN(_add_516_n141 ) );
NAND2_X2 _add_516_U241  ( .A1(H4[24]), .A2(SHA1_result[56]), .ZN(_add_516_n155 ) );
INV_X4 _add_516_U240  ( .A(H4[24]), .ZN(_add_516_n173 ) );
INV_X4 _add_516_U239  ( .A(SHA1_result[56]), .ZN(_add_516_n174 ) );
NAND2_X2 _add_516_U238  ( .A1(_add_516_n173 ), .A2(_add_516_n174 ), .ZN(_add_516_n157 ) );
NAND2_X2 _add_516_U237  ( .A1(_add_516_n155 ), .A2(_add_516_n157 ), .ZN(_add_516_n172 ) );
XNOR2_X2 _add_516_U236  ( .A(_add_516_n141 ), .B(_add_516_n172 ), .ZN(N1004));
NAND2_X2 _add_516_U235  ( .A1(_add_516_n11 ), .A2(_add_516_n29 ), .ZN(_add_516_n171 ) );
NAND2_X2 _add_516_U234  ( .A1(_add_516_n169 ), .A2(_add_516_n170 ), .ZN(_add_516_n168 ) );
NAND2_X2 _add_516_U233  ( .A1(_add_516_n168 ), .A2(_add_516_n157 ), .ZN(_add_516_n167 ) );
NAND2_X2 _add_516_U232  ( .A1(_add_516_n155 ), .A2(_add_516_n167 ), .ZN(_add_516_n165 ) );
NAND2_X2 _add_516_U231  ( .A1(H4[25]), .A2(SHA1_result[57]), .ZN(_add_516_n156 ) );
NAND2_X2 _add_516_U230  ( .A1(_add_516_n156 ), .A2(_add_516_n30 ), .ZN(_add_516_n166 ) );
XNOR2_X2 _add_516_U229  ( .A(_add_516_n165 ), .B(_add_516_n166 ), .ZN(N1005));
NAND2_X2 _add_516_U228  ( .A1(_add_516_n156 ), .A2(_add_516_n155 ), .ZN(_add_516_n164 ) );
NAND2_X2 _add_516_U227  ( .A1(_add_516_n164 ), .A2(_add_516_n30 ), .ZN(_add_516_n163 ) );
NAND2_X2 _add_516_U226  ( .A1(_add_516_n162 ), .A2(_add_516_n163 ), .ZN(_add_516_n158 ) );
NAND2_X2 _add_516_U225  ( .A1(H4[26]), .A2(SHA1_result[58]), .ZN(_add_516_n154 ) );
INV_X4 _add_516_U224  ( .A(H4[26]), .ZN(_add_516_n160 ) );
INV_X4 _add_516_U223  ( .A(SHA1_result[58]), .ZN(_add_516_n161 ) );
NAND2_X2 _add_516_U222  ( .A1(_add_516_n160 ), .A2(_add_516_n161 ), .ZN(_add_516_n146 ) );
NAND2_X2 _add_516_U221  ( .A1(_add_516_n154 ), .A2(_add_516_n146 ), .ZN(_add_516_n159 ) );
XNOR2_X2 _add_516_U220  ( .A(_add_516_n158 ), .B(_add_516_n159 ), .ZN(N1006));
NAND2_X2 _add_516_U219  ( .A1(_add_516_n9 ), .A2(_add_516_n141 ), .ZN(_add_516_n151 ) );
NAND3_X2 _add_516_U218  ( .A1(_add_516_n154 ), .A2(_add_516_n155 ), .A3(_add_516_n156 ), .ZN(_add_516_n145 ) );
NAND2_X2 _add_516_U217  ( .A1(_add_516_n153 ), .A2(_add_516_n154 ), .ZN(_add_516_n144 ) );
NAND2_X2 _add_516_U216  ( .A1(_add_516_n151 ), .A2(_add_516_n152 ), .ZN(_add_516_n147 ) );
INV_X4 _add_516_U215  ( .A(H4[27]), .ZN(_add_516_n149 ) );
INV_X4 _add_516_U214  ( .A(SHA1_result[59]), .ZN(_add_516_n150 ) );
NAND2_X2 _add_516_U213  ( .A1(_add_516_n149 ), .A2(_add_516_n150 ), .ZN(_add_516_n132 ) );
NAND2_X2 _add_516_U212  ( .A1(H4[27]), .A2(SHA1_result[59]), .ZN(_add_516_n143 ) );
NAND2_X2 _add_516_U211  ( .A1(_add_516_n132 ), .A2(_add_516_n143 ), .ZN(_add_516_n148 ) );
XNOR2_X2 _add_516_U210  ( .A(_add_516_n147 ), .B(_add_516_n148 ), .ZN(N1007));
NAND4_X2 _add_516_U209  ( .A1(_add_516_n144 ), .A2(_add_516_n145 ), .A3(_add_516_n146 ), .A4(_add_516_n132 ), .ZN(_add_516_n142 ) );
NAND2_X2 _add_516_U208  ( .A1(_add_516_n142 ), .A2(_add_516_n143 ), .ZN(_add_516_n133 ) );
INV_X4 _add_516_U207  ( .A(_add_516_n133 ), .ZN(_add_516_n138 ) );
AND2_X2 _add_516_U206  ( .A1(_add_516_n9 ), .A2(_add_516_n132 ), .ZN(_add_516_n140 ) );
NAND2_X2 _add_516_U205  ( .A1(_add_516_n140 ), .A2(_add_516_n141 ), .ZN(_add_516_n139 ) );
NAND2_X2 _add_516_U204  ( .A1(_add_516_n138 ), .A2(_add_516_n139 ), .ZN(_add_516_n134 ) );
INV_X4 _add_516_U203  ( .A(H4[28]), .ZN(_add_516_n136 ) );
INV_X4 _add_516_U202  ( .A(SHA1_result[60]), .ZN(_add_516_n137 ) );
NAND2_X2 _add_516_U201  ( .A1(_add_516_n136 ), .A2(_add_516_n137 ), .ZN(_add_516_n131 ) );
NAND2_X2 _add_516_U200  ( .A1(H4[28]), .A2(SHA1_result[60]), .ZN(_add_516_n89 ) );
NAND2_X2 _add_516_U199  ( .A1(_add_516_n131 ), .A2(_add_516_n89 ), .ZN(_add_516_n135 ) );
XNOR2_X2 _add_516_U198  ( .A(_add_516_n134 ), .B(_add_516_n135 ), .ZN(N1008));
NAND2_X2 _add_516_U197  ( .A1(_add_516_n133 ), .A2(_add_516_n131 ), .ZN(_add_516_n90 ) );
INV_X4 _add_516_U196  ( .A(_add_516_n82 ), .ZN(_add_516_n123 ) );
NAND2_X2 _add_516_U195  ( .A1(_add_516_n26 ), .A2(_add_516_n123 ), .ZN(_add_516_n109 ) );
INV_X4 _add_516_U194  ( .A(_add_516_n130 ), .ZN(_add_516_n129 ) );
NAND2_X2 _add_516_U193  ( .A1(_add_516_n129 ), .A2(_add_516_n123 ), .ZN(_add_516_n93 ) );
NAND4_X2 _add_516_U192  ( .A1(_add_516_n89 ), .A2(_add_516_n90 ), .A3(_add_516_n109 ), .A4(_add_516_n93 ), .ZN(_add_516_n122 ) );
NAND2_X2 _add_516_U191  ( .A1(_add_516_n8 ), .A2(_add_516_n128 ), .ZN(_add_516_n127 ) );
NAND2_X2 _add_516_U190  ( .A1(H4[29]), .A2(SHA1_result[61]), .ZN(_add_516_n92 ) );
INV_X4 _add_516_U189  ( .A(H4[29]), .ZN(_add_516_n120 ) );
INV_X4 _add_516_U188  ( .A(SHA1_result[61]), .ZN(_add_516_n121 ) );
NAND2_X2 _add_516_U187  ( .A1(_add_516_n120 ), .A2(_add_516_n121 ), .ZN(_add_516_n108 ) );
NAND2_X2 _add_516_U186  ( .A1(_add_516_n92 ), .A2(_add_516_n108 ), .ZN(_add_516_n119 ) );
XNOR2_X2 _add_516_U185  ( .A(_add_516_n72 ), .B(_add_516_n116 ), .ZN(N982));
INV_X4 _add_516_U184  ( .A(_add_516_n92 ), .ZN(_add_516_n114 ) );
INV_X4 _add_516_U183  ( .A(_add_516_n108 ), .ZN(_add_516_n95 ) );
INV_X4 _add_516_U182  ( .A(_add_516_n90 ), .ZN(_add_516_n113 ) );
NAND2_X2 _add_516_U181  ( .A1(_add_516_n113 ), .A2(_add_516_n108 ), .ZN(_add_516_n112 ) );
NAND2_X2 _add_516_U180  ( .A1(_add_516_n111 ), .A2(_add_516_n112 ), .ZN(_add_516_n104 ) );
INV_X4 _add_516_U179  ( .A(_add_516_n93 ), .ZN(_add_516_n110 ) );
NAND2_X2 _add_516_U178  ( .A1(_add_516_n110 ), .A2(_add_516_n108 ), .ZN(_add_516_n106 ) );
INV_X4 _add_516_U177  ( .A(_add_516_n109 ), .ZN(_add_516_n83 ) );
NAND2_X2 _add_516_U176  ( .A1(_add_516_n83 ), .A2(_add_516_n108 ), .ZN(_add_516_n107 ) );
NAND2_X2 _add_516_U175  ( .A1(_add_516_n106 ), .A2(_add_516_n107 ), .ZN(_add_516_n105 ) );
NAND2_X2 _add_516_U174  ( .A1(_add_516_n80 ), .A2(_add_516_n103 ), .ZN(_add_516_n102 ) );
NAND2_X2 _add_516_U173  ( .A1(_add_516_n101 ), .A2(_add_516_n102 ), .ZN(_add_516_n97 ) );
NAND2_X2 _add_516_U172  ( .A1(H4[30]), .A2(SHA1_result[62]), .ZN(_add_516_n87 ) );
INV_X4 _add_516_U171  ( .A(H4[30]), .ZN(_add_516_n99 ) );
INV_X4 _add_516_U170  ( .A(SHA1_result[62]), .ZN(_add_516_n100 ) );
NAND2_X2 _add_516_U169  ( .A1(_add_516_n99 ), .A2(_add_516_n100 ), .ZN(_add_516_n96 ) );
NAND2_X2 _add_516_U168  ( .A1(_add_516_n87 ), .A2(_add_516_n96 ), .ZN(_add_516_n98 ) );
XNOR2_X2 _add_516_U167  ( .A(_add_516_n97 ), .B(_add_516_n98 ), .ZN(N1010));
INV_X4 _add_516_U166  ( .A(_add_516_n96 ), .ZN(_add_516_n94 ) );
NAND2_X2 _add_516_U165  ( .A1(_add_516_n92 ), .A2(_add_516_n93 ), .ZN(_add_516_n91 ) );
NAND2_X2 _add_516_U164  ( .A1(_add_516_n79 ), .A2(_add_516_n91 ), .ZN(_add_516_n75 ) );
INV_X4 _add_516_U163  ( .A(_add_516_n79 ), .ZN(_add_516_n88 ) );
INV_X4 _add_516_U162  ( .A(_add_516_n87 ), .ZN(_add_516_n86 ) );
NAND2_X2 _add_516_U161  ( .A1(_add_516_n83 ), .A2(_add_516_n79 ), .ZN(_add_516_n77 ) );
NAND4_X2 _add_516_U160  ( .A1(_add_516_n79 ), .A2(_add_516_n123 ), .A3(_add_516_n124 ), .A4(_add_516_n80 ), .ZN(_add_516_n78 ) );
NAND4_X2 _add_516_U159  ( .A1(_add_516_n75 ), .A2(_add_516_n76 ), .A3(_add_516_n77 ), .A4(_add_516_n78 ), .ZN(_add_516_n73 ) );
XNOR2_X2 _add_516_U158  ( .A(H4[31]), .B(SHA1_result[63]), .ZN(_add_516_n74 ) );
XNOR2_X2 _add_516_U157  ( .A(_add_516_n73 ), .B(_add_516_n74 ), .ZN(N1011));
NAND2_X2 _add_516_U156  ( .A1(_add_516_n68 ), .A2(_add_516_n69 ), .ZN(_add_516_n67 ) );
INV_X4 _add_516_U155  ( .A(_add_516_n58 ), .ZN(_add_516_n65 ) );
XNOR2_X2 _add_516_U154  ( .A(_add_516_n41 ), .B(_add_516_n66 ), .ZN(N984) );
INV_X4 _add_516_U153  ( .A(_add_516_n52 ), .ZN(_add_516_n63 ) );
XNOR2_X2 _add_516_U152  ( .A(_add_516_n61 ), .B(_add_516_n62 ), .ZN(N985) );
NAND2_X2 _add_516_U151  ( .A1(_add_516_n41 ), .A2(_add_516_n58 ), .ZN(_add_516_n57 ) );
NAND2_X2 _add_516_U150  ( .A1(_add_516_n56 ), .A2(_add_516_n57 ), .ZN(_add_516_n53 ) );
NAND2_X2 _add_516_U149  ( .A1(_add_516_n53 ), .A2(_add_516_n52 ), .ZN(_add_516_n54 ) );
NAND2_X2 _add_516_U148  ( .A1(H4[6]), .A2(SHA1_result[38]), .ZN(_add_516_n50 ) );
NAND2_X2 _add_516_U147  ( .A1(_add_516_n50 ), .A2(_add_516_n254 ), .ZN(_add_516_n55 ) );
XNOR2_X2 _add_516_U146  ( .A(_add_516_n54 ), .B(_add_516_n55 ), .ZN(N986) );
NAND2_X2 _add_516_U145  ( .A1(_add_516_n27 ), .A2(_add_516_n50 ), .ZN(_add_516_n49 ) );
INV_X4 _add_516_U144  ( .A(_add_516_n47 ), .ZN(_add_516_n46 ) );
XNOR2_X2 _add_516_U143  ( .A(_add_516_n43 ), .B(_add_516_n44 ), .ZN(N987) );
XNOR2_X2 _add_516_U142  ( .A(_add_516_n35 ), .B(_add_516_n36 ), .ZN(N988) );
NAND2_X2 _add_516_U141  ( .A1(_add_516_n33 ), .A2(_add_516_n34 ), .ZN(_add_516_n32 ) );
XNOR2_X2 _add_516_U140  ( .A(_add_516_n31 ), .B(_add_516_n32 ), .ZN(N989) );
INV_X4 _add_516_U139  ( .A(_add_516_n68 ), .ZN(_add_516_n335 ) );
NAND3_X2 _add_516_U138  ( .A1(SHA1_result[48]), .A2(_add_516_n241 ), .A3(H4[16]), .ZN(_add_516_n237 ) );
NOR2_X2 _add_516_U137  ( .A1(SHA1_result[32]), .A2(H4[0]), .ZN(_add_516_n216 ) );
NOR2_X2 _add_516_U136  ( .A1(_add_516_n4 ), .A2(_add_516_n216 ), .ZN(N980));
NAND3_X2 _add_516_U135  ( .A1(SHA1_result[52]), .A2(H4[20]), .A3(_add_516_n202 ), .ZN(_add_516_n196 ) );
NAND3_X2 _add_516_U134  ( .A1(SHA1_result[34]), .A2(H4[2]), .A3(_add_516_n69 ), .ZN(_add_516_n275 ) );
NOR2_X2 _add_516_U133  ( .A1(H4[25]), .A2(SHA1_result[57]), .ZN(_add_516_n153 ) );
OR2_X2 _add_516_U132  ( .A1(H4[25]), .A2(SHA1_result[57]), .ZN(_add_516_n30 ) );
NOR2_X2 _add_516_U131  ( .A1(SHA1_result[39]), .A2(H4[7]), .ZN(_add_516_n256 ) );
NOR2_X2 _add_516_U130  ( .A1(SHA1_result[38]), .A2(H4[6]), .ZN(_add_516_n255 ) );
NAND3_X2 _add_516_U129  ( .A1(SHA1_result[38]), .A2(H4[6]), .A3(_add_516_n388 ), .ZN(_add_516_n253 ) );
NOR2_X2 _add_516_U128  ( .A1(SHA1_result[48]), .A2(H4[16]), .ZN(_add_516_n225 ) );
NOR2_X2 _add_516_U127  ( .A1(SHA1_result[39]), .A2(H4[7]), .ZN(_add_516_n45 ) );
NOR2_X2 _add_516_U126  ( .A1(SHA1_result[37]), .A2(H4[5]), .ZN(_add_516_n60 ) );
NOR2_X2 _add_516_U125  ( .A1(SHA1_result[33]), .A2(H4[1]), .ZN(_add_516_n117 ) );
NOR2_X2 _add_516_U124  ( .A1(SHA1_result[52]), .A2(H4[20]), .ZN(_add_516_n191 ) );
NOR2_X2 _add_516_U123  ( .A1(SHA1_result[36]), .A2(H4[4]), .ZN(_add_516_n59 ) );
NOR2_X2 _add_516_U122  ( .A1(SHA1_result[34]), .A2(H4[2]), .ZN(_add_516_n71 ) );
NOR2_X2 _add_516_U121  ( .A1(SHA1_result[38]), .A2(H4[6]), .ZN(_add_516_n51 ) );
NOR2_X2 _add_516_U120  ( .A1(SHA1_result[37]), .A2(H4[5]), .ZN(_add_516_n374 ) );
NOR2_X2 _add_516_U119  ( .A1(SHA1_result[38]), .A2(H4[6]), .ZN(_add_516_n375 ) );
OR2_X2 _add_516_U118  ( .A1(_add_516_n81 ), .A2(_add_516_n126 ), .ZN(_add_516_n29 ) );
NAND3_X2 _add_516_U117  ( .A1(_add_516_n288 ), .A2(_add_516_n2 ), .A3(_add_516_n315 ), .ZN(_add_516_n329 ) );
NOR2_X2 _add_516_U116  ( .A1(_add_516_n294 ), .A2(_add_516_n71 ), .ZN(_add_516_n378 ) );
NAND3_X2 _add_516_U115  ( .A1(_add_516_n376 ), .A2(_add_516_n377 ), .A3(_add_516_n378 ), .ZN(_add_516_n337 ) );
NAND3_X2 _add_516_U114  ( .A1(_add_516_n305 ), .A2(_add_516_n279 ), .A3(_add_516_n303 ), .ZN(_add_516_n306 ) );
AND2_X2 _add_516_U113  ( .A1(_add_516_n306 ), .A2(_add_516_n272 ), .ZN(_add_516_n300 ) );
NAND3_X2 _add_516_U112  ( .A1(_add_516_n236 ), .A2(_add_516_n241 ), .A3(_add_516_n128 ), .ZN(_add_516_n235 ) );
NOR2_X2 _add_516_U111  ( .A1(_add_516_n37 ), .A2(_add_516_n364 ), .ZN(_add_516_n362 ) );
NOR2_X2 _add_516_U110  ( .A1(_add_516_n171 ), .A2(_add_516_n10 ), .ZN(_add_516_n170 ) );
NAND3_X2 _add_516_U109  ( .A1(_add_516_n288 ), .A2(_add_516_n2 ), .A3(_add_516_n315 ), .ZN(_add_516_n326 ) );
NAND3_X2 _add_516_U108  ( .A1(_add_516_n365 ), .A2(_add_516_n304 ), .A3(_add_516_n18 ), .ZN(_add_516_n31 ) );
NOR2_X2 _add_516_U107  ( .A1(_add_516_n266 ), .A2(_add_516_n280 ), .ZN(_add_516_n284 ) );
NOR3_X2 _add_516_U106  ( .A1(_add_516_n14 ), .A2(_add_516_n51 ), .A3(_add_516_n45 ), .ZN(_add_516_n291 ) );
NAND3_X2 _add_516_U105  ( .A1(_add_516_n157 ), .A2(_add_516_n30 ), .A3(_add_516_n141 ), .ZN(_add_516_n162 ) );
NAND3_X2 _add_516_U104  ( .A1(_add_516_n3 ), .A2(_add_516_n388 ), .A3(_add_516_n254 ), .ZN(_add_516_n252 ) );
NAND3_X2 _add_516_U103  ( .A1(_add_516_n252 ), .A2(_add_516_n47 ), .A3(_add_516_n253 ), .ZN(_add_516_n249 ) );
OR2_X4 _add_516_U102  ( .A1(_add_516_n117 ), .A2(_add_516_n379 ), .ZN(_add_516_n28 ) );
AND2_X2 _add_516_U101  ( .A1(_add_516_n118 ), .A2(_add_516_n28 ), .ZN(_add_516_n72 ) );
NOR2_X2 _add_516_U100  ( .A1(_add_516_n95 ), .A2(_add_516_n89 ), .ZN(_add_516_n115 ) );
OR2_X2 _add_516_U99  ( .A1(_add_516_n51 ), .A2(_add_516_n52 ), .ZN(_add_516_n27 ) );
NOR2_X2 _add_516_U98  ( .A1(_add_516_n41 ), .A2(_add_516_n59 ), .ZN(_add_516_n64 ) );
AND3_X2 _add_516_U97  ( .A1(_add_516_n180 ), .A2(_add_516_n181 ), .A3(_add_516_n182 ), .ZN(_add_516_n26 ) );
NOR2_X2 _add_516_U96  ( .A1(_add_516_n71 ), .A2(_add_516_n72 ), .ZN(_add_516_n70 ) );
NOR2_X2 _add_516_U95  ( .A1(_add_516_n104 ), .A2(_add_516_n105 ), .ZN(_add_516_n101 ) );
NOR2_X2 _add_516_U94  ( .A1(_add_516_n266 ), .A2(_add_516_n319 ), .ZN(_add_516_n318 ) );
NAND3_X2 _add_516_U93  ( .A1(_add_516_n146 ), .A2(_add_516_n145 ), .A3(_add_516_n144 ), .ZN(_add_516_n152 ) );
NOR2_X2 _add_516_U92  ( .A1(_add_516_n88 ), .A2(_add_516_n90 ), .ZN(_add_516_n84 ) );
NOR2_X2 _add_516_U91  ( .A1(_add_516_n88 ), .A2(_add_516_n89 ), .ZN(_add_516_n85 ) );
NOR3_X2 _add_516_U90  ( .A1(_add_516_n84 ), .A2(_add_516_n85 ), .A3(_add_516_n86 ), .ZN(_add_516_n76 ) );
NOR3_X2 _add_516_U89  ( .A1(_add_516_n15 ), .A2(_add_516_n317 ), .A3(_add_516_n318 ), .ZN(_add_516_n313 ) );
NOR2_X2 _add_516_U88  ( .A1(_add_516_n266 ), .A2(_add_516_n280 ), .ZN(_add_516_n316 ) );
NOR2_X2 _add_516_U87  ( .A1(_add_516_n51 ), .A2(_add_516_n53 ), .ZN(_add_516_n48 ) );
NAND3_X2 _add_516_U86  ( .A1(_add_516_n194 ), .A2(_add_516_n195 ), .A3(_add_516_n196 ), .ZN(_add_516_n182 ) );
NOR2_X2 _add_516_U85  ( .A1(_add_516_n215 ), .A2(_add_516_n4 ), .ZN(_add_516_n293 ) );
NOR3_X2 _add_516_U84  ( .A1(_add_516_n13 ), .A2(_add_516_n293 ), .A3(_add_516_n294 ), .ZN(_add_516_n292 ) );
NOR3_X2 _add_516_U83  ( .A1(_add_516_n287 ), .A2(_add_516_n258 ), .A3(_add_516_n68 ), .ZN(_add_516_n283 ) );
NOR3_X2 _add_516_U82  ( .A1(_add_516_n296 ), .A2(_add_516_n280 ), .A3(_add_516_n276 ), .ZN(_add_516_n289 ) );
NAND3_X2 _add_516_U81  ( .A1(_add_516_n131 ), .A2(_add_516_n132 ), .A3(_add_516_n9 ), .ZN(_add_516_n82 ) );
NOR2_X2 _add_516_U80  ( .A1(_add_516_n114 ), .A2(_add_516_n115 ), .ZN(_add_516_n111 ) );
NOR3_X2 _add_516_U79  ( .A1(_add_516_n295 ), .A2(_add_516_n286 ), .A3(_add_516_n266 ), .ZN(_add_516_n290 ) );
NOR2_X2 _add_516_U78  ( .A1(_add_516_n255 ), .A2(_add_516_n256 ), .ZN(_add_516_n385 ) );
NOR3_X2 _add_516_U77  ( .A1(_add_516_n191 ), .A2(_add_516_n192 ), .A3(_add_516_n193 ), .ZN(_add_516_n183 ) );
NOR3_X2 _add_516_U76  ( .A1(_add_516_n223 ), .A2(_add_516_n224 ), .A3(_add_516_n225 ), .ZN(_add_516_n213 ) );
NOR2_X2 _add_516_U75  ( .A1(_add_516_n12 ), .A2(_add_516_n71 ), .ZN(_add_516_n116 ) );
NOR2_X2 _add_516_U74  ( .A1(_add_516_n48 ), .A2(_add_516_n49 ), .ZN(_add_516_n43 ) );
NOR2_X2 _add_516_U73  ( .A1(_add_516_n45 ), .A2(_add_516_n46 ), .ZN(_add_516_n44 ) );
OR2_X4 _add_516_U72  ( .A1(_add_516_n70 ), .A2(_add_516_n12 ), .ZN(_add_516_n25 ) );
XNOR2_X2 _add_516_U71  ( .A(_add_516_n25 ), .B(_add_516_n67 ), .ZN(N983) );
NOR2_X2 _add_516_U70  ( .A1(_add_516_n64 ), .A2(_add_516_n65 ), .ZN(_add_516_n61 ) );
NOR2_X2 _add_516_U69  ( .A1(_add_516_n63 ), .A2(_add_516_n60 ), .ZN(_add_516_n62 ) );
NOR2_X2 _add_516_U68  ( .A1(_add_516_n215 ), .A2(_add_516_n117 ), .ZN(_add_516_n214 ) );
NOR2_X2 _add_516_U67  ( .A1(_add_516_n59 ), .A2(_add_516_n65 ), .ZN(_add_516_n66 ) );
NAND3_X2 _add_516_U66  ( .A1(_add_516_n3 ), .A2(_add_516_n384 ), .A3(_add_516_n385 ), .ZN(_add_516_n383 ) );
NAND3_X2 _add_516_U65  ( .A1(_add_516_n253 ), .A2(_add_516_n47 ), .A3(_add_516_n383 ), .ZN(_add_516_n40 ) );
NOR2_X2 _add_516_U64  ( .A1(_add_516_n59 ), .A2(_add_516_n60 ), .ZN(_add_516_n56 ) );
NOR2_X2 _add_516_U63  ( .A1(_add_516_n348 ), .A2(_add_516_n349 ), .ZN(_add_516_n344 ) );
NOR2_X2 _add_516_U62  ( .A1(_add_516_n94 ), .A2(_add_516_n95 ), .ZN(_add_516_n79 ) );
AND2_X4 _add_516_U61  ( .A1(_add_516_n68 ), .A2(_add_516_n337 ), .ZN(_add_516_n24 ) );
AND2_X2 _add_516_U60  ( .A1(_add_516_n275 ), .A2(_add_516_n24 ), .ZN(_add_516_n41 ) );
OR2_X4 _add_516_U59  ( .A1(_add_516_n16 ), .A2(_add_516_n263 ), .ZN(_add_516_n23 ) );
OR2_X4 _add_516_U58  ( .A1(_add_516_n269 ), .A2(_add_516_n270 ), .ZN(_add_516_n22 ) );
NAND2_X2 _add_516_U57  ( .A1(_add_516_n22 ), .A2(_add_516_n23 ), .ZN(_add_516_n21 ) );
OR2_X4 _add_516_U56  ( .A1(_add_516_n122 ), .A2(_add_516_n17 ), .ZN(_add_516_n20 ) );
XNOR2_X2 _add_516_U55  ( .A(_add_516_n20 ), .B(_add_516_n119 ), .ZN(N1009));
NOR2_X2 _add_516_U54  ( .A1(_add_516_n374 ), .A2(_add_516_n375 ), .ZN(_add_516_n373 ) );
NAND3_X2 _add_516_U53  ( .A1(_add_516_n5 ), .A2(_add_516_n388 ), .A3(_add_516_n373 ), .ZN(_add_516_n42 ) );
NOR3_X2 _add_516_U52  ( .A1(_add_516_n203 ), .A2(_add_516_n193 ), .A3(_add_516_n191 ), .ZN(_add_516_n200 ) );
OR2_X4 _add_516_U51  ( .A1(_add_516_n200 ), .A2(_add_516_n201 ), .ZN(_add_516_n19 ) );
XNOR2_X2 _add_516_U50  ( .A(_add_516_n19 ), .B(_add_516_n197 ), .ZN(N1002));
NAND3_X2 _add_516_U49  ( .A1(_add_516_n126 ), .A2(_add_516_n125 ), .A3(_add_516_n212 ), .ZN(_add_516_n190 ) );
NAND3_X2 _add_516_U48  ( .A1(_add_516_n125 ), .A2(_add_516_n126 ), .A3(_add_516_n127 ), .ZN(_add_516_n80 ) );
NOR2_X2 _add_516_U47  ( .A1(_add_516_n286 ), .A2(_add_516_n266 ), .ZN(_add_516_n307 ) );
NOR3_X2 _add_516_U46  ( .A1(_add_516_n257 ), .A2(_add_516_n258 ), .A3(_add_516_n259 ), .ZN(_add_516_n248 ) );
NOR2_X2 _add_516_U45  ( .A1(_add_516_n279 ), .A2(_add_516_n38 ), .ZN(_add_516_n278 ) );
NOR2_X2 _add_516_U44  ( .A1(_add_516_n258 ), .A2(_add_516_n276 ), .ZN(_add_516_n271 ) );
NOR2_X2 _add_516_U43  ( .A1(_add_516_n258 ), .A2(_add_516_n279 ), .ZN(_add_516_n346 ) );
NOR2_X2 _add_516_U42  ( .A1(_add_516_n342 ), .A2(_add_516_n333 ), .ZN(_add_516_n338 ) );
NOR2_X2 _add_516_U41  ( .A1(_add_516_n321 ), .A2(_add_516_n276 ), .ZN(_add_516_n339 ) );
NAND3_X2 _add_516_U40  ( .A1(_add_516_n8 ), .A2(_add_516_n124 ), .A3(_add_516_n128 ), .ZN(_add_516_n169 ) );
NOR3_X2 _add_516_U39  ( .A1(_add_516_n82 ), .A2(_add_516_n95 ), .A3(_add_516_n81 ), .ZN(_add_516_n103 ) );
OR2_X2 _add_516_U38  ( .A1(_add_516_n41 ), .A2(_add_516_n363 ), .ZN(_add_516_n18 ) );
NOR2_X2 _add_516_U37  ( .A1(_add_516_n41 ), .A2(_add_516_n42 ), .ZN(_add_516_n353 ) );
NOR2_X2 _add_516_U36  ( .A1(_add_516_n353 ), .A2(_add_516_n40 ), .ZN(_add_516_n350 ) );
NOR2_X2 _add_516_U35  ( .A1(_add_516_n350 ), .A2(_add_516_n330 ), .ZN(_add_516_n342 ) );
NOR2_X2 _add_516_U34  ( .A1(_add_516_n41 ), .A2(_add_516_n42 ), .ZN(_add_516_n39 ) );
NOR2_X2 _add_516_U33  ( .A1(_add_516_n39 ), .A2(_add_516_n40 ), .ZN(_add_516_n35 ) );
NOR2_X2 _add_516_U32  ( .A1(_add_516_n37 ), .A2(_add_516_n38 ), .ZN(_add_516_n36 ) );
NOR3_X2 _add_516_U31  ( .A1(_add_516_n286 ), .A2(_add_516_n279 ), .A3(_add_516_n38 ), .ZN(_add_516_n285 ) );
NOR2_X2 _add_516_U30  ( .A1(_add_516_n38 ), .A2(_add_516_n279 ), .ZN(_add_516_n352 ) );
NOR2_X2 _add_516_U29  ( .A1(_add_516_n258 ), .A2(_add_516_n259 ), .ZN(_add_516_n351 ) );
NOR2_X2 _add_516_U28  ( .A1(_add_516_n335 ), .A2(_add_516_n336 ), .ZN(_add_516_n334 ) );
NOR2_X2 _add_516_U27  ( .A1(_add_516_n334 ), .A2(_add_516_n42 ), .ZN(_add_516_n332 ) );
NOR2_X2 _add_516_U26  ( .A1(_add_516_n176 ), .A2(_add_516_n10 ), .ZN(_add_516_n175 ) );
AND3_X2 _add_516_U25  ( .A1(_add_516_n123 ), .A2(_add_516_n124 ), .A3(_add_516_n80 ), .ZN(_add_516_n17 ) );
NOR2_X2 _add_516_U24  ( .A1(_add_516_n262 ), .A2(_add_516_n21 ), .ZN(_add_516_n245 ) );
NOR2_X2 _add_516_U23  ( .A1(_add_516_n247 ), .A2(_add_516_n6 ), .ZN(_add_516_n246 ) );
NAND3_X2 _add_516_U22  ( .A1(_add_516_n7 ), .A2(_add_516_n245 ), .A3(_add_516_n246 ), .ZN(_add_516_n128 ) );
AND2_X4 _add_516_U21  ( .A1(_add_516_n267 ), .A2(_add_516_n268 ), .ZN(_add_516_n16 ) );
AND2_X4 _add_516_U20  ( .A1(_add_516_n316 ), .A2(_add_516_n321 ), .ZN(_add_516_n15 ) );
OR2_X4 _add_516_U19  ( .A1(_add_516_n59 ), .A2(_add_516_n60 ), .ZN(_add_516_n14 ) );
OR2_X4 _add_516_U18  ( .A1(_add_516_n71 ), .A2(_add_516_n117 ), .ZN(_add_516_n13 ) );
AND2_X4 _add_516_U17  ( .A1(H4[2]), .A2(SHA1_result[34]), .ZN(_add_516_n12 ));
AND2_X4 _add_516_U16  ( .A1(_add_516_n179 ), .A2(_add_516_n130 ), .ZN(_add_516_n11 ) );
AND3_X4 _add_516_U15  ( .A1(_add_516_n177 ), .A2(_add_516_n178 ), .A3(_add_516_n124 ), .ZN(_add_516_n10 ) );
NAND2_X1 _add_516_U14  ( .A1(H4[12]), .A2(n14817), .ZN(_add_516_n308 ) );
AND3_X4 _add_516_U13  ( .A1(_add_516_n157 ), .A2(_add_516_n146 ), .A3(_add_516_n30 ), .ZN(_add_516_n9 ) );
AND2_X4 _add_516_U12  ( .A1(_add_516_n213 ), .A2(_add_516_n178 ), .ZN(_add_516_n8 ) );
AND2_X4 _add_516_U11  ( .A1(_add_516_n298 ), .A2(_add_516_n299 ), .ZN(_add_516_n7 ) );
AND4_X4 _add_516_U10  ( .A1(_add_516_n248 ), .A2(_add_516_n249 ), .A3(_add_516_n250 ), .A4(_add_516_n1 ), .ZN(_add_516_n6 ) );
OR2_X4 _add_516_U9  ( .A1(SHA1_result[36]), .A2(H4[4]), .ZN(_add_516_n5 ) );
AND2_X4 _add_516_U8  ( .A1(H4[0]), .A2(SHA1_result[32]), .ZN(_add_516_n4 ));
OR2_X4 _add_516_U7  ( .A1(SHA1_result[37]), .A2(H4[5]), .ZN(_add_516_n3 ) );
NOR2_X1 _add_516_U6  ( .A1(SHA1_result[49]), .A2(H4[17]), .ZN(_add_516_n223 ) );
NOR2_X1 _add_516_U5  ( .A1(SHA1_result[45]), .A2(H4[13]), .ZN(_add_516_n280 ) );
OR3_X4 _add_516_U4  ( .A1(_add_516_n40 ), .A2(_add_516_n332 ), .A3(_add_516_n333 ), .ZN(_add_516_n2 ) );
NOR2_X1 _add_516_U3  ( .A1(n14830), .A2(H4[14]), .ZN(_add_516_n266 ) );
AND3_X4 _add_516_U2  ( .A1(_add_516_n288 ), .A2(_add_516_n277 ), .A3(_add_516_n307 ), .ZN(_add_516_n1 ) );
NAND2_X2 _add_515_U407  ( .A1(H3[0]), .A2(SHA1_result[64]), .ZN(_add_515_n223 ) );
INV_X4 _add_515_U406  ( .A(H3[0]), .ZN(_add_515_n374 ) );
INV_X4 _add_515_U405  ( .A(SHA1_result[64]), .ZN(_add_515_n375 ) );
NAND2_X2 _add_515_U404  ( .A1(_add_515_n374 ), .A2(_add_515_n375 ), .ZN(_add_515_n360 ) );
NAND2_X2 _add_515_U403  ( .A1(SHA1_result[70]), .A2(H3[6]), .ZN(_add_515_n373 ) );
NAND2_X2 _add_515_U402  ( .A1(H3[7]), .A2(SHA1_result[71]), .ZN(_add_515_n46 ) );
NAND2_X2 _add_515_U401  ( .A1(H3[4]), .A2(SHA1_result[68]), .ZN(_add_515_n62 ) );
NAND2_X2 _add_515_U400  ( .A1(H3[5]), .A2(SHA1_result[69]), .ZN(_add_515_n53 ) );
NAND2_X2 _add_515_U399  ( .A1(_add_515_n62 ), .A2(_add_515_n53 ), .ZN(_add_515_n369 ) );
NAND2_X2 _add_515_U398  ( .A1(_add_515_n263 ), .A2(_add_515_n369 ), .ZN(_add_515_n368 ) );
INV_X4 _add_515_U397  ( .A(_add_515_n39 ), .ZN(_add_515_n324 ) );
INV_X4 _add_515_U396  ( .A(H3[3]), .ZN(_add_515_n366 ) );
INV_X4 _add_515_U395  ( .A(SHA1_result[67]), .ZN(_add_515_n367 ) );
NAND2_X2 _add_515_U394  ( .A1(_add_515_n366 ), .A2(_add_515_n367 ), .ZN(_add_515_n361 ) );
INV_X4 _add_515_U393  ( .A(_add_515_n361 ), .ZN(_add_515_n65 ) );
INV_X4 _add_515_U392  ( .A(H3[1]), .ZN(_add_515_n364 ) );
INV_X4 _add_515_U391  ( .A(SHA1_result[65]), .ZN(_add_515_n365 ) );
NAND2_X2 _add_515_U390  ( .A1(_add_515_n364 ), .A2(_add_515_n365 ), .ZN(_add_515_n116 ) );
NAND2_X2 _add_515_U389  ( .A1(_add_515_n363 ), .A2(_add_515_n116 ), .ZN(_add_515_n284 ) );
INV_X4 _add_515_U388  ( .A(_add_515_n284 ), .ZN(_add_515_n362 ) );
NAND2_X2 _add_515_U387  ( .A1(H3[1]), .A2(SHA1_result[65]), .ZN(_add_515_n117 ) );
NAND2_X2 _add_515_U386  ( .A1(_add_515_n223 ), .A2(_add_515_n117 ), .ZN(_add_515_n286 ) );
NAND2_X2 _add_515_U385  ( .A1(_add_515_n362 ), .A2(_add_515_n286 ), .ZN(_add_515_n359 ) );
NAND2_X2 _add_515_U384  ( .A1(H3[3]), .A2(SHA1_result[67]), .ZN(_add_515_n292 ) );
INV_X4 _add_515_U383  ( .A(_add_515_n292 ), .ZN(_add_515_n66 ) );
INV_X4 _add_515_U382  ( .A(_add_515_n59 ), .ZN(_add_515_n40 ) );
INV_X4 _add_515_U381  ( .A(_add_515_n45 ), .ZN(_add_515_n354 ) );
INV_X4 _add_515_U380  ( .A(_add_515_n48 ), .ZN(_add_515_n355 ) );
INV_X4 _add_515_U379  ( .A(H3[4]), .ZN(_add_515_n357 ) );
INV_X4 _add_515_U378  ( .A(SHA1_result[68]), .ZN(_add_515_n358 ) );
NAND2_X2 _add_515_U377  ( .A1(_add_515_n357 ), .A2(_add_515_n358 ), .ZN(_add_515_n61 ) );
INV_X4 _add_515_U376  ( .A(_add_515_n61 ), .ZN(_add_515_n58 ) );
NAND2_X2 _add_515_U375  ( .A1(H3[9]), .A2(SHA1_result[73]), .ZN(_add_515_n34 ) );
NAND2_X2 _add_515_U374  ( .A1(_add_515_n13 ), .A2(_add_515_n34 ), .ZN(_add_515_n348 ) );
INV_X4 _add_515_U373  ( .A(H3[10]), .ZN(_add_515_n350 ) );
INV_X4 _add_515_U372  ( .A(SHA1_result[74]), .ZN(_add_515_n351 ) );
NAND2_X2 _add_515_U371  ( .A1(_add_515_n350 ), .A2(_add_515_n351 ), .ZN(_add_515_n258 ) );
NAND2_X2 _add_515_U370  ( .A1(H3[10]), .A2(SHA1_result[74]), .ZN(_add_515_n273 ) );
NAND2_X2 _add_515_U369  ( .A1(_add_515_n258 ), .A2(_add_515_n273 ), .ZN(_add_515_n349 ) );
XNOR2_X2 _add_515_U368  ( .A(_add_515_n348 ), .B(_add_515_n349 ), .ZN(N958));
INV_X4 _add_515_U367  ( .A(_add_515_n258 ), .ZN(_add_515_n280 ) );
NAND2_X2 _add_515_U366  ( .A1(_add_515_n30 ), .A2(_add_515_n34 ), .ZN(_add_515_n347 ) );
NAND2_X2 _add_515_U365  ( .A1(_add_515_n346 ), .A2(_add_515_n347 ), .ZN(_add_515_n345 ) );
NAND2_X2 _add_515_U364  ( .A1(_add_515_n345 ), .A2(_add_515_n273 ), .ZN(_add_515_n343 ) );
NAND2_X2 _add_515_U363  ( .A1(H3[11]), .A2(SHA1_result[75]), .ZN(_add_515_n272 ) );
NAND2_X2 _add_515_U362  ( .A1(_add_515_n272 ), .A2(_add_515_n257 ), .ZN(_add_515_n344 ) );
XNOR2_X2 _add_515_U361  ( .A(_add_515_n343 ), .B(_add_515_n344 ), .ZN(N959));
INV_X4 _add_515_U360  ( .A(_add_515_n33 ), .ZN(_add_515_n274 ) );
INV_X4 _add_515_U359  ( .A(_add_515_n37 ), .ZN(_add_515_n259 ) );
INV_X4 _add_515_U358  ( .A(_add_515_n257 ), .ZN(_add_515_n279 ) );
INV_X4 _add_515_U357  ( .A(_add_515_n273 ), .ZN(_add_515_n338 ) );
INV_X4 _add_515_U356  ( .A(_add_515_n272 ), .ZN(_add_515_n339 ) );
NAND2_X2 _add_515_U355  ( .A1(H3[8]), .A2(SHA1_result[72]), .ZN(_add_515_n277 ) );
NAND2_X2 _add_515_U354  ( .A1(H3[9]), .A2(SHA1_result[73]), .ZN(_add_515_n278 ) );
NAND2_X2 _add_515_U353  ( .A1(_add_515_n277 ), .A2(_add_515_n278 ), .ZN(_add_515_n337 ) );
NAND2_X2 _add_515_U352  ( .A1(_add_515_n336 ), .A2(_add_515_n337 ), .ZN(_add_515_n335 ) );
NAND2_X2 _add_515_U351  ( .A1(_add_515_n334 ), .A2(_add_515_n335 ), .ZN(_add_515_n333 ) );
NAND2_X2 _add_515_U350  ( .A1(_add_515_n333 ), .A2(_add_515_n257 ), .ZN(_add_515_n325 ) );
INV_X4 _add_515_U349  ( .A(_add_515_n325 ), .ZN(_add_515_n332 ) );
NAND2_X2 _add_515_U348  ( .A1(H3[12]), .A2(SHA1_result[76]), .ZN(_add_515_n299 ) );
INV_X4 _add_515_U347  ( .A(_add_515_n299 ), .ZN(_add_515_n312 ) );
INV_X4 _add_515_U346  ( .A(H3[12]), .ZN(_add_515_n329 ) );
INV_X4 _add_515_U345  ( .A(SHA1_result[76]), .ZN(_add_515_n330 ) );
NAND2_X2 _add_515_U344  ( .A1(_add_515_n329 ), .A2(_add_515_n330 ), .ZN(_add_515_n321 ) );
INV_X4 _add_515_U343  ( .A(_add_515_n321 ), .ZN(_add_515_n304 ) );
XNOR2_X2 _add_515_U342  ( .A(_add_515_n327 ), .B(_add_515_n328 ), .ZN(N960));
NAND2_X2 _add_515_U341  ( .A1(_add_515_n326 ), .A2(_add_515_n325 ), .ZN(_add_515_n320 ) );
NAND2_X2 _add_515_U340  ( .A1(_add_515_n324 ), .A2(_add_515_n325 ), .ZN(_add_515_n323 ) );
XNOR2_X2 _add_515_U339  ( .A(_add_515_n318 ), .B(_add_515_n319 ), .ZN(N961));
NAND2_X2 _add_515_U338  ( .A1(H3[14]), .A2(SHA1_result[78]), .ZN(_add_515_n301 ) );
INV_X4 _add_515_U337  ( .A(_add_515_n301 ), .ZN(_add_515_n315 ) );
XNOR2_X2 _add_515_U336  ( .A(_add_515_n313 ), .B(_add_515_n314 ), .ZN(N962));
NAND2_X2 _add_515_U335  ( .A1(_add_515_n1 ), .A2(_add_515_n28 ), .ZN(_add_515_n308 ) );
NAND2_X2 _add_515_U334  ( .A1(_add_515_n311 ), .A2(_add_515_n312 ), .ZN(_add_515_n309 ) );
NAND2_X2 _add_515_U333  ( .A1(_add_515_n27 ), .A2(_add_515_n311 ), .ZN(_add_515_n310 ) );
NAND4_X2 _add_515_U332  ( .A1(_add_515_n308 ), .A2(_add_515_n301 ), .A3(_add_515_n309 ), .A4(_add_515_n310 ), .ZN(_add_515_n306 ) );
NAND2_X2 _add_515_U331  ( .A1(H3[15]), .A2(SHA1_result[79]), .ZN(_add_515_n266 ) );
NAND2_X2 _add_515_U330  ( .A1(_add_515_n29 ), .A2(_add_515_n266 ), .ZN(_add_515_n307 ) );
XNOR2_X2 _add_515_U329  ( .A(_add_515_n306 ), .B(_add_515_n307 ), .ZN(N963));
NAND2_X2 _add_515_U328  ( .A1(H3[16]), .A2(SHA1_result[80]), .ZN(_add_515_n247 ) );
NAND2_X2 _add_515_U327  ( .A1(_add_515_n247 ), .A2(_add_515_n249 ), .ZN(_add_515_n250 ) );
NAND2_X2 _add_515_U326  ( .A1(_add_515_n257 ), .A2(_add_515_n258 ), .ZN(_add_515_n297 ) );
NAND4_X2 _add_515_U325  ( .A1(_add_515_n294 ), .A2(_add_515_n274 ), .A3(_add_515_n290 ), .A4(_add_515_n295 ), .ZN(_add_515_n287 ) );
NAND2_X2 _add_515_U324  ( .A1(_add_515_n257 ), .A2(_add_515_n258 ), .ZN(_add_515_n293 ) );
INV_X4 _add_515_U323  ( .A(_add_515_n265 ), .ZN(_add_515_n290 ) );
NAND4_X2 _add_515_U322  ( .A1(_add_515_n289 ), .A2(_add_515_n274 ), .A3(_add_515_n290 ), .A4(_add_515_n291 ), .ZN(_add_515_n288 ) );
NAND2_X2 _add_515_U321  ( .A1(_add_515_n287 ), .A2(_add_515_n288 ), .ZN(_add_515_n267 ) );
INV_X4 _add_515_U320  ( .A(_add_515_n286 ), .ZN(_add_515_n285 ) );
NAND2_X2 _add_515_U319  ( .A1(_add_515_n277 ), .A2(_add_515_n278 ), .ZN(_add_515_n276 ) );
NAND4_X2 _add_515_U318  ( .A1(_add_515_n274 ), .A2(_add_515_n275 ), .A3(_add_515_n276 ), .A4(_add_515_n290 ), .ZN(_add_515_n269 ) );
NAND2_X2 _add_515_U317  ( .A1(_add_515_n272 ), .A2(_add_515_n273 ), .ZN(_add_515_n271 ) );
NAND2_X2 _add_515_U316  ( .A1(_add_515_n269 ), .A2(_add_515_n270 ), .ZN(_add_515_n268 ) );
INV_X4 _add_515_U315  ( .A(_add_515_n266 ), .ZN(_add_515_n253 ) );
INV_X4 _add_515_U314  ( .A(_add_515_n62 ), .ZN(_add_515_n57 ) );
INV_X4 _add_515_U313  ( .A(_add_515_n53 ), .ZN(_add_515_n55 ) );
INV_X4 _add_515_U312  ( .A(_add_515_n263 ), .ZN(_add_515_n262 ) );
XNOR2_X2 _add_515_U311  ( .A(_add_515_n250 ), .B(_add_515_n125 ), .ZN(N964));
INV_X4 _add_515_U310  ( .A(_add_515_n241 ), .ZN(_add_515_n249 ) );
NAND2_X2 _add_515_U309  ( .A1(_add_515_n125 ), .A2(_add_515_n249 ), .ZN(_add_515_n248 ) );
NAND2_X2 _add_515_U308  ( .A1(_add_515_n247 ), .A2(_add_515_n248 ), .ZN(_add_515_n244 ) );
INV_X4 _add_515_U307  ( .A(_add_515_n240 ), .ZN(_add_515_n246 ) );
NAND2_X2 _add_515_U306  ( .A1(H3[17]), .A2(SHA1_result[81]), .ZN(_add_515_n243 ) );
NAND2_X2 _add_515_U305  ( .A1(_add_515_n246 ), .A2(_add_515_n243 ), .ZN(_add_515_n245 ) );
XNOR2_X2 _add_515_U304  ( .A(_add_515_n244 ), .B(_add_515_n245 ), .ZN(N965));
NAND2_X2 _add_515_U303  ( .A1(_add_515_n242 ), .A2(_add_515_n243 ), .ZN(_add_515_n230 ) );
INV_X4 _add_515_U302  ( .A(_add_515_n230 ), .ZN(_add_515_n238 ) );
NAND2_X2 _add_515_U301  ( .A1(_add_515_n233 ), .A2(_add_515_n125 ), .ZN(_add_515_n239 ) );
NAND2_X2 _add_515_U300  ( .A1(_add_515_n238 ), .A2(_add_515_n239 ), .ZN(_add_515_n234 ) );
NAND2_X2 _add_515_U299  ( .A1(H3[18]), .A2(SHA1_result[82]), .ZN(_add_515_n229 ) );
INV_X4 _add_515_U298  ( .A(H3[18]), .ZN(_add_515_n236 ) );
INV_X4 _add_515_U297  ( .A(SHA1_result[82]), .ZN(_add_515_n237 ) );
NAND2_X2 _add_515_U296  ( .A1(_add_515_n236 ), .A2(_add_515_n237 ), .ZN(_add_515_n231 ) );
NAND2_X2 _add_515_U295  ( .A1(_add_515_n229 ), .A2(_add_515_n231 ), .ZN(_add_515_n235 ) );
XNOR2_X2 _add_515_U294  ( .A(_add_515_n234 ), .B(_add_515_n235 ), .ZN(N966));
INV_X4 _add_515_U293  ( .A(_add_515_n125 ), .ZN(_add_515_n232 ) );
NAND2_X2 _add_515_U292  ( .A1(_add_515_n233 ), .A2(_add_515_n231 ), .ZN(_add_515_n219 ) );
NAND2_X2 _add_515_U291  ( .A1(_add_515_n230 ), .A2(_add_515_n231 ), .ZN(_add_515_n228 ) );
NAND2_X2 _add_515_U290  ( .A1(_add_515_n228 ), .A2(_add_515_n229 ), .ZN(_add_515_n184 ) );
INV_X4 _add_515_U289  ( .A(H3[19]), .ZN(_add_515_n225 ) );
INV_X4 _add_515_U288  ( .A(SHA1_result[83]), .ZN(_add_515_n226 ) );
NAND2_X2 _add_515_U287  ( .A1(_add_515_n225 ), .A2(_add_515_n226 ), .ZN(_add_515_n185 ) );
NAND2_X2 _add_515_U286  ( .A1(H3[19]), .A2(SHA1_result[83]), .ZN(_add_515_n220 ) );
NAND2_X2 _add_515_U285  ( .A1(_add_515_n185 ), .A2(_add_515_n220 ), .ZN(_add_515_n224 ) );
INV_X4 _add_515_U284  ( .A(_add_515_n223 ), .ZN(_add_515_n222 ) );
NAND2_X2 _add_515_U283  ( .A1(_add_515_n117 ), .A2(_add_515_n116 ), .ZN(_add_515_n221 ) );
XNOR2_X2 _add_515_U282  ( .A(_add_515_n222 ), .B(_add_515_n221 ), .ZN(N949));
INV_X4 _add_515_U281  ( .A(_add_515_n220 ), .ZN(_add_515_n126 ) );
INV_X4 _add_515_U280  ( .A(_add_515_n219 ), .ZN(_add_515_n218 ) );
NAND2_X2 _add_515_U279  ( .A1(_add_515_n9 ), .A2(_add_515_n125 ), .ZN(_add_515_n217 ) );
NAND2_X2 _add_515_U278  ( .A1(_add_515_n216 ), .A2(_add_515_n217 ), .ZN(_add_515_n192 ) );
INV_X4 _add_515_U277  ( .A(_add_515_n192 ), .ZN(_add_515_n214 ) );
NAND2_X2 _add_515_U276  ( .A1(H3[20]), .A2(SHA1_result[84]), .ZN(_add_515_n207 ) );
INV_X4 _add_515_U275  ( .A(_add_515_n207 ), .ZN(_add_515_n212 ) );
XNOR2_X2 _add_515_U274  ( .A(_add_515_n214 ), .B(_add_515_n215 ), .ZN(N968));
NAND2_X2 _add_515_U273  ( .A1(H3[21]), .A2(SHA1_result[85]), .ZN(_add_515_n206 ) );
INV_X4 _add_515_U272  ( .A(_add_515_n206 ), .ZN(_add_515_n210 ) );
XNOR2_X2 _add_515_U271  ( .A(_add_515_n208 ), .B(_add_515_n209 ), .ZN(N969));
NAND2_X2 _add_515_U270  ( .A1(_add_515_n206 ), .A2(_add_515_n207 ), .ZN(_add_515_n203 ) );
INV_X4 _add_515_U269  ( .A(_add_515_n205 ), .ZN(_add_515_n204 ) );
NAND2_X2 _add_515_U268  ( .A1(_add_515_n203 ), .A2(_add_515_n204 ), .ZN(_add_515_n194 ) );
NAND2_X2 _add_515_U267  ( .A1(_add_515_n193 ), .A2(_add_515_n192 ), .ZN(_add_515_n200 ) );
NAND2_X2 _add_515_U266  ( .A1(_add_515_n194 ), .A2(_add_515_n200 ), .ZN(_add_515_n196 ) );
INV_X4 _add_515_U265  ( .A(H3[22]), .ZN(_add_515_n198 ) );
INV_X4 _add_515_U264  ( .A(SHA1_result[86]), .ZN(_add_515_n199 ) );
NAND2_X2 _add_515_U263  ( .A1(_add_515_n198 ), .A2(_add_515_n199 ), .ZN(_add_515_n181 ) );
NAND2_X2 _add_515_U262  ( .A1(H3[22]), .A2(SHA1_result[86]), .ZN(_add_515_n195 ) );
NAND2_X2 _add_515_U261  ( .A1(_add_515_n181 ), .A2(_add_515_n195 ), .ZN(_add_515_n197 ) );
XNOR2_X2 _add_515_U260  ( .A(_add_515_n196 ), .B(_add_515_n197 ), .ZN(N970));
NAND2_X2 _add_515_U259  ( .A1(_add_515_n194 ), .A2(_add_515_n195 ), .ZN(_add_515_n183 ) );
NAND2_X2 _add_515_U258  ( .A1(_add_515_n183 ), .A2(_add_515_n181 ), .ZN(_add_515_n190 ) );
NAND2_X2 _add_515_U257  ( .A1(_add_515_n6 ), .A2(_add_515_n192 ), .ZN(_add_515_n191 ) );
NAND2_X2 _add_515_U256  ( .A1(_add_515_n190 ), .A2(_add_515_n191 ), .ZN(_add_515_n186 ) );
INV_X4 _add_515_U255  ( .A(H3[23]), .ZN(_add_515_n188 ) );
INV_X4 _add_515_U254  ( .A(SHA1_result[87]), .ZN(_add_515_n189 ) );
NAND2_X2 _add_515_U253  ( .A1(_add_515_n188 ), .A2(_add_515_n189 ), .ZN(_add_515_n182 ) );
NAND2_X2 _add_515_U252  ( .A1(H3[23]), .A2(SHA1_result[87]), .ZN(_add_515_n133 ) );
NAND2_X2 _add_515_U251  ( .A1(_add_515_n182 ), .A2(_add_515_n133 ), .ZN(_add_515_n187 ) );
XNOR2_X2 _add_515_U250  ( .A(_add_515_n186 ), .B(_add_515_n187 ), .ZN(N971));
NAND2_X2 _add_515_U249  ( .A1(_add_515_n6 ), .A2(_add_515_n182 ), .ZN(_add_515_n98 ) );
INV_X4 _add_515_U248  ( .A(_add_515_n98 ), .ZN(_add_515_n109 ) );
NAND3_X2 _add_515_U247  ( .A1(_add_515_n184 ), .A2(_add_515_n185 ), .A3(_add_515_n109 ), .ZN(_add_515_n147 ) );
NAND2_X2 _add_515_U246  ( .A1(_add_515_n126 ), .A2(_add_515_n109 ), .ZN(_add_515_n146 ) );
NAND2_X2 _add_515_U245  ( .A1(H3[24]), .A2(SHA1_result[88]), .ZN(_add_515_n172 ) );
INV_X4 _add_515_U244  ( .A(_add_515_n172 ), .ZN(_add_515_n177 ) );
INV_X4 _add_515_U243  ( .A(H3[24]), .ZN(_add_515_n179 ) );
INV_X4 _add_515_U242  ( .A(SHA1_result[88]), .ZN(_add_515_n180 ) );
XNOR2_X2 _add_515_U241  ( .A(_add_515_n161 ), .B(_add_515_n178 ), .ZN(N972));
NAND2_X2 _add_515_U240  ( .A1(H3[25]), .A2(SHA1_result[89]), .ZN(_add_515_n171 ) );
INV_X4 _add_515_U239  ( .A(_add_515_n171 ), .ZN(_add_515_n175 ) );
XNOR2_X2 _add_515_U238  ( .A(_add_515_n173 ), .B(_add_515_n174 ), .ZN(N973));
NAND2_X2 _add_515_U237  ( .A1(_add_515_n171 ), .A2(_add_515_n172 ), .ZN(_add_515_n160 ) );
INV_X4 _add_515_U236  ( .A(_add_515_n160 ), .ZN(_add_515_n170 ) );
NAND2_X2 _add_515_U235  ( .A1(H3[26]), .A2(SHA1_result[90]), .ZN(_add_515_n158 ) );
INV_X4 _add_515_U234  ( .A(H3[26]), .ZN(_add_515_n166 ) );
INV_X4 _add_515_U233  ( .A(SHA1_result[90]), .ZN(_add_515_n167 ) );
NAND2_X2 _add_515_U232  ( .A1(_add_515_n166 ), .A2(_add_515_n167 ), .ZN(_add_515_n156 ) );
NAND2_X2 _add_515_U231  ( .A1(_add_515_n158 ), .A2(_add_515_n156 ), .ZN(_add_515_n165 ) );
INV_X4 _add_515_U230  ( .A(_add_515_n156 ), .ZN(_add_515_n164 ) );
INV_X4 _add_515_U229  ( .A(_add_515_n143 ), .ZN(_add_515_n162 ) );
INV_X4 _add_515_U228  ( .A(_add_515_n158 ), .ZN(_add_515_n159 ) );
NAND2_X2 _add_515_U227  ( .A1(_add_515_n157 ), .A2(_add_515_n158 ), .ZN(_add_515_n155 ) );
NAND2_X2 _add_515_U226  ( .A1(_add_515_n155 ), .A2(_add_515_n156 ), .ZN(_add_515_n154 ) );
NAND2_X2 _add_515_U225  ( .A1(H3[27]), .A2(SHA1_result[91]), .ZN(_add_515_n139 ) );
INV_X4 _add_515_U224  ( .A(H3[27]), .ZN(_add_515_n150 ) );
INV_X4 _add_515_U223  ( .A(SHA1_result[91]), .ZN(_add_515_n151 ) );
NAND2_X2 _add_515_U222  ( .A1(_add_515_n150 ), .A2(_add_515_n151 ), .ZN(_add_515_n141 ) );
NAND2_X2 _add_515_U221  ( .A1(_add_515_n139 ), .A2(_add_515_n141 ), .ZN(_add_515_n149 ) );
INV_X4 _add_515_U220  ( .A(_add_515_n148 ), .ZN(_add_515_n144 ) );
NAND4_X2 _add_515_U219  ( .A1(_add_515_n133 ), .A2(_add_515_n146 ), .A3(_add_515_n129 ), .A4(_add_515_n147 ), .ZN(_add_515_n145 ) );
NAND2_X2 _add_515_U218  ( .A1(_add_515_n143 ), .A2(_add_515_n141 ), .ZN(_add_515_n132 ) );
NAND2_X2 _add_515_U217  ( .A1(_add_515_n140 ), .A2(_add_515_n141 ), .ZN(_add_515_n138 ) );
NAND2_X2 _add_515_U216  ( .A1(_add_515_n138 ), .A2(_add_515_n139 ), .ZN(_add_515_n89 ) );
NAND2_X2 _add_515_U215  ( .A1(H3[28]), .A2(SHA1_result[92]), .ZN(_add_515_n84 ) );
INV_X4 _add_515_U214  ( .A(H3[28]), .ZN(_add_515_n135 ) );
INV_X4 _add_515_U213  ( .A(SHA1_result[92]), .ZN(_add_515_n136 ) );
NAND2_X2 _add_515_U212  ( .A1(_add_515_n135 ), .A2(_add_515_n136 ), .ZN(_add_515_n91 ) );
NAND2_X2 _add_515_U211  ( .A1(_add_515_n84 ), .A2(_add_515_n91 ), .ZN(_add_515_n134 ) );
NAND2_X2 _add_515_U210  ( .A1(_add_515_n89 ), .A2(_add_515_n91 ), .ZN(_add_515_n127 ) );
INV_X4 _add_515_U209  ( .A(_add_515_n133 ), .ZN(_add_515_n130 ) );
INV_X4 _add_515_U208  ( .A(_add_515_n132 ), .ZN(_add_515_n131 ) );
NAND2_X2 _add_515_U207  ( .A1(_add_515_n131 ), .A2(_add_515_n91 ), .ZN(_add_515_n97 ) );
INV_X4 _add_515_U206  ( .A(_add_515_n97 ), .ZN(_add_515_n122 ) );
NAND2_X2 _add_515_U205  ( .A1(_add_515_n130 ), .A2(_add_515_n122 ), .ZN(_add_515_n94 ) );
INV_X4 _add_515_U204  ( .A(_add_515_n129 ), .ZN(_add_515_n128 ) );
NAND2_X2 _add_515_U203  ( .A1(_add_515_n128 ), .A2(_add_515_n122 ), .ZN(_add_515_n85 ) );
NAND4_X2 _add_515_U202  ( .A1(_add_515_n127 ), .A2(_add_515_n84 ), .A3(_add_515_n94 ), .A4(_add_515_n85 ), .ZN(_add_515_n121 ) );
NAND2_X2 _add_515_U201  ( .A1(_add_515_n9 ), .A2(_add_515_n125 ), .ZN(_add_515_n124 ) );
NAND2_X2 _add_515_U200  ( .A1(_add_515_n123 ), .A2(_add_515_n124 ), .ZN(_add_515_n95 ) );
NAND2_X2 _add_515_U199  ( .A1(H3[29]), .A2(SHA1_result[93]), .ZN(_add_515_n82 ) );
INV_X4 _add_515_U198  ( .A(H3[29]), .ZN(_add_515_n119 ) );
INV_X4 _add_515_U197  ( .A(SHA1_result[93]), .ZN(_add_515_n120 ) );
NAND2_X2 _add_515_U196  ( .A1(_add_515_n119 ), .A2(_add_515_n120 ), .ZN(_add_515_n110 ) );
NAND2_X2 _add_515_U195  ( .A1(_add_515_n82 ), .A2(_add_515_n110 ), .ZN(_add_515_n118 ) );
INV_X4 _add_515_U194  ( .A(_add_515_n116 ), .ZN(_add_515_n115 ) );
XNOR2_X2 _add_515_U193  ( .A(_add_515_n69 ), .B(_add_515_n114 ), .ZN(N950));
INV_X4 _add_515_U192  ( .A(_add_515_n85 ), .ZN(_add_515_n113 ) );
NAND2_X2 _add_515_U191  ( .A1(_add_515_n113 ), .A2(_add_515_n110 ), .ZN(_add_515_n105 ) );
INV_X4 _add_515_U190  ( .A(_add_515_n110 ), .ZN(_add_515_n99 ) );
INV_X4 _add_515_U189  ( .A(_add_515_n82 ), .ZN(_add_515_n112 ) );
NAND2_X2 _add_515_U188  ( .A1(_add_515_n92 ), .A2(_add_515_n110 ), .ZN(_add_515_n107 ) );
NAND4_X2 _add_515_U187  ( .A1(_add_515_n122 ), .A2(_add_515_n95 ), .A3(_add_515_n109 ), .A4(_add_515_n110 ), .ZN(_add_515_n108 ) );
NAND4_X2 _add_515_U186  ( .A1(_add_515_n105 ), .A2(_add_515_n106 ), .A3(_add_515_n107 ), .A4(_add_515_n108 ), .ZN(_add_515_n101 ) );
NAND2_X2 _add_515_U185  ( .A1(H3[30]), .A2(SHA1_result[94]), .ZN(_add_515_n81 ) );
INV_X4 _add_515_U184  ( .A(H3[30]), .ZN(_add_515_n103 ) );
INV_X4 _add_515_U183  ( .A(SHA1_result[94]), .ZN(_add_515_n104 ) );
NAND2_X2 _add_515_U182  ( .A1(_add_515_n103 ), .A2(_add_515_n104 ), .ZN(_add_515_n100 ) );
NAND2_X2 _add_515_U181  ( .A1(_add_515_n81 ), .A2(_add_515_n100 ), .ZN(_add_515_n102 ) );
XNOR2_X2 _add_515_U180  ( .A(_add_515_n101 ), .B(_add_515_n102 ), .ZN(N978));
INV_X4 _add_515_U179  ( .A(_add_515_n100 ), .ZN(_add_515_n77 ) );
INV_X4 _add_515_U178  ( .A(_add_515_n93 ), .ZN(_add_515_n83 ) );
NAND2_X2 _add_515_U177  ( .A1(_add_515_n95 ), .A2(_add_515_n96 ), .ZN(_add_515_n72 ) );
INV_X4 _add_515_U176  ( .A(_add_515_n94 ), .ZN(_add_515_n92 ) );
NAND2_X2 _add_515_U175  ( .A1(_add_515_n92 ), .A2(_add_515_n93 ), .ZN(_add_515_n86 ) );
INV_X4 _add_515_U174  ( .A(_add_515_n91 ), .ZN(_add_515_n90 ) );
NAND2_X2 _add_515_U173  ( .A1(_add_515_n88 ), .A2(_add_515_n89 ), .ZN(_add_515_n87 ) );
NAND2_X2 _add_515_U172  ( .A1(_add_515_n86 ), .A2(_add_515_n87 ), .ZN(_add_515_n74 ) );
NAND2_X2 _add_515_U171  ( .A1(_add_515_n81 ), .A2(_add_515_n82 ), .ZN(_add_515_n80 ) );
NOR3_X2 _add_515_U170  ( .A1(_add_515_n74 ), .A2(_add_515_n75 ), .A3(_add_515_n76 ), .ZN(_add_515_n73 ) );
NAND2_X2 _add_515_U169  ( .A1(_add_515_n72 ), .A2(_add_515_n73 ), .ZN(_add_515_n70 ) );
XNOR2_X2 _add_515_U168  ( .A(H3[31]), .B(SHA1_result[95]), .ZN(_add_515_n71 ) );
XNOR2_X2 _add_515_U167  ( .A(_add_515_n70 ), .B(_add_515_n71 ), .ZN(N979) );
XNOR2_X2 _add_515_U166  ( .A(_add_515_n63 ), .B(_add_515_n64 ), .ZN(N951) );
NAND2_X2 _add_515_U165  ( .A1(_add_515_n61 ), .A2(_add_515_n62 ), .ZN(_add_515_n60 ) );
XNOR2_X2 _add_515_U164  ( .A(_add_515_n59 ), .B(_add_515_n60 ), .ZN(N952) );
XNOR2_X2 _add_515_U163  ( .A(_add_515_n52 ), .B(_add_515_n54 ), .ZN(N953) );
XNOR2_X2 _add_515_U162  ( .A(_add_515_n49 ), .B(_add_515_n50 ), .ZN(N954) );
INV_X4 _add_515_U161  ( .A(_add_515_n46 ), .ZN(_add_515_n44 ) );
XNOR2_X2 _add_515_U160  ( .A(_add_515_n42 ), .B(_add_515_n43 ), .ZN(N955) );
XNOR2_X2 _add_515_U159  ( .A(_add_515_n35 ), .B(_add_515_n36 ), .ZN(N956) );
INV_X4 _add_515_U158  ( .A(_add_515_n34 ), .ZN(_add_515_n32 ) );
XNOR2_X2 _add_515_U157  ( .A(_add_515_n30 ), .B(_add_515_n31 ), .ZN(N957) );
OR2_X2 _add_515_U156  ( .A1(SHA1_result[79]), .A2(H3[15]), .ZN(_add_515_n29 ) );
NAND3_X2 _add_515_U155  ( .A1(SHA1_result[80]), .A2(_add_515_n246 ), .A3(H3[16]), .ZN(_add_515_n242 ) );
NOR2_X2 _add_515_U154  ( .A1(SHA1_result[84]), .A2(H3[20]), .ZN(_add_515_n202 ) );
NOR2_X2 _add_515_U153  ( .A1(SHA1_result[85]), .A2(H3[21]), .ZN(_add_515_n201 ) );
NOR2_X2 _add_515_U152  ( .A1(_add_515_n201 ), .A2(_add_515_n202 ), .ZN(_add_515_n193 ) );
NAND3_X2 _add_515_U151  ( .A1(SHA1_result[66]), .A2(H3[2]), .A3(_add_515_n361 ), .ZN(_add_515_n296 ) );
NOR2_X2 _add_515_U150  ( .A1(H3[25]), .A2(SHA1_result[89]), .ZN(_add_515_n157 ) );
NOR2_X2 _add_515_U149  ( .A1(SHA1_result[85]), .A2(H3[21]), .ZN(_add_515_n205 ) );
NOR2_X2 _add_515_U148  ( .A1(SHA1_result[81]), .A2(H3[17]), .ZN(_add_515_n240 ) );
NOR2_X2 _add_515_U147  ( .A1(SHA1_result[84]), .A2(H3[20]), .ZN(_add_515_n213 ) );
NOR2_X2 _add_515_U146  ( .A1(SHA1_result[70]), .A2(H3[6]), .ZN(_add_515_n370 ) );
NOR2_X2 _add_515_U145  ( .A1(SHA1_result[71]), .A2(H3[7]), .ZN(_add_515_n372 ) );
NOR2_X2 _add_515_U144  ( .A1(SHA1_result[69]), .A2(H3[5]), .ZN(_add_515_n371 ) );
NOR3_X2 _add_515_U143  ( .A1(_add_515_n370 ), .A2(_add_515_n371 ), .A3(_add_515_n372 ), .ZN(_add_515_n263 ) );
NOR2_X2 _add_515_U142  ( .A1(SHA1_result[80]), .A2(H3[16]), .ZN(_add_515_n241 ) );
NOR2_X2 _add_515_U141  ( .A1(H3[25]), .A2(SHA1_result[89]), .ZN(_add_515_n163 ) );
OR2_X2 _add_515_U140  ( .A1(H3[11]), .A2(SHA1_result[75]), .ZN(_add_515_n257 ) );
NOR2_X2 _add_515_U139  ( .A1(SHA1_result[72]), .A2(H3[8]), .ZN(_add_515_n37 ) );
NOR2_X2 _add_515_U138  ( .A1(SHA1_result[79]), .A2(H3[15]), .ZN(_add_515_n300 ) );
NOR2_X2 _add_515_U137  ( .A1(SHA1_result[71]), .A2(H3[7]), .ZN(_add_515_n45 ) );
NOR2_X2 _add_515_U136  ( .A1(SHA1_result[70]), .A2(H3[6]), .ZN(_add_515_n48 ) );
NOR2_X2 _add_515_U135  ( .A1(SHA1_result[69]), .A2(H3[5]), .ZN(_add_515_n51 ) );
NOR2_X2 _add_515_U134  ( .A1(SHA1_result[66]), .A2(H3[2]), .ZN(_add_515_n68 ) );
NOR2_X2 _add_515_U133  ( .A1(SHA1_result[77]), .A2(H3[13]), .ZN(_add_515_n303 ) );
NOR2_X2 _add_515_U132  ( .A1(SHA1_result[73]), .A2(H3[9]), .ZN(_add_515_n33 ) );
AND3_X2 _add_515_U131  ( .A1(_add_515_n320 ), .A2(_add_515_n321 ), .A3(_add_515_n16 ), .ZN(_add_515_n27 ) );
NAND3_X2 _add_515_U130  ( .A1(_add_515_n29 ), .A2(_add_515_n28 ), .A3(_add_515_n1 ), .ZN(_add_515_n298 ) );
NAND3_X2 _add_515_U129  ( .A1(_add_515_n296 ), .A2(_add_515_n359 ), .A3(_add_515_n292 ), .ZN(_add_515_n59 ) );
NOR2_X2 _add_515_U128  ( .A1(_add_515_n68 ), .A2(_add_515_n69 ), .ZN(_add_515_n67 ) );
NOR2_X2 _add_515_U127  ( .A1(_add_515_n67 ), .A2(_add_515_n11 ), .ZN(_add_515_n63 ) );
NOR2_X2 _add_515_U126  ( .A1(_add_515_n65 ), .A2(_add_515_n66 ), .ZN(_add_515_n64 ) );
NOR2_X2 _add_515_U125  ( .A1(_add_515_n316 ), .A2(_add_515_n1 ), .ZN(_add_515_n313 ) );
NOR2_X2 _add_515_U124  ( .A1(_add_515_n315 ), .A2(_add_515_n305 ), .ZN(_add_515_n314 ) );
NOR2_X2 _add_515_U123  ( .A1(_add_515_n38 ), .A2(_add_515_n39 ), .ZN(_add_515_n35 ) );
NOR2_X2 _add_515_U122  ( .A1(_add_515_n5 ), .A2(_add_515_n37 ), .ZN(_add_515_n36 ) );
NOR2_X2 _add_515_U121  ( .A1(_add_515_n293 ), .A2(_add_515_n37 ), .ZN(_add_515_n289 ) );
NOR2_X2 _add_515_U120  ( .A1(_add_515_n33 ), .A2(_add_515_n280 ), .ZN(_add_515_n346 ) );
NOR2_X2 _add_515_U119  ( .A1(_add_515_n157 ), .A2(_add_515_n170 ), .ZN(_add_515_n169 ) );
NOR2_X2 _add_515_U118  ( .A1(_add_515_n312 ), .A2(_add_515_n27 ), .ZN(_add_515_n317 ) );
NOR2_X2 _add_515_U117  ( .A1(_add_515_n303 ), .A2(_add_515_n317 ), .ZN(_add_515_n316 ) );
NOR2_X2 _add_515_U116  ( .A1(_add_515_n83 ), .A2(_add_515_n84 ), .ZN(_add_515_n79 ) );
NOR2_X2 _add_515_U115  ( .A1(_add_515_n79 ), .A2(_add_515_n80 ), .ZN(_add_515_n78 ) );
NOR2_X2 _add_515_U114  ( .A1(_add_515_n77 ), .A2(_add_515_n78 ), .ZN(_add_515_n76 ) );
NOR2_X2 _add_515_U113  ( .A1(_add_515_n159 ), .A2(_add_515_n160 ), .ZN(_add_515_n153 ) );
NOR2_X2 _add_515_U112  ( .A1(_add_515_n153 ), .A2(_add_515_n154 ), .ZN(_add_515_n140 ) );
NOR2_X2 _add_515_U111  ( .A1(_add_515_n213 ), .A2(_add_515_n214 ), .ZN(_add_515_n211 ) );
NOR2_X2 _add_515_U110  ( .A1(_add_515_n144 ), .A2(_add_515_n145 ), .ZN(_add_515_n142 ) );
NOR2_X2 _add_515_U109  ( .A1(_add_515_n142 ), .A2(_add_515_n132 ), .ZN(_add_515_n137 ) );
NOR2_X2 _add_515_U108  ( .A1(_add_515_n280 ), .A2(_add_515_n33 ), .ZN(_add_515_n336 ) );
OR2_X4 _add_515_U107  ( .A1(_add_515_n51 ), .A2(_add_515_n52 ), .ZN(_add_515_n26 ) );
AND2_X2 _add_515_U106  ( .A1(_add_515_n53 ), .A2(_add_515_n26 ), .ZN(_add_515_n49 ) );
NOR2_X2 _add_515_U105  ( .A1(_add_515_n48 ), .A2(_add_515_n49 ), .ZN(_add_515_n47 ) );
NOR2_X2 _add_515_U104  ( .A1(_add_515_n240 ), .A2(_add_515_n241 ), .ZN(_add_515_n233 ) );
NOR2_X2 _add_515_U103  ( .A1(_add_515_n305 ), .A2(_add_515_n303 ), .ZN(_add_515_n311 ) );
NOR2_X2 _add_515_U102  ( .A1(_add_515_n99 ), .A2(_add_515_n84 ), .ZN(_add_515_n111 ) );
AND3_X2 _add_515_U101  ( .A1(_add_515_n91 ), .A2(_add_515_n110 ), .A3(_add_515_n89 ), .ZN(_add_515_n25 ) );
NOR2_X2 _add_515_U100  ( .A1(_add_515_n57 ), .A2(_add_515_n55 ), .ZN(_add_515_n264 ) );
NAND3_X2 _add_515_U99  ( .A1(_add_515_n264 ), .A2(_add_515_n46 ), .A3(_add_515_n2 ), .ZN(_add_515_n260 ) );
NAND3_X2 _add_515_U98  ( .A1(_add_515_n181 ), .A2(_add_515_n182 ), .A3(_add_515_n183 ), .ZN(_add_515_n129 ) );
OR2_X4 _add_515_U97  ( .A1(_add_515_n115 ), .A2(_add_515_n223 ), .ZN(_add_515_n24 ) );
AND2_X2 _add_515_U96  ( .A1(_add_515_n117 ), .A2(_add_515_n24 ), .ZN(_add_515_n69 ) );
NAND3_X2 _add_515_U95  ( .A1(_add_515_n46 ), .A2(_add_515_n2 ), .A3(_add_515_n262 ), .ZN(_add_515_n261 ) );
NAND3_X2 _add_515_U94  ( .A1(_add_515_n290 ), .A2(_add_515_n260 ), .A3(_add_515_n261 ), .ZN(_add_515_n255 ) );
NAND3_X2 _add_515_U93  ( .A1(_add_515_n257 ), .A2(_add_515_n258 ), .A3(_add_515_n259 ), .ZN(_add_515_n256 ) );
NOR3_X2 _add_515_U92  ( .A1(_add_515_n255 ), .A2(_add_515_n33 ), .A3(_add_515_n256 ), .ZN(_add_515_n254 ) );
NAND3_X2 _add_515_U91  ( .A1(_add_515_n2 ), .A2(_add_515_n46 ), .A3(_add_515_n368 ), .ZN(_add_515_n39 ) );
OR2_X4 _add_515_U90  ( .A1(_add_515_n137 ), .A2(_add_515_n89 ), .ZN(_add_515_n23 ) );
XNOR2_X2 _add_515_U89  ( .A(_add_515_n23 ), .B(_add_515_n134 ), .ZN(N976) );
NOR3_X2 _add_515_U88  ( .A1(_add_515_n25 ), .A2(_add_515_n111 ), .A3(_add_515_n112 ), .ZN(_add_515_n106 ) );
OR2_X4 _add_515_U87  ( .A1(_add_515_n227 ), .A2(_add_515_n184 ), .ZN(_add_515_n22 ) );
XNOR2_X2 _add_515_U86  ( .A(_add_515_n22 ), .B(_add_515_n224 ), .ZN(N967) );
NOR2_X2 _add_515_U85  ( .A1(_add_515_n212 ), .A2(_add_515_n213 ), .ZN(_add_515_n215 ) );
NOR2_X2 _add_515_U84  ( .A1(_add_515_n11 ), .A2(_add_515_n68 ), .ZN(_add_515_n114 ) );
NOR2_X2 _add_515_U83  ( .A1(_add_515_n55 ), .A2(_add_515_n51 ), .ZN(_add_515_n54 ) );
NOR2_X2 _add_515_U82  ( .A1(_add_515_n10 ), .A2(_add_515_n48 ), .ZN(_add_515_n50 ) );
OR2_X4 _add_515_U81  ( .A1(_add_515_n121 ), .A2(_add_515_n17 ), .ZN(_add_515_n21 ) );
XNOR2_X2 _add_515_U80  ( .A(_add_515_n21 ), .B(_add_515_n118 ), .ZN(N977) );
NOR2_X2 _add_515_U79  ( .A1(_add_515_n312 ), .A2(_add_515_n27 ), .ZN(_add_515_n318 ) );
NOR2_X2 _add_515_U78  ( .A1(_add_515_n1 ), .A2(_add_515_n303 ), .ZN(_add_515_n319 ) );
NOR2_X2 _add_515_U77  ( .A1(_add_515_n47 ), .A2(_add_515_n10 ), .ZN(_add_515_n42 ) );
NOR2_X2 _add_515_U76  ( .A1(_add_515_n44 ), .A2(_add_515_n45 ), .ZN(_add_515_n43 ) );
NOR2_X2 _add_515_U75  ( .A1(_add_515_n211 ), .A2(_add_515_n212 ), .ZN(_add_515_n208 ) );
NOR2_X2 _add_515_U74  ( .A1(_add_515_n205 ), .A2(_add_515_n210 ), .ZN(_add_515_n209 ) );
NOR2_X2 _add_515_U73  ( .A1(_add_515_n32 ), .A2(_add_515_n33 ), .ZN(_add_515_n31 ) );
NOR2_X2 _add_515_U72  ( .A1(_add_515_n177 ), .A2(_add_515_n8 ), .ZN(_add_515_n178 ) );
NOR3_X2 _add_515_U71  ( .A1(_add_515_n40 ), .A2(_add_515_n41 ), .A3(_add_515_n37 ), .ZN(_add_515_n353 ) );
NOR2_X2 _add_515_U70  ( .A1(_add_515_n324 ), .A2(_add_515_n37 ), .ZN(_add_515_n352 ) );
NOR3_X2 _add_515_U69  ( .A1(_add_515_n352 ), .A2(_add_515_n353 ), .A3(_add_515_n5 ), .ZN(_add_515_n30 ) );
NOR3_X2 _add_515_U68  ( .A1(_add_515_n163 ), .A2(_add_515_n164 ), .A3(_add_515_n8 ), .ZN(_add_515_n143 ) );
NOR2_X2 _add_515_U67  ( .A1(_add_515_n338 ), .A2(_add_515_n339 ), .ZN(_add_515_n334 ) );
NOR2_X2 _add_515_U66  ( .A1(_add_515_n279 ), .A2(_add_515_n284 ), .ZN(_add_515_n282 ) );
NOR3_X2 _add_515_U65  ( .A1(_add_515_n285 ), .A2(_add_515_n33 ), .A3(_add_515_n280 ), .ZN(_add_515_n281 ) );
OR2_X4 _add_515_U64  ( .A1(_add_515_n152 ), .A2(_add_515_n140 ), .ZN(_add_515_n20 ) );
XNOR2_X2 _add_515_U63  ( .A(_add_515_n20 ), .B(_add_515_n149 ), .ZN(N975) );
OR2_X4 _add_515_U62  ( .A1(_add_515_n168 ), .A2(_add_515_n169 ), .ZN(_add_515_n19 ) );
XNOR2_X2 _add_515_U61  ( .A(_add_515_n19 ), .B(_add_515_n165 ), .ZN(N974) );
NOR2_X2 _add_515_U60  ( .A1(_add_515_n176 ), .A2(_add_515_n177 ), .ZN(_add_515_n173 ) );
NOR2_X2 _add_515_U59  ( .A1(_add_515_n163 ), .A2(_add_515_n175 ), .ZN(_add_515_n174 ) );
NOR2_X2 _add_515_U58  ( .A1(_add_515_n41 ), .A2(_add_515_n296 ), .ZN(_add_515_n295 ) );
NOR2_X2 _add_515_U57  ( .A1(_add_515_n41 ), .A2(_add_515_n292 ), .ZN(_add_515_n291 ) );
NOR2_X2 _add_515_U56  ( .A1(_add_515_n8 ), .A2(_add_515_n161 ), .ZN(_add_515_n176 ) );
NAND3_X2 _add_515_U55  ( .A1(_add_515_n271 ), .A2(_add_515_n257 ), .A3(_add_515_n290 ), .ZN(_add_515_n270 ) );
NOR3_X2 _add_515_U54  ( .A1(_add_515_n161 ), .A2(_add_515_n163 ), .A3(_add_515_n8 ), .ZN(_add_515_n168 ) );
NOR2_X2 _add_515_U53  ( .A1(_add_515_n297 ), .A2(_add_515_n37 ), .ZN(_add_515_n294 ) );
NOR2_X2 _add_515_U52  ( .A1(_add_515_n303 ), .A2(_add_515_n304 ), .ZN(_add_515_n302 ) );
NAND3_X2 _add_515_U51  ( .A1(_add_515_n28 ), .A2(_add_515_n29 ), .A3(_add_515_n302 ), .ZN(_add_515_n265 ) );
NOR2_X2 _add_515_U50  ( .A1(_add_515_n65 ), .A2(_add_515_n68 ), .ZN(_add_515_n363 ) );
NOR2_X2 _add_515_U49  ( .A1(_add_515_n58 ), .A2(_add_515_n51 ), .ZN(_add_515_n356 ) );
NAND3_X2 _add_515_U48  ( .A1(_add_515_n354 ), .A2(_add_515_n355 ), .A3(_add_515_n356 ), .ZN(_add_515_n41 ) );
AND4_X4 _add_515_U47  ( .A1(_add_515_n129 ), .A2(_add_515_n133 ), .A3(_add_515_n146 ), .A4(_add_515_n148 ), .ZN(_add_515_n18 ) );
AND2_X2 _add_515_U46  ( .A1(_add_515_n147 ), .A2(_add_515_n18 ), .ZN(_add_515_n161 ) );
NOR2_X2 _add_515_U45  ( .A1(_add_515_n232 ), .A2(_add_515_n219 ), .ZN(_add_515_n227 ) );
NOR2_X2 _add_515_U44  ( .A1(_add_515_n280 ), .A2(_add_515_n279 ), .ZN(_add_515_n341 ) );
NAND3_X2 _add_515_U43  ( .A1(_add_515_n274 ), .A2(_add_515_n259 ), .A3(_add_515_n341 ), .ZN(_add_515_n326 ) );
NOR2_X2 _add_515_U42  ( .A1(_add_515_n331 ), .A2(_add_515_n332 ), .ZN(_add_515_n327 ) );
NOR2_X2 _add_515_U41  ( .A1(_add_515_n312 ), .A2(_add_515_n304 ), .ZN(_add_515_n328 ) );
NOR3_X2 _add_515_U40  ( .A1(_add_515_n97 ), .A2(_add_515_n83 ), .A3(_add_515_n98 ), .ZN(_add_515_n96 ) );
NOR2_X2 _add_515_U39  ( .A1(_add_515_n126 ), .A2(_add_515_n12 ), .ZN(_add_515_n216 ) );
NOR2_X2 _add_515_U38  ( .A1(_add_515_n40 ), .A2(_add_515_n58 ), .ZN(_add_515_n56 ) );
NOR2_X2 _add_515_U37  ( .A1(_add_515_n56 ), .A2(_add_515_n57 ), .ZN(_add_515_n52 ) );
NOR2_X2 _add_515_U36  ( .A1(_add_515_n90 ), .A2(_add_515_n83 ), .ZN(_add_515_n88 ) );
NOR2_X2 _add_515_U35  ( .A1(_add_515_n40 ), .A2(_add_515_n41 ), .ZN(_add_515_n342 ) );
NOR2_X2 _add_515_U34  ( .A1(_add_515_n342 ), .A2(_add_515_n39 ), .ZN(_add_515_n340 ) );
NOR2_X2 _add_515_U33  ( .A1(_add_515_n340 ), .A2(_add_515_n326 ), .ZN(_add_515_n331 ) );
NOR2_X2 _add_515_U32  ( .A1(_add_515_n40 ), .A2(_add_515_n41 ), .ZN(_add_515_n38 ) );
NOR2_X2 _add_515_U31  ( .A1(_add_515_n40 ), .A2(_add_515_n41 ), .ZN(_add_515_n322 ) );
NOR2_X2 _add_515_U30  ( .A1(_add_515_n77 ), .A2(_add_515_n99 ), .ZN(_add_515_n93 ) );
NOR2_X2 _add_515_U29  ( .A1(_add_515_n126 ), .A2(_add_515_n12 ), .ZN(_add_515_n123 ) );
NOR2_X2 _add_515_U28  ( .A1(_add_515_n279 ), .A2(_add_515_n280 ), .ZN(_add_515_n275 ) );
NAND3_X2 _add_515_U27  ( .A1(_add_515_n9 ), .A2(_add_515_n109 ), .A3(_add_515_n125 ), .ZN(_add_515_n148 ) );
NOR2_X2 _add_515_U26  ( .A1(_add_515_n41 ), .A2(_add_515_n265 ), .ZN(_add_515_n283 ) );
NOR2_X2 _add_515_U25  ( .A1(_add_515_n161 ), .A2(_add_515_n162 ), .ZN(_add_515_n152 ) );
NOR3_X2 _add_515_U24  ( .A1(_add_515_n267 ), .A2(_add_515_n7 ), .A3(_add_515_n268 ), .ZN(_add_515_n251 ) );
NOR2_X2 _add_515_U23  ( .A1(_add_515_n253 ), .A2(_add_515_n254 ), .ZN(_add_515_n252 ) );
NAND3_X2 _add_515_U22  ( .A1(_add_515_n4 ), .A2(_add_515_n251 ), .A3(_add_515_n252 ), .ZN(_add_515_n125 ) );
AND3_X2 _add_515_U21  ( .A1(_add_515_n122 ), .A2(_add_515_n109 ), .A3(_add_515_n95 ), .ZN(_add_515_n17 ) );
NOR2_X2 _add_515_U20  ( .A1(_add_515_n83 ), .A2(_add_515_n85 ), .ZN(_add_515_n75 ) );
OR2_X4 _add_515_U19  ( .A1(_add_515_n322 ), .A2(_add_515_n323 ), .ZN(_add_515_n16 ) );
AND2_X4 _add_515_U18  ( .A1(_add_515_n223 ), .A2(_add_515_n360 ), .ZN(N948));
OR2_X4 _add_515_U17  ( .A1(_add_515_n300 ), .A2(_add_515_n301 ), .ZN(_add_515_n14 ) );
OR2_X4 _add_515_U16  ( .A1(_add_515_n30 ), .A2(_add_515_n33 ), .ZN(_add_515_n13 ) );
AND2_X4 _add_515_U15  ( .A1(_add_515_n184 ), .A2(_add_515_n185 ), .ZN(_add_515_n12 ) );
AND2_X4 _add_515_U14  ( .A1(H3[2]), .A2(SHA1_result[66]), .ZN(_add_515_n11 ));
AND2_X4 _add_515_U13  ( .A1(H3[6]), .A2(SHA1_result[70]), .ZN(_add_515_n10 ));
AND2_X4 _add_515_U12  ( .A1(_add_515_n218 ), .A2(_add_515_n185 ), .ZN(_add_515_n9 ) );
AND2_X4 _add_515_U11  ( .A1(_add_515_n179 ), .A2(_add_515_n180 ), .ZN(_add_515_n8 ) );
AND4_X4 _add_515_U10  ( .A1(_add_515_n281 ), .A2(_add_515_n259 ), .A3(_add_515_n282 ), .A4(_add_515_n283 ), .ZN(_add_515_n7 ) );
OR2_X4 _add_515_U9  ( .A1(SHA1_result[78]), .A2(H3[14]), .ZN(_add_515_n28 ));
NOR2_X1 _add_515_U8  ( .A1(SHA1_result[78]), .A2(H3[14]), .ZN(_add_515_n305 ) );
AND2_X4 _add_515_U7  ( .A1(_add_515_n193 ), .A2(_add_515_n181 ), .ZN(_add_515_n6 ) );
AND2_X4 _add_515_U6  ( .A1(H3[8]), .A2(SHA1_result[72]), .ZN(_add_515_n5 ));
AND3_X4 _add_515_U5  ( .A1(_add_515_n14 ), .A2(_add_515_n298 ), .A3(_add_515_n3 ), .ZN(_add_515_n4 ) );
OR2_X4 _add_515_U4  ( .A1(_add_515_n265 ), .A2(_add_515_n299 ), .ZN(_add_515_n3 ) );
OR2_X4 _add_515_U3  ( .A1(_add_515_n45 ), .A2(_add_515_n373 ), .ZN(_add_515_n2 ) );
AND2_X4 _add_515_U2  ( .A1(H3[13]), .A2(SHA1_result[77]), .ZN(_add_515_n1 ));
INV_X4 _add_1_root_add_136_4_U441  ( .A(_add_1_root_add_136_4_n389 ), .ZN(_add_1_root_add_136_4_n75 ) );
NOR2_X4 _add_1_root_add_136_4_U440  ( .A1(Wt[1]), .A2(N65), .ZN(_add_1_root_add_136_4_n144 ) );
NAND2_X2 _add_1_root_add_136_4_U439  ( .A1(N65), .A2(Wt[1]), .ZN(_add_1_root_add_136_4_n410 ) );
INV_X4 _add_1_root_add_136_4_U438  ( .A(_add_1_root_add_136_4_n409 ), .ZN(_add_1_root_add_136_4_n94 ) );
INV_X4 _add_1_root_add_136_4_U437  ( .A(_add_1_root_add_136_4_n382 ), .ZN(_add_1_root_add_136_4_n398 ) );
INV_X4 _add_1_root_add_136_4_U436  ( .A(_add_1_root_add_136_4_n407 ), .ZN(_add_1_root_add_136_4_n404 ) );
NOR2_X4 _add_1_root_add_136_4_U435  ( .A1(_add_1_root_add_136_4_n103 ), .A2(_add_1_root_add_136_4_n403 ), .ZN(_add_1_root_add_136_4_n392 ) );
INV_X4 _add_1_root_add_136_4_U434  ( .A(_add_1_root_add_136_4_n17 ), .ZN(_add_1_root_add_136_4_n85 ) );
NAND3_X4 _add_1_root_add_136_4_U433  ( .A1(_add_1_root_add_136_4_n42 ), .A2(Wt[5]), .A3(_add_1_root_add_136_4_n66 ), .ZN(_add_1_root_add_136_4_n324 ) );
NOR2_X4 _add_1_root_add_136_4_U432  ( .A1(N70), .A2(Wt[6]), .ZN(_add_1_root_add_136_4_n401 ) );
NAND2_X2 _add_1_root_add_136_4_U431  ( .A1(Wt[4]), .A2(N68), .ZN(_add_1_root_add_136_4_n402 ) );
NAND3_X4 _add_1_root_add_136_4_U430  ( .A1(_add_1_root_add_136_4_n324 ),.A2(_add_1_root_add_136_4_n399 ), .A3(_add_1_root_add_136_4_n12 ),.ZN(_add_1_root_add_136_4_n84 ) );
NAND3_X4 _add_1_root_add_136_4_U429  ( .A1(_add_1_root_add_136_4_n84 ), .A2(_add_1_root_add_136_4_n85 ), .A3(_add_1_root_add_136_4_n398 ), .ZN(_add_1_root_add_136_4_n390 ) );
XNOR2_X2 _add_1_root_add_136_4_U428  ( .A(_add_1_root_add_136_4_n394 ), .B(_add_1_root_add_136_4_n395 ), .ZN(N138) );
NAND4_X2 _add_1_root_add_136_4_U427  ( .A1(_add_1_root_add_136_4_n391 ),.A2(_add_1_root_add_136_4_n389 ), .A3(_add_1_root_add_136_4_n375 ),.A4(_add_1_root_add_136_4_n390 ), .ZN(_add_1_root_add_136_4_n388 ) );
INV_X4 _add_1_root_add_136_4_U426  ( .A(_add_1_root_add_136_4_n372 ), .ZN(_add_1_root_add_136_4_n384 ) );
NAND2_X2 _add_1_root_add_136_4_U425  ( .A1(Wt[12]), .A2(N76), .ZN(_add_1_root_add_136_4_n335 ) );
NAND2_X2 _add_1_root_add_136_4_U424  ( .A1(_add_1_root_add_136_4_n338 ),.A2(_add_1_root_add_136_4_n335 ), .ZN(_add_1_root_add_136_4_n370 ) );
XNOR2_X2 _add_1_root_add_136_4_U423  ( .A(_add_1_root_add_136_4_n369 ), .B(_add_1_root_add_136_4_n370 ), .ZN(N140) );
NAND2_X2 _add_1_root_add_136_4_U422  ( .A1(N77), .A2(Wt[13]), .ZN(_add_1_root_add_136_4_n360 ) );
NOR2_X4 _add_1_root_add_136_4_U421  ( .A1(Wt[13]), .A2(N77), .ZN(_add_1_root_add_136_4_n233 ) );
NAND2_X2 _add_1_root_add_136_4_U420  ( .A1(_add_1_root_add_136_4_n360 ),.A2(_add_1_root_add_136_4_n367 ), .ZN(_add_1_root_add_136_4_n366 ) );
XNOR2_X2 _add_1_root_add_136_4_U419  ( .A(_add_1_root_add_136_4_n365 ), .B(_add_1_root_add_136_4_n366 ), .ZN(N141) );
INV_X4 _add_1_root_add_136_4_U418  ( .A(_add_1_root_add_136_4_n338 ), .ZN(_add_1_root_add_136_4_n363 ) );
INV_X4 _add_1_root_add_136_4_U417  ( .A(_add_1_root_add_136_4_n355 ), .ZN(_add_1_root_add_136_4_n361 ) );
INV_X4 _add_1_root_add_136_4_U416  ( .A(_add_1_root_add_136_4_n360 ), .ZN(_add_1_root_add_136_4_n358 ) );
NOR3_X4 _add_1_root_add_136_4_U415  ( .A1(_add_1_root_add_136_4_n357 ), .A2(_add_1_root_add_136_4_n358 ), .A3(_add_1_root_add_136_4_n359 ), .ZN(_add_1_root_add_136_4_n352 ) );
NAND2_X2 _add_1_root_add_136_4_U414  ( .A1(_add_1_root_add_136_4_n33 ), .A2(_add_1_root_add_136_4_n355 ), .ZN(_add_1_root_add_136_4_n354 ) );
NAND3_X4 _add_1_root_add_136_4_U413  ( .A1(_add_1_root_add_136_4_n352 ),.A2(_add_1_root_add_136_4_n353 ), .A3(_add_1_root_add_136_4_n354 ),.ZN(_add_1_root_add_136_4_n350 ) );
XNOR2_X2 _add_1_root_add_136_4_U412  ( .A(_add_1_root_add_136_4_n350 ), .B(_add_1_root_add_136_4_n351 ), .ZN(N142) );
NAND2_X2 _add_1_root_add_136_4_U411  ( .A1(N79), .A2(Wt[15]), .ZN(_add_1_root_add_136_4_n339 ) );
INV_X4 _add_1_root_add_136_4_U410  ( .A(N79), .ZN(_add_1_root_add_136_4_n344 ) );
INV_X4 _add_1_root_add_136_4_U409  ( .A(Wt[15]), .ZN(_add_1_root_add_136_4_n345 ) );
XNOR2_X2 _add_1_root_add_136_4_U408  ( .A(_add_1_root_add_136_4_n343 ), .B(_add_1_root_add_136_4_n16 ), .ZN(N143) );
NAND3_X4 _add_1_root_add_136_4_U407  ( .A1(N77), .A2(_add_1_root_add_136_4_n341 ), .A3(Wt[13]), .ZN(_add_1_root_add_136_4_n340 ) );
NAND3_X4 _add_1_root_add_136_4_U406  ( .A1(_add_1_root_add_136_4_n340 ),.A2(_add_1_root_add_136_4_n339 ), .A3(_add_1_root_add_136_4_n348 ),.ZN(_add_1_root_add_136_4_n315 ) );
NAND2_X2 _add_1_root_add_136_4_U405  ( .A1(_add_1_root_add_136_4_n315 ),.A2(_add_1_root_add_136_4_n314 ), .ZN(_add_1_root_add_136_4_n317 ) );
NAND2_X2 _add_1_root_add_136_4_U404  ( .A1(_add_1_root_add_136_4_n338 ),.A2(_add_1_root_add_136_4_n59 ), .ZN(_add_1_root_add_136_4_n336 ) );
NAND3_X4 _add_1_root_add_136_4_U403  ( .A1(_add_1_root_add_136_4_n337 ),.A2(_add_1_root_add_136_4_n335 ), .A3(_add_1_root_add_136_4_n336 ),.ZN(_add_1_root_add_136_4_n220 ) );
INV_X4 _add_1_root_add_136_4_U402  ( .A(_add_1_root_add_136_4_n314 ), .ZN(_add_1_root_add_136_4_n232 ) );
INV_X4 _add_1_root_add_136_4_U401  ( .A(_add_1_root_add_136_4_n335 ), .ZN(_add_1_root_add_136_4_n225 ) );
NAND2_X2 _add_1_root_add_136_4_U400  ( .A1(Wt[1]), .A2(N65), .ZN(_add_1_root_add_136_4_n331 ) );
NAND2_X2 _add_1_root_add_136_4_U399  ( .A1(_add_1_root_add_136_4_n327 ),.A2(_add_1_root_add_136_4_n328 ), .ZN(_add_1_root_add_136_4_n326 ) );
NAND2_X2 _add_1_root_add_136_4_U398  ( .A1(_add_1_root_add_136_4_n325 ),.A2(_add_1_root_add_136_4_n326 ), .ZN(_add_1_root_add_136_4_n226 ) );
NAND3_X4 _add_1_root_add_136_4_U397  ( .A1(_add_1_root_add_136_4_n320 ),.A2(_add_1_root_add_136_4_n226 ), .A3(_add_1_root_add_136_4_n319 ),.ZN(_add_1_root_add_136_4_n286 ) );
NAND3_X4 _add_1_root_add_136_4_U396  ( .A1(_add_1_root_add_136_4_n220 ),.A2(_add_1_root_add_136_4_n286 ), .A3(_add_1_root_add_136_4_n318 ),.ZN(_add_1_root_add_136_4_n312 ) );
NAND2_X2 _add_1_root_add_136_4_U395  ( .A1(_add_1_root_add_136_4_n317 ),.A2(_add_1_root_add_136_4_n312 ), .ZN(_add_1_root_add_136_4_n316 ) );
NAND2_X2 _add_1_root_add_136_4_U394  ( .A1(N80), .A2(Wt[16]), .ZN(_add_1_root_add_136_4_n300 ) );
INV_X4 _add_1_root_add_136_4_U393  ( .A(_add_1_root_add_136_4_n300 ), .ZN(_add_1_root_add_136_4_n313 ) );
INV_X4 _add_1_root_add_136_4_U392  ( .A(_add_1_root_add_136_4_n312 ), .ZN(_add_1_root_add_136_4_n310 ) );
INV_X4 _add_1_root_add_136_4_U391  ( .A(N81), .ZN(_add_1_root_add_136_4_n306 ) );
INV_X4 _add_1_root_add_136_4_U390  ( .A(Wt[17]), .ZN(_add_1_root_add_136_4_n307 ) );
NAND2_X2 _add_1_root_add_136_4_U389  ( .A1(_add_1_root_add_136_4_n7 ), .A2(Wt[17]), .ZN(_add_1_root_add_136_4_n242 ) );
XNOR2_X2 _add_1_root_add_136_4_U388  ( .A(_add_1_root_add_136_4_n304 ), .B(_add_1_root_add_136_4_n305 ), .ZN(N145) );
NOR2_X4 _add_1_root_add_136_4_U387  ( .A1(_add_1_root_add_136_4_n303 ), .A2(_add_1_root_add_136_4_n1 ), .ZN(_add_1_root_add_136_4_n234 ) );
NOR2_X4 _add_1_root_add_136_4_U386  ( .A1(N82), .A2(Wt[18]), .ZN(_add_1_root_add_136_4_n275 ) );
XNOR2_X2 _add_1_root_add_136_4_U385  ( .A(_add_1_root_add_136_4_n259 ), .B(_add_1_root_add_136_4_n297 ), .ZN(N146) );
INV_X4 _add_1_root_add_136_4_U384  ( .A(_add_1_root_add_136_4_n272 ), .ZN(_add_1_root_add_136_4_n293 ) );
XNOR2_X2 _add_1_root_add_136_4_U383  ( .A(_add_1_root_add_136_4_n291 ), .B(_add_1_root_add_136_4_n292 ), .ZN(N147) );
NAND2_X2 _add_1_root_add_136_4_U382  ( .A1(N65), .A2(Wt[1]), .ZN(_add_1_root_add_136_4_n143 ) );
XNOR2_X2 _add_1_root_add_136_4_U381  ( .A(_add_1_root_add_136_4_n333 ), .B(_add_1_root_add_136_4_n287 ), .ZN(N129) );
NOR2_X4 _add_1_root_add_136_4_U380  ( .A1(_add_1_root_add_136_4_n279 ), .A2(_add_1_root_add_136_4_n280 ), .ZN(_add_1_root_add_136_4_n276 ) );
INV_X4 _add_1_root_add_136_4_U379  ( .A(N84), .ZN(_add_1_root_add_136_4_n277 ) );
INV_X4 _add_1_root_add_136_4_U378  ( .A(Wt[20]), .ZN(_add_1_root_add_136_4_n278 ) );
NAND2_X2 _add_1_root_add_136_4_U377  ( .A1(N84), .A2(Wt[20]), .ZN(_add_1_root_add_136_4_n258 ) );
XNOR2_X2 _add_1_root_add_136_4_U376  ( .A(_add_1_root_add_136_4_n276 ), .B(_add_1_root_add_136_4_n21 ), .ZN(N148) );
NAND2_X2 _add_1_root_add_136_4_U375  ( .A1(_add_1_root_add_136_4_n271 ),.A2(_add_1_root_add_136_4_n258 ), .ZN(_add_1_root_add_136_4_n270 ) );
INV_X4 _add_1_root_add_136_4_U374  ( .A(Wt[21]), .ZN(_add_1_root_add_136_4_n268 ) );
INV_X4 _add_1_root_add_136_4_U373  ( .A(_add_1_root_add_136_4_n45 ), .ZN(_add_1_root_add_136_4_n247 ) );
XNOR2_X2 _add_1_root_add_136_4_U372  ( .A(_add_1_root_add_136_4_n265 ), .B(_add_1_root_add_136_4_n266 ), .ZN(N149) );
INV_X4 _add_1_root_add_136_4_U371  ( .A(_add_1_root_add_136_4_n258 ), .ZN(_add_1_root_add_136_4_n257 ) );
INV_X4 _add_1_root_add_136_4_U370  ( .A(_add_1_root_add_136_4_n203 ), .ZN(_add_1_root_add_136_4_n215 ) );
INV_X4 _add_1_root_add_136_4_U369  ( .A(N86), .ZN(_add_1_root_add_136_4_n250 ) );
INV_X4 _add_1_root_add_136_4_U368  ( .A(Wt[22]), .ZN(_add_1_root_add_136_4_n251 ) );
XNOR2_X2 _add_1_root_add_136_4_U367  ( .A(_add_1_root_add_136_4_n248 ), .B(_add_1_root_add_136_4_n249 ), .ZN(N150) );
INV_X4 _add_1_root_add_136_4_U366  ( .A(_add_1_root_add_136_4_n245 ), .ZN(_add_1_root_add_136_4_n244 ) );
NOR2_X4 _add_1_root_add_136_4_U365  ( .A1(_add_1_root_add_136_4_n215 ), .A2(_add_1_root_add_136_4_n24 ), .ZN(_add_1_root_add_136_4_n218 ) );
INV_X4 _add_1_root_add_136_4_U364  ( .A(_add_1_root_add_136_4_n205 ), .ZN(_add_1_root_add_136_4_n235 ) );
NOR2_X4 _add_1_root_add_136_4_U363  ( .A1(_add_1_root_add_136_4_n22 ), .A2(_add_1_root_add_136_4_n235 ), .ZN(_add_1_root_add_136_4_n219 ) );
INV_X4 _add_1_root_add_136_4_U362  ( .A(_add_1_root_add_136_4_n234 ), .ZN(_add_1_root_add_136_4_n230 ) );
INV_X4 _add_1_root_add_136_4_U361  ( .A(_add_1_root_add_136_4_n226 ), .ZN(_add_1_root_add_136_4_n224 ) );
NAND3_X4 _add_1_root_add_136_4_U360  ( .A1(_add_1_root_add_136_4_n219 ),.A2(_add_1_root_add_136_4_n218 ), .A3(_add_1_root_add_136_4_n201 ),.ZN(_add_1_root_add_136_4_n138 ) );
NAND2_X2 _add_1_root_add_136_4_U359  ( .A1(N87), .A2(Wt[23]), .ZN(_add_1_root_add_136_4_n209 ) );
INV_X4 _add_1_root_add_136_4_U358  ( .A(_add_1_root_add_136_4_n209 ), .ZN(_add_1_root_add_136_4_n217 ) );
XNOR2_X2 _add_1_root_add_136_4_U357  ( .A(_add_1_root_add_136_4_n130 ), .B(_add_1_root_add_136_4_n216 ), .ZN(N151) );
NAND4_X2 _add_1_root_add_136_4_U356  ( .A1(_add_1_root_add_136_4_n204 ),.A2(_add_1_root_add_136_4_n214 ), .A3(_add_1_root_add_136_4_n37 ),.A4(_add_1_root_add_136_4_n201 ), .ZN(_add_1_root_add_136_4_n211 ) );
INV_X4 _add_1_root_add_136_4_U355  ( .A(_add_1_root_add_136_4_n213 ), .ZN(_add_1_root_add_136_4_n212 ) );
NAND2_X2 _add_1_root_add_136_4_U354  ( .A1(N88), .A2(Wt[24]), .ZN(_add_1_root_add_136_4_n187 ) );
INV_X4 _add_1_root_add_136_4_U353  ( .A(_add_1_root_add_136_4_n187 ), .ZN(_add_1_root_add_136_4_n208 ) );
NAND4_X2 _add_1_root_add_136_4_U352  ( .A1(_add_1_root_add_136_4_n202 ),.A2(_add_1_root_add_136_4_n203 ), .A3(_add_1_root_add_136_4_n204 ),.A4(_add_1_root_add_136_4_n37 ), .ZN(_add_1_root_add_136_4_n199 ) );
INV_X4 _add_1_root_add_136_4_U351  ( .A(_add_1_root_add_136_4_n198 ), .ZN(_add_1_root_add_136_4_n197 ) );
INV_X4 _add_1_root_add_136_4_U350  ( .A(N89), .ZN(_add_1_root_add_136_4_n190 ) );
INV_X4 _add_1_root_add_136_4_U349  ( .A(Wt[25]), .ZN(_add_1_root_add_136_4_n191 ) );
XNOR2_X2 _add_1_root_add_136_4_U348  ( .A(_add_1_root_add_136_4_n188 ), .B(_add_1_root_add_136_4_n189 ), .ZN(N153) );
INV_X4 _add_1_root_add_136_4_U347  ( .A(Wt[26]), .ZN(_add_1_root_add_136_4_n182 ) );
NAND2_X2 _add_1_root_add_136_4_U346  ( .A1(Wt[26]), .A2(N90), .ZN(_add_1_root_add_136_4_n176 ) );
NAND2_X2 _add_1_root_add_136_4_U345  ( .A1(_add_1_root_add_136_4_n177 ),.A2(_add_1_root_add_136_4_n163 ), .ZN(_add_1_root_add_136_4_n167 ) );
NAND2_X2 _add_1_root_add_136_4_U344  ( .A1(_add_1_root_add_136_4_n166 ),.A2(_add_1_root_add_136_4_n138 ), .ZN(_add_1_root_add_136_4_n170 ) );
INV_X4 _add_1_root_add_136_4_U343  ( .A(_add_1_root_add_136_4_n176 ), .ZN(_add_1_root_add_136_4_n175 ) );
NAND2_X2 _add_1_root_add_136_4_U342  ( .A1(_add_1_root_add_136_4_n170 ),.A2(_add_1_root_add_136_4_n171 ), .ZN(_add_1_root_add_136_4_n168 ) );
NAND2_X2 _add_1_root_add_136_4_U341  ( .A1(N91), .A2(Wt[27]), .ZN(_add_1_root_add_136_4_n128 ) );
NAND2_X2 _add_1_root_add_136_4_U340  ( .A1(_add_1_root_add_136_4_n164 ),.A2(_add_1_root_add_136_4_n128 ), .ZN(_add_1_root_add_136_4_n169 ) );
XNOR2_X2 _add_1_root_add_136_4_U339  ( .A(_add_1_root_add_136_4_n168 ), .B(_add_1_root_add_136_4_n169 ), .ZN(N155) );
INV_X4 _add_1_root_add_136_4_U338  ( .A(_add_1_root_add_136_4_n167 ), .ZN(_add_1_root_add_136_4_n166 ) );
NAND2_X2 _add_1_root_add_136_4_U337  ( .A1(_add_1_root_add_136_4_n166 ),.A2(_add_1_root_add_136_4_n164 ), .ZN(_add_1_root_add_136_4_n131 ) );
INV_X4 _add_1_root_add_136_4_U336  ( .A(_add_1_root_add_136_4_n162 ), .ZN(_add_1_root_add_136_4_n125 ) );
INV_X4 _add_1_root_add_136_4_U335  ( .A(N92), .ZN(_add_1_root_add_136_4_n159 ) );
INV_X4 _add_1_root_add_136_4_U334  ( .A(Wt[28]), .ZN(_add_1_root_add_136_4_n160 ) );
NAND2_X2 _add_1_root_add_136_4_U333  ( .A1(_add_1_root_add_136_4_n159 ),.A2(_add_1_root_add_136_4_n160 ), .ZN(_add_1_root_add_136_4_n153 ) );
INV_X4 _add_1_root_add_136_4_U332  ( .A(_add_1_root_add_136_4_n153 ), .ZN(_add_1_root_add_136_4_n139 ) );
NAND2_X2 _add_1_root_add_136_4_U331  ( .A1(N92), .A2(Wt[28]), .ZN(_add_1_root_add_136_4_n141 ) );
INV_X4 _add_1_root_add_136_4_U330  ( .A(_add_1_root_add_136_4_n141 ), .ZN(_add_1_root_add_136_4_n154 ) );
XNOR2_X2 _add_1_root_add_136_4_U329  ( .A(_add_1_root_add_136_4_n157 ), .B(_add_1_root_add_136_4_n158 ), .ZN(N156) );
INV_X4 _add_1_root_add_136_4_U328  ( .A(_add_1_root_add_136_4_n131 ), .ZN(_add_1_root_add_136_4_n137 ) );
NAND2_X2 _add_1_root_add_136_4_U327  ( .A1(_add_1_root_add_136_4_n125 ),.A2(_add_1_root_add_136_4_n153 ), .ZN(_add_1_root_add_136_4_n152 ) );
NAND2_X2 _add_1_root_add_136_4_U326  ( .A1(_add_1_root_add_136_4_n151 ),.A2(_add_1_root_add_136_4_n152 ), .ZN(_add_1_root_add_136_4_n150 ) );
NAND2_X2 _add_1_root_add_136_4_U325  ( .A1(N93), .A2(Wt[29]), .ZN(_add_1_root_add_136_4_n140 ) );
INV_X4 _add_1_root_add_136_4_U324  ( .A(_add_1_root_add_136_4_n140 ), .ZN(_add_1_root_add_136_4_n148 ) );
XNOR2_X2 _add_1_root_add_136_4_U323  ( .A(_add_1_root_add_136_4_n146 ), .B(_add_1_root_add_136_4_n147 ), .ZN(N157) );
NAND2_X2 _add_1_root_add_136_4_U322  ( .A1(N66), .A2(Wt[2]), .ZN(_add_1_root_add_136_4_n110 ) );
NAND2_X2 _add_1_root_add_136_4_U321  ( .A1(_add_1_root_add_136_4_n145 ),.A2(_add_1_root_add_136_4_n110 ), .ZN(_add_1_root_add_136_4_n142 ) );
NAND2_X2 _add_1_root_add_136_4_U320  ( .A1(_add_1_root_add_136_4_n53 ), .A2(_add_1_root_add_136_4_n143 ), .ZN(_add_1_root_add_136_4_n113 ) );
XNOR2_X2 _add_1_root_add_136_4_U319  ( .A(_add_1_root_add_136_4_n142 ), .B(_add_1_root_add_136_4_n113 ), .ZN(N130) );
NAND2_X2 _add_1_root_add_136_4_U318  ( .A1(_add_1_root_add_136_4_n57 ), .A2(_add_1_root_add_136_4_n140 ), .ZN(_add_1_root_add_136_4_n126 ) );
INV_X4 _add_1_root_add_136_4_U317  ( .A(_add_1_root_add_136_4_n126 ), .ZN(_add_1_root_add_136_4_n134 ) );
NAND2_X2 _add_1_root_add_136_4_U316  ( .A1(_add_1_root_add_136_4_n123 ),.A2(_add_1_root_add_136_4_n29 ), .ZN(_add_1_root_add_136_4_n135 ) );
NAND2_X2 _add_1_root_add_136_4_U315  ( .A1(N94), .A2(Wt[30]), .ZN(_add_1_root_add_136_4_n120 ) );
NAND2_X2 _add_1_root_add_136_4_U314  ( .A1(_add_1_root_add_136_4_n124 ),.A2(_add_1_root_add_136_4_n120 ), .ZN(_add_1_root_add_136_4_n133 ) );
XNOR2_X2 _add_1_root_add_136_4_U313  ( .A(_add_1_root_add_136_4_n132 ), .B(_add_1_root_add_136_4_n133 ), .ZN(N158) );
INV_X4 _add_1_root_add_136_4_U312  ( .A(_add_1_root_add_136_4_n128 ), .ZN(_add_1_root_add_136_4_n127 ) );
NAND2_X2 _add_1_root_add_136_4_U311  ( .A1(_add_1_root_add_136_4_n126 ),.A2(_add_1_root_add_136_4_n124 ), .ZN(_add_1_root_add_136_4_n121 ) );
NAND4_X2 _add_1_root_add_136_4_U310  ( .A1(_add_1_root_add_136_4_n119 ),.A2(_add_1_root_add_136_4_n120 ), .A3(_add_1_root_add_136_4_n121 ),.A4(_add_1_root_add_136_4_n122 ), .ZN(_add_1_root_add_136_4_n118 ) );
INV_X4 _add_1_root_add_136_4_U309  ( .A(N95), .ZN(_add_1_root_add_136_4_n116 ) );
XNOR2_X2 _add_1_root_add_136_4_U308  ( .A(_add_1_root_add_136_4_n116 ), .B(Wt[31]), .ZN(_add_1_root_add_136_4_n115 ) );
XNOR2_X2 _add_1_root_add_136_4_U307  ( .A(_add_1_root_add_136_4_n114 ), .B(_add_1_root_add_136_4_n115 ), .ZN(N159) );
INV_X4 _add_1_root_add_136_4_U306  ( .A(_add_1_root_add_136_4_n113 ), .ZN(_add_1_root_add_136_4_n112 ) );
INV_X4 _add_1_root_add_136_4_U305  ( .A(_add_1_root_add_136_4_n110 ), .ZN(_add_1_root_add_136_4_n109 ) );
XNOR2_X2 _add_1_root_add_136_4_U304  ( .A(_add_1_root_add_136_4_n105 ), .B(_add_1_root_add_136_4_n106 ), .ZN(N131) );
NAND2_X2 _add_1_root_add_136_4_U303  ( .A1(N68), .A2(Wt[4]), .ZN(_add_1_root_add_136_4_n96 ) );
INV_X4 _add_1_root_add_136_4_U302  ( .A(_add_1_root_add_136_4_n96 ), .ZN(_add_1_root_add_136_4_n102 ) );
XNOR2_X2 _add_1_root_add_136_4_U301  ( .A(_add_1_root_add_136_4_n103 ), .B(_add_1_root_add_136_4_n104 ), .ZN(N132) );
XNOR2_X2 _add_1_root_add_136_4_U300  ( .A(_add_1_root_add_136_4_n98 ), .B(_add_1_root_add_136_4_n99 ), .ZN(N133) );
NAND2_X2 _add_1_root_add_136_4_U299  ( .A1(_add_1_root_add_136_4_n88 ), .A2(_add_1_root_add_136_4_n14 ), .ZN(_add_1_root_add_136_4_n90 ) );
XNOR2_X2 _add_1_root_add_136_4_U298  ( .A(_add_1_root_add_136_4_n89 ), .B(_add_1_root_add_136_4_n90 ), .ZN(N134) );
XNOR2_X2 _add_1_root_add_136_4_U297  ( .A(_add_1_root_add_136_4_n86 ), .B(_add_1_root_add_136_4_n9 ), .ZN(N135) );
NAND2_X2 _add_1_root_add_136_4_U296  ( .A1(_add_1_root_add_136_4_n85 ), .A2(_add_1_root_add_136_4_n84 ), .ZN(_add_1_root_add_136_4_n81 ) );
NAND2_X2 _add_1_root_add_136_4_U295  ( .A1(_add_1_root_add_136_4_n81 ), .A2(_add_1_root_add_136_4_n82 ), .ZN(_add_1_root_add_136_4_n78 ) );
INV_X4 _add_1_root_add_136_4_U294  ( .A(_add_1_root_add_136_4_n375 ), .ZN(_add_1_root_add_136_4_n80 ) );
XNOR2_X2 _add_1_root_add_136_4_U293  ( .A(_add_1_root_add_136_4_n78 ), .B(_add_1_root_add_136_4_n79 ), .ZN(_add_1_root_add_136_4_n77 ) );
INV_X4 _add_1_root_add_136_4_U292  ( .A(_add_1_root_add_136_4_n77 ), .ZN(N136) );
XNOR2_X2 _add_1_root_add_136_4_U291  ( .A(_add_1_root_add_136_4_n73 ), .B(_add_1_root_add_136_4_n74 ), .ZN(N137) );
NAND2_X4 _add_1_root_add_136_4_U290  ( .A1(_add_1_root_add_136_4_n299 ),.A2(_add_1_root_add_136_4_n300 ), .ZN(_add_1_root_add_136_4_n238 ) );
NAND2_X4 _add_1_root_add_136_4_U289  ( .A1(_add_1_root_add_136_4_n267 ),.A2(_add_1_root_add_136_4_n268 ), .ZN(_add_1_root_add_136_4_n239 ) );
NAND3_X2 _add_1_root_add_136_4_U288  ( .A1(_add_1_root_add_136_4_n11 ), .A2(_add_1_root_add_136_4_n228 ), .A3(_add_1_root_add_136_4_n338 ), .ZN(_add_1_root_add_136_4_n337 ) );
INV_X2 _add_1_root_add_136_4_U287  ( .A(_add_1_root_add_136_4_n233 ), .ZN(_add_1_root_add_136_4_n367 ) );
NOR3_X2 _add_1_root_add_136_4_U286  ( .A1(_add_1_root_add_136_4_n23 ), .A2(_add_1_root_add_136_4_n232 ), .A3(_add_1_root_add_136_4_n25 ), .ZN(_add_1_root_add_136_4_n318 ) );
NAND2_X2 _add_1_root_add_136_4_U285  ( .A1(Wt[14]), .A2(N78), .ZN(_add_1_root_add_136_4_n348 ) );
NAND2_X4 _add_1_root_add_136_4_U284  ( .A1(_add_1_root_add_136_4_n238 ),.A2(_add_1_root_add_136_4_n38 ), .ZN(_add_1_root_add_136_4_n264 ) );
NAND2_X4 _add_1_root_add_136_4_U283  ( .A1(_add_1_root_add_136_4_n306 ),.A2(_add_1_root_add_136_4_n307 ), .ZN(_add_1_root_add_136_4_n237 ) );
NAND2_X1 _add_1_root_add_136_4_U282  ( .A1(_add_1_root_add_136_4_n38 ), .A2(_add_1_root_add_136_4_n242 ), .ZN(_add_1_root_add_136_4_n305 ) );
INV_X4 _add_1_root_add_136_4_U281  ( .A(_add_1_root_add_136_4_n94 ), .ZN(_add_1_root_add_136_4_n408 ) );
INV_X4 _add_1_root_add_136_4_U280  ( .A(_add_1_root_add_136_4_n225 ), .ZN(_add_1_root_add_136_4_n319 ) );
NOR2_X2 _add_1_root_add_136_4_U279  ( .A1(N93), .A2(Wt[29]), .ZN(_add_1_root_add_136_4_n72 ) );
NOR3_X1 _add_1_root_add_136_4_U278  ( .A1(_add_1_root_add_136_4_n333 ), .A2(_add_1_root_add_136_4_n144 ), .A3(_add_1_root_add_136_4_n330 ), .ZN(_add_1_root_add_136_4_n332 ) );
NOR2_X2 _add_1_root_add_136_4_U277  ( .A1(_add_1_root_add_136_4_n332 ), .A2(_add_1_root_add_136_4_n109 ), .ZN(_add_1_root_add_136_4_n327 ) );
AND2_X2 _add_1_root_add_136_4_U276  ( .A1(N74), .A2(Wt[10]), .ZN(_add_1_root_add_136_4_n70 ) );
NOR2_X2 _add_1_root_add_136_4_U275  ( .A1(_add_1_root_add_136_4_n117 ), .A2(_add_1_root_add_136_4_n118 ), .ZN(_add_1_root_add_136_4_n114 ) );
AND2_X2 _add_1_root_add_136_4_U274  ( .A1(N82), .A2(Wt[18]), .ZN(_add_1_root_add_136_4_n69 ) );
NOR2_X1 _add_1_root_add_136_4_U273  ( .A1(_add_1_root_add_136_4_n330 ), .A2(_add_1_root_add_136_4_n331 ), .ZN(_add_1_root_add_136_4_n329 ) );
NOR2_X2 _add_1_root_add_136_4_U272  ( .A1(Wt[24]), .A2(N88), .ZN(_add_1_root_add_136_4_n195 ) );
AND2_X2 _add_1_root_add_136_4_U271  ( .A1(N89), .A2(Wt[25]), .ZN(_add_1_root_add_136_4_n68 ) );
NOR2_X1 _add_1_root_add_136_4_U270  ( .A1(Wt[2]), .A2(N66), .ZN(_add_1_root_add_136_4_n111 ) );
NOR2_X2 _add_1_root_add_136_4_U269  ( .A1(_add_1_root_add_136_4_n289 ), .A2(_add_1_root_add_136_4_n290 ), .ZN(N128) );
OR2_X2 _add_1_root_add_136_4_U268  ( .A1(N91), .A2(Wt[27]), .ZN(_add_1_root_add_136_4_n164 ) );
NOR2_X1 _add_1_root_add_136_4_U267  ( .A1(_add_1_root_add_136_4_n70 ), .A2(_add_1_root_add_136_4_n393 ), .ZN(_add_1_root_add_136_4_n395 ) );
OR2_X4 _add_1_root_add_136_4_U266  ( .A1(_add_1_root_add_136_4_n183 ), .A2(_add_1_root_add_136_4_n208 ), .ZN(_add_1_root_add_136_4_n64 ) );
XNOR2_X2 _add_1_root_add_136_4_U265  ( .A(_add_1_root_add_136_4_n207 ), .B(_add_1_root_add_136_4_n64 ), .ZN(N152) );
OR2_X4 _add_1_root_add_136_4_U264  ( .A1(_add_1_root_add_136_4_n381 ), .A2(_add_1_root_add_136_4_n384 ), .ZN(_add_1_root_add_136_4_n62 ) );
XNOR2_X2 _add_1_root_add_136_4_U263  ( .A(_add_1_root_add_136_4_n383 ), .B(_add_1_root_add_136_4_n62 ), .ZN(N139) );
NOR2_X2 _add_1_root_add_136_4_U262  ( .A1(_add_1_root_add_136_4_n101 ), .A2(_add_1_root_add_136_4_n102 ), .ZN(_add_1_root_add_136_4_n98 ) );
NOR2_X2 _add_1_root_add_136_4_U261  ( .A1(_add_1_root_add_136_4_n100 ), .A2(_add_1_root_add_136_4_n407 ), .ZN(_add_1_root_add_136_4_n99 ) );
NAND2_X2 _add_1_root_add_136_4_U260  ( .A1(_add_1_root_add_136_4_n324 ),.A2(_add_1_root_add_136_4_n12 ), .ZN(_add_1_root_add_136_4_n322 ) );
NOR2_X2 _add_1_root_add_136_4_U259  ( .A1(_add_1_root_add_136_4_n199 ), .A2(_add_1_root_add_136_4_n200 ), .ZN(_add_1_root_add_136_4_n196 ) );
NOR2_X2 _add_1_root_add_136_4_U258  ( .A1(_add_1_root_add_136_4_n196 ), .A2(_add_1_root_add_136_4_n197 ), .ZN(_add_1_root_add_136_4_n192 ) );
NOR2_X1 _add_1_root_add_136_4_U257  ( .A1(_add_1_root_add_136_4_n68 ), .A2(_add_1_root_add_136_4_n193 ), .ZN(_add_1_root_add_136_4_n185 ) );
NOR2_X2 _add_1_root_add_136_4_U256  ( .A1(_add_1_root_add_136_4_n259 ), .A2(_add_1_root_add_136_4_n260 ), .ZN(_add_1_root_add_136_4_n252 ) );
NOR2_X2 _add_1_root_add_136_4_U255  ( .A1(_add_1_root_add_136_4_n262 ), .A2(_add_1_root_add_136_4_n298 ), .ZN(_add_1_root_add_136_4_n273 ) );
NOR2_X2 _add_1_root_add_136_4_U254  ( .A1(_add_1_root_add_136_4_n111 ), .A2(_add_1_root_add_136_4_n112 ), .ZN(_add_1_root_add_136_4_n108 ) );
NOR2_X2 _add_1_root_add_136_4_U253  ( .A1(_add_1_root_add_136_4_n139 ), .A2(_add_1_root_add_136_4_n128 ), .ZN(_add_1_root_add_136_4_n155 ) );
NOR2_X2 _add_1_root_add_136_4_U252  ( .A1(_add_1_root_add_136_4_n154 ), .A2(_add_1_root_add_136_4_n155 ), .ZN(_add_1_root_add_136_4_n151 ) );
NOR3_X1 _add_1_root_add_136_4_U251  ( .A1(_add_1_root_add_136_4_n129 ), .A2(_add_1_root_add_136_4_n130 ), .A3(_add_1_root_add_136_4_n131 ), .ZN(_add_1_root_add_136_4_n117 ) );
NOR2_X1 _add_1_root_add_136_4_U250  ( .A1(_add_1_root_add_136_4_n8 ), .A2(_add_1_root_add_136_4_n293 ), .ZN(_add_1_root_add_136_4_n292 ) );
NAND3_X1 _add_1_root_add_136_4_U249  ( .A1(_add_1_root_add_136_4_n123 ),.A2(_add_1_root_add_136_4_n124 ), .A3(_add_1_root_add_136_4_n125 ),.ZN(_add_1_root_add_136_4_n122 ) );
NAND3_X1 _add_1_root_add_136_4_U248  ( .A1(_add_1_root_add_136_4_n127 ),.A2(_add_1_root_add_136_4_n124 ), .A3(_add_1_root_add_136_4_n123 ),.ZN(_add_1_root_add_136_4_n119 ) );
NOR2_X2 _add_1_root_add_136_4_U247  ( .A1(_add_1_root_add_136_4_n68 ), .A2(_add_1_root_add_136_4_n175 ), .ZN(_add_1_root_add_136_4_n172 ) );
NOR2_X1 _add_1_root_add_136_4_U246  ( .A1(_add_1_root_add_136_4_n247 ), .A2(_add_1_root_add_136_4_n10 ), .ZN(_add_1_root_add_136_4_n266 ) );
NOR2_X2 _add_1_root_add_136_4_U245  ( .A1(_add_1_root_add_136_4_n217 ), .A2(_add_1_root_add_136_4_n213 ), .ZN(_add_1_root_add_136_4_n216 ) );
NOR2_X2 _add_1_root_add_136_4_U244  ( .A1(_add_1_root_add_136_4_n149 ), .A2(_add_1_root_add_136_4_n150 ), .ZN(_add_1_root_add_136_4_n146 ) );
NOR2_X2 _add_1_root_add_136_4_U243  ( .A1(_add_1_root_add_136_4_n148 ), .A2(_add_1_root_add_136_4_n72 ), .ZN(_add_1_root_add_136_4_n147 ) );
NAND3_X2 _add_1_root_add_136_4_U242  ( .A1(_add_1_root_add_136_4_n134 ),.A2(_add_1_root_add_136_4_n135 ), .A3(_add_1_root_add_136_4_n136 ),.ZN(_add_1_root_add_136_4_n132 ) );
NOR2_X2 _add_1_root_add_136_4_U241  ( .A1(_add_1_root_add_136_4_n313 ), .A2(_add_1_root_add_136_4_n35 ), .ZN(_add_1_root_add_136_4_n308 ) );
NOR2_X2 _add_1_root_add_136_4_U240  ( .A1(_add_1_root_add_136_4_n192 ), .A2(_add_1_root_add_136_4_n193 ), .ZN(_add_1_root_add_136_4_n188 ) );
NOR2_X1 _add_1_root_add_136_4_U239  ( .A1(_add_1_root_add_136_4_n94 ), .A2(_add_1_root_add_136_4_n107 ), .ZN(_add_1_root_add_136_4_n106 ) );
NOR2_X2 _add_1_root_add_136_4_U238  ( .A1(_add_1_root_add_136_4_n108 ), .A2(_add_1_root_add_136_4_n109 ), .ZN(_add_1_root_add_136_4_n105 ) );
NAND3_X2 _add_1_root_add_136_4_U237  ( .A1(_add_1_root_add_136_4_n19 ), .A2(_add_1_root_add_136_4_n40 ), .A3(_add_1_root_add_136_4_n355 ), .ZN(_add_1_root_add_136_4_n353 ) );
NOR2_X2 _add_1_root_add_136_4_U236  ( .A1(_add_1_root_add_136_4_n224 ), .A2(_add_1_root_add_136_4_n225 ), .ZN(_add_1_root_add_136_4_n223 ) );
NAND3_X2 _add_1_root_add_136_4_U235  ( .A1(_add_1_root_add_136_4_n221 ),.A2(_add_1_root_add_136_4_n222 ), .A3(_add_1_root_add_136_4_n220 ),.ZN(_add_1_root_add_136_4_n201 ) );
OR2_X4 _add_1_root_add_136_4_U234  ( .A1(_add_1_root_add_136_4_n1 ), .A2(_add_1_root_add_136_4_n313 ), .ZN(_add_1_root_add_136_4_n56 ) );
XNOR2_X2 _add_1_root_add_136_4_U233  ( .A(_add_1_root_add_136_4_n316 ), .B(_add_1_root_add_136_4_n56 ), .ZN(N144) );
NAND3_X2 _add_1_root_add_136_4_U232  ( .A1(_add_1_root_add_136_4_n220 ),.A2(_add_1_root_add_136_4_n20 ), .A3(_add_1_root_add_136_4_n286 ),.ZN(_add_1_root_add_136_4_n301 ) );
NOR2_X1 _add_1_root_add_136_4_U231  ( .A1(_add_1_root_add_136_4_n130 ), .A2(_add_1_root_add_136_4_n131 ), .ZN(_add_1_root_add_136_4_n161 ) );
INV_X8 _add_1_root_add_136_4_U230  ( .A(_add_1_root_add_136_4_n138 ), .ZN(_add_1_root_add_136_4_n130 ) );
OR2_X4 _add_1_root_add_136_4_U229  ( .A1(N94), .A2(Wt[30]), .ZN(_add_1_root_add_136_4_n124 ) );
NOR2_X1 _add_1_root_add_136_4_U228  ( .A1(Wt[0]), .A2(N64), .ZN(_add_1_root_add_136_4_n290 ) );
OR2_X4 _add_1_root_add_136_4_U227  ( .A1(N76), .A2(Wt[12]), .ZN(_add_1_root_add_136_4_n338 ) );
NOR2_X2 _add_1_root_add_136_4_U226  ( .A1(_add_1_root_add_136_4_n93 ), .A2(_add_1_root_add_136_4_n94 ), .ZN(_add_1_root_add_136_4_n92 ) );
NOR2_X1 _add_1_root_add_136_4_U225  ( .A1(_add_1_root_add_136_4_n183 ), .A2(_add_1_root_add_136_4_n213 ), .ZN(_add_1_root_add_136_4_n198 ) );
INV_X1 _add_1_root_add_136_4_U224  ( .A(_add_1_root_add_136_4_n143 ), .ZN(_add_1_root_add_136_4_n288 ) );
NOR2_X1 _add_1_root_add_136_4_U223  ( .A1(_add_1_root_add_136_4_n288 ), .A2(_add_1_root_add_136_4_n144 ), .ZN(_add_1_root_add_136_4_n287 ) );
OR2_X1 _add_1_root_add_136_4_U222  ( .A1(_add_1_root_add_136_4_n72 ), .A2(_add_1_root_add_136_4_n141 ), .ZN(_add_1_root_add_136_4_n57 ) );
NOR3_X4 _add_1_root_add_136_4_U221  ( .A1(_add_1_root_add_136_4_n54 ), .A2(_add_1_root_add_136_4_n381 ), .A3(_add_1_root_add_136_4_n382 ), .ZN(_add_1_root_add_136_4_n59 ) );
NAND2_X2 _add_1_root_add_136_4_U220  ( .A1(_add_1_root_add_136_4_n333 ),.A2(_add_1_root_add_136_4_n410 ), .ZN(_add_1_root_add_136_4_n51 ) );
NAND2_X4 _add_1_root_add_136_4_U219  ( .A1(_add_1_root_add_136_4_n390 ),.A2(_add_1_root_add_136_4_n375 ), .ZN(_add_1_root_add_136_4_n397 ) );
NOR2_X1 _add_1_root_add_136_4_U218  ( .A1(_add_1_root_add_136_4_n31 ), .A2(_add_1_root_add_136_4_n102 ), .ZN(_add_1_root_add_136_4_n104 ) );
NAND3_X2 _add_1_root_add_136_4_U217  ( .A1(Wt[23]), .A2(_add_1_root_add_136_4_n194 ), .A3(N87), .ZN(_add_1_root_add_136_4_n186 ) );
INV_X4 _add_1_root_add_136_4_U216  ( .A(_add_1_root_add_136_4_n144 ), .ZN(_add_1_root_add_136_4_n50 ) );
NAND3_X2 _add_1_root_add_136_4_U215  ( .A1(_add_1_root_add_136_4_n97 ), .A2(_add_1_root_add_136_4_n95 ), .A3(_add_1_root_add_136_4_n96 ), .ZN(_add_1_root_add_136_4_n93 ) );
NOR2_X1 _add_1_root_add_136_4_U214  ( .A1(_add_1_root_add_136_4_n43 ), .A2(_add_1_root_add_136_4_n107 ), .ZN(_add_1_root_add_136_4_n325 ) );
NAND3_X2 _add_1_root_add_136_4_U213  ( .A1(Wt[2]), .A2(N66), .A3(_add_1_root_add_136_4_n411 ), .ZN(_add_1_root_add_136_4_n95 ) );
NOR2_X2 _add_1_root_add_136_4_U212  ( .A1(_add_1_root_add_136_4_n376 ), .A2(_add_1_root_add_136_4_n380 ), .ZN(_add_1_root_add_136_4_n379 ) );
NAND2_X2 _add_1_root_add_136_4_U211  ( .A1(_add_1_root_add_136_4_n36 ), .A2(Wt[10]), .ZN(_add_1_root_add_136_4_n386 ) );
NOR2_X2 _add_1_root_add_136_4_U210  ( .A1(Wt[10]), .A2(_add_1_root_add_136_4_n36 ), .ZN(_add_1_root_add_136_4_n393 ) );
NOR2_X1 _add_1_root_add_136_4_U209  ( .A1(N74), .A2(Wt[10]), .ZN(_add_1_root_add_136_4_n380 ) );
NAND2_X4 _add_1_root_add_136_4_U208  ( .A1(_add_1_root_add_136_4_n274 ),.A2(_add_1_root_add_136_4_n256 ), .ZN(_add_1_root_add_136_4_n261 ) );
NAND2_X4 _add_1_root_add_136_4_U207  ( .A1(_add_1_root_add_136_4_n48 ), .A2(_add_1_root_add_136_4_n49 ), .ZN(N154) );
NAND2_X4 _add_1_root_add_136_4_U206  ( .A1(_add_1_root_add_136_4_n178 ),.A2(_add_1_root_add_136_4_n179 ), .ZN(_add_1_root_add_136_4_n48 ) );
NOR2_X4 _add_1_root_add_136_4_U205  ( .A1(_add_1_root_add_136_4_n323 ), .A2(_add_1_root_add_136_4_n65 ), .ZN(_add_1_root_add_136_4_n399 ) );
OR2_X4 _add_1_root_add_136_4_U204  ( .A1(_add_1_root_add_136_4_n144 ), .A2(_add_1_root_add_136_4_n333 ), .ZN(_add_1_root_add_136_4_n53 ) );
INV_X2 _add_1_root_add_136_4_U203  ( .A(_add_1_root_add_136_4_n229 ), .ZN(_add_1_root_add_136_4_n236 ) );
NAND2_X4 _add_1_root_add_136_4_U202  ( .A1(_add_1_root_add_136_4_n87 ), .A2(_add_1_root_add_136_4_n88 ), .ZN(_add_1_root_add_136_4_n86 ) );
NOR3_X4 _add_1_root_add_136_4_U201  ( .A1(_add_1_root_add_136_4_n400 ), .A2(_add_1_root_add_136_4_n401 ), .A3(_add_1_root_add_136_4_n402 ), .ZN(_add_1_root_add_136_4_n323 ) );
NOR3_X4 _add_1_root_add_136_4_U200  ( .A1(_add_1_root_add_136_4_n322 ), .A2(_add_1_root_add_136_4_n47 ), .A3(_add_1_root_add_136_4_n65 ), .ZN(_add_1_root_add_136_4_n321 ) );
INV_X4 _add_1_root_add_136_4_U199  ( .A(N85), .ZN(_add_1_root_add_136_4_n267 ) );
INV_X8 _add_1_root_add_136_4_U198  ( .A(_add_1_root_add_136_4_n254 ), .ZN(_add_1_root_add_136_4_n243 ) );
NOR2_X4 _add_1_root_add_136_4_U197  ( .A1(_add_1_root_add_136_4_n243 ), .A2(_add_1_root_add_136_4_n244 ), .ZN(_add_1_root_add_136_4_n206 ) );
NOR2_X2 _add_1_root_add_136_4_U196  ( .A1(Wt[8]), .A2(N72), .ZN(_add_1_root_add_136_4_n382 ) );
NAND2_X4 _add_1_root_add_136_4_U195  ( .A1(_add_1_root_add_136_4_n277 ),.A2(_add_1_root_add_136_4_n278 ), .ZN(_add_1_root_add_136_4_n256 ) );
NOR2_X4 _add_1_root_add_136_4_U194  ( .A1(Wt[2]), .A2(N66), .ZN(_add_1_root_add_136_4_n330 ) );
NAND2_X1 _add_1_root_add_136_4_U193  ( .A1(N86), .A2(Wt[22]), .ZN(_add_1_root_add_136_4_n203 ) );
NAND2_X2 _add_1_root_add_136_4_U192  ( .A1(_add_1_root_add_136_4_n11 ), .A2(_add_1_root_add_136_4_n2 ), .ZN(_add_1_root_add_136_4_n362 ) );
NOR2_X4 _add_1_root_add_136_4_U191  ( .A1(_add_1_root_add_136_4_n269 ), .A2(_add_1_root_add_136_4_n270 ), .ZN(_add_1_root_add_136_4_n265 ) );
NOR2_X4 _add_1_root_add_136_4_U190  ( .A1(N67), .A2(Wt[3]), .ZN(_add_1_root_add_136_4_n107 ) );
NAND2_X4 _add_1_root_add_136_4_U189  ( .A1(_add_1_root_add_136_4_n250 ),.A2(_add_1_root_add_136_4_n251 ), .ZN(_add_1_root_add_136_4_n240 ) );
INV_X8 _add_1_root_add_136_4_U188  ( .A(_add_1_root_add_136_4_n240 ), .ZN(_add_1_root_add_136_4_n246 ) );
NOR2_X4 _add_1_root_add_136_4_U187  ( .A1(_add_1_root_add_136_4_n392 ), .A2(_add_1_root_add_136_4_n397 ), .ZN(_add_1_root_add_136_4_n73 ) );
NOR2_X2 _add_1_root_add_136_4_U186  ( .A1(_add_1_root_add_136_4_n232 ), .A2(_add_1_root_add_136_4_n233 ), .ZN(_add_1_root_add_136_4_n302 ) );
OR3_X2 _add_1_root_add_136_4_U185  ( .A1(_add_1_root_add_136_4_n25 ), .A2(_add_1_root_add_136_4_n232 ), .A3(_add_1_root_add_136_4_n231 ), .ZN(_add_1_root_add_136_4_n60 ) );
NOR2_X4 _add_1_root_add_136_4_U184  ( .A1(_add_1_root_add_136_4_n25 ), .A2(_add_1_root_add_136_4_n363 ), .ZN(_add_1_root_add_136_4_n355 ) );
NAND2_X4 _add_1_root_add_136_4_U183  ( .A1(_add_1_root_add_136_4_n89 ), .A2(_add_1_root_add_136_4_n14 ), .ZN(_add_1_root_add_136_4_n87 ) );
NOR2_X4 _add_1_root_add_136_4_U182  ( .A1(_add_1_root_add_136_4_n295 ), .A2(_add_1_root_add_136_4_n69 ), .ZN(_add_1_root_add_136_4_n291 ) );
INV_X1 _add_1_root_add_136_4_U181  ( .A(_add_1_root_add_136_4_n294 ), .ZN(_add_1_root_add_136_4_n46 ) );
INV_X8 _add_1_root_add_136_4_U180  ( .A(_add_1_root_add_136_4_n261 ), .ZN(_add_1_root_add_136_4_n241 ) );
NAND3_X4 _add_1_root_add_136_4_U179  ( .A1(_add_1_root_add_136_4_n241 ),.A2(_add_1_root_add_136_4_n240 ), .A3(_add_1_root_add_136_4_n239 ),.ZN(_add_1_root_add_136_4_n229 ) );
NAND2_X4 _add_1_root_add_136_4_U178  ( .A1(_add_1_root_add_136_4_n46 ), .A2(Wt[19]), .ZN(_add_1_root_add_136_4_n272 ) );
NAND2_X1 _add_1_root_add_136_4_U177  ( .A1(_add_1_root_add_136_4_n239 ),.A2(_add_1_root_add_136_4_n241 ), .ZN(_add_1_root_add_136_4_n260 ) );
NAND3_X2 _add_1_root_add_136_4_U176  ( .A1(_add_1_root_add_136_4_n315 ),.A2(_add_1_root_add_136_4_n311 ), .A3(_add_1_root_add_136_4_n314 ),.ZN(_add_1_root_add_136_4_n299 ) );
OR2_X2 _add_1_root_add_136_4_U175  ( .A1(_add_1_root_add_136_4_n8 ), .A2(_add_1_root_add_136_4_n281 ), .ZN(_add_1_root_add_136_4_n71 ) );
NAND3_X2 _add_1_root_add_136_4_U174  ( .A1(_add_1_root_add_136_4_n236 ),.A2(_add_1_root_add_136_4_n38 ), .A3(_add_1_root_add_136_4_n238 ),.ZN(_add_1_root_add_136_4_n205 ) );
NOR2_X4 _add_1_root_add_136_4_U173  ( .A1(_add_1_root_add_136_4_n23 ), .A2(_add_1_root_add_136_4_n349 ), .ZN(_add_1_root_add_136_4_n346 ) );
NAND3_X2 _add_1_root_add_136_4_U172  ( .A1(_add_1_root_add_136_4_n356 ),.A2(_add_1_root_add_136_4_n15 ), .A3(_add_1_root_add_136_4_n362 ),.ZN(_add_1_root_add_136_4_n369 ) );
INV_X8 _add_1_root_add_136_4_U171  ( .A(_add_1_root_add_136_4_n83 ), .ZN(_add_1_root_add_136_4_n103 ) );
NOR2_X2 _add_1_root_add_136_4_U170  ( .A1(_add_1_root_add_136_4_n103 ), .A2(_add_1_root_add_136_4_n31 ), .ZN(_add_1_root_add_136_4_n101 ) );
INV_X4 _add_1_root_add_136_4_U169  ( .A(_add_1_root_add_136_4_n392 ), .ZN(_add_1_root_add_136_4_n391 ) );
NAND2_X4 _add_1_root_add_136_4_U168  ( .A1(_add_1_root_add_136_4_n334 ),.A2(_add_1_root_add_136_4_n398 ), .ZN(_add_1_root_add_136_4_n403 ) );
NAND2_X2 _add_1_root_add_136_4_U167  ( .A1(_add_1_root_add_136_4_n267 ),.A2(_add_1_root_add_136_4_n268 ), .ZN(_add_1_root_add_136_4_n45 ) );
NAND2_X4 _add_1_root_add_136_4_U166  ( .A1(_add_1_root_add_136_4_n210 ),.A2(_add_1_root_add_136_4_n209 ), .ZN(_add_1_root_add_136_4_n207 ) );
NAND2_X4 _add_1_root_add_136_4_U165  ( .A1(_add_1_root_add_136_4_n255 ),.A2(_add_1_root_add_136_4_n271 ), .ZN(_add_1_root_add_136_4_n254 ) );
NOR2_X4 _add_1_root_add_136_4_U164  ( .A1(N71), .A2(Wt[7]), .ZN(_add_1_root_add_136_4_n406 ) );
NOR2_X4 _add_1_root_add_136_4_U163  ( .A1(N73), .A2(Wt[9]), .ZN(_add_1_root_add_136_4_n376 ) );
NOR2_X4 _add_1_root_add_136_4_U162  ( .A1(_add_1_root_add_136_4_n246 ), .A2(_add_1_root_add_136_4_n247 ), .ZN(_add_1_root_add_136_4_n245 ) );
NOR2_X2 _add_1_root_add_136_4_U161  ( .A1(_add_1_root_add_136_4_n233 ), .A2(_add_1_root_add_136_4_n335 ), .ZN(_add_1_root_add_136_4_n359 ) );
NOR2_X2 _add_1_root_add_136_4_U160  ( .A1(_add_1_root_add_136_4_n215 ), .A2(_add_1_root_add_136_4_n206 ), .ZN(_add_1_root_add_136_4_n214 ) );
NOR2_X4 _add_1_root_add_136_4_U159  ( .A1(_add_1_root_add_136_4_n227 ), .A2(_add_1_root_add_136_4_n3 ), .ZN(_add_1_root_add_136_4_n320 ) );
NOR2_X4 _add_1_root_add_136_4_U158  ( .A1(_add_1_root_add_136_4_n406 ), .A2(_add_1_root_add_136_4_n401 ), .ZN(_add_1_root_add_136_4_n405 ) );
NAND2_X1 _add_1_root_add_136_4_U157  ( .A1(Wt[3]), .A2(N67), .ZN(_add_1_root_add_136_4_n409 ) );
INV_X4 _add_1_root_add_136_4_U156  ( .A(_add_1_root_add_136_4_n41 ), .ZN(_add_1_root_add_136_4_n42 ) );
NOR2_X1 _add_1_root_add_136_4_U155  ( .A1(_add_1_root_add_136_4_n94 ), .A2(_add_1_root_add_136_4_n329 ), .ZN(_add_1_root_add_136_4_n328 ) );
NAND3_X2 _add_1_root_add_136_4_U154  ( .A1(_add_1_root_add_136_4_n52 ), .A2(_add_1_root_add_136_4_n51 ), .A3(_add_1_root_add_136_4_n50 ), .ZN(_add_1_root_add_136_4_n97 ) );
NAND3_X2 _add_1_root_add_136_4_U153  ( .A1(_add_1_root_add_136_4_n95 ), .A2(_add_1_root_add_136_4_n97 ), .A3(_add_1_root_add_136_4_n408 ), .ZN(_add_1_root_add_136_4_n83 ) );
NAND2_X4 _add_1_root_add_136_4_U152  ( .A1(_add_1_root_add_136_4_n309 ),.A2(_add_1_root_add_136_4_n308 ), .ZN(_add_1_root_add_136_4_n304 ) );
NOR2_X2 _add_1_root_add_136_4_U151  ( .A1(_add_1_root_add_136_4_n75 ), .A2(_add_1_root_add_136_4_n76 ), .ZN(_add_1_root_add_136_4_n74 ) );
NOR2_X4 _add_1_root_add_136_4_U150  ( .A1(_add_1_root_add_136_4_n361 ), .A2(_add_1_root_add_136_4_n362 ), .ZN(_add_1_root_add_136_4_n357 ) );
NOR2_X1 _add_1_root_add_136_4_U149  ( .A1(_add_1_root_add_136_4_n103 ), .A2(_add_1_root_add_136_4_n43 ), .ZN(_add_1_root_add_136_4_n39 ) );
INV_X2 _add_1_root_add_136_4_U148  ( .A(_add_1_root_add_136_4_n303 ), .ZN(_add_1_root_add_136_4_n38 ) );
INV_X4 _add_1_root_add_136_4_U147  ( .A(_add_1_root_add_136_4_n235 ), .ZN(_add_1_root_add_136_4_n37 ) );
INV_X2 _add_1_root_add_136_4_U146  ( .A(_add_1_root_add_136_4_n201 ), .ZN(_add_1_root_add_136_4_n200 ) );
BUF_X16 _add_1_root_add_136_4_U145  ( .A(N74), .Z(_add_1_root_add_136_4_n36 ) );
NAND2_X4 _add_1_root_add_136_4_U144  ( .A1(_add_1_root_add_136_4_n344 ),.A2(_add_1_root_add_136_4_n345 ), .ZN(_add_1_root_add_136_4_n314 ) );
AND3_X2 _add_1_root_add_136_4_U143  ( .A1(_add_1_root_add_136_4_n314 ), .A2(_add_1_root_add_136_4_n311 ), .A3(_add_1_root_add_136_4_n315 ), .ZN(_add_1_root_add_136_4_n35 ) );
NAND2_X1 _add_1_root_add_136_4_U142  ( .A1(_add_1_root_add_136_4_n4 ), .A2(Wt[6]), .ZN(_add_1_root_add_136_4_n88 ) );
INV_X1 _add_1_root_add_136_4_U141  ( .A(_add_1_root_add_136_4_n130 ), .ZN(_add_1_root_add_136_4_n34 ) );
NAND2_X4 _add_1_root_add_136_4_U140  ( .A1(_add_1_root_add_136_4_n211 ),.A2(_add_1_root_add_136_4_n212 ), .ZN(_add_1_root_add_136_4_n210 ) );
NAND2_X4 _add_1_root_add_136_4_U139  ( .A1(_add_1_root_add_136_4_n186 ),.A2(_add_1_root_add_136_4_n187 ), .ZN(_add_1_root_add_136_4_n193 ) );
NOR2_X1 _add_1_root_add_136_4_U138  ( .A1(_add_1_root_add_136_4_n184 ), .A2(_add_1_root_add_136_4_n68 ), .ZN(_add_1_root_add_136_4_n189 ) );
NAND2_X1 _add_1_root_add_136_4_U137  ( .A1(_add_1_root_add_136_4_n223 ),.A2(_add_1_root_add_136_4_n320 ), .ZN(_add_1_root_add_136_4_n222 ) );
INV_X2 _add_1_root_add_136_4_U136  ( .A(_add_1_root_add_136_4_n231 ), .ZN(_add_1_root_add_136_4_n364 ) );
NAND2_X4 _add_1_root_add_136_4_U135  ( .A1(_add_1_root_add_136_4_n264 ),.A2(_add_1_root_add_136_4_n242 ), .ZN(_add_1_root_add_136_4_n298 ) );
NAND2_X4 _add_1_root_add_136_4_U134  ( .A1(_add_1_root_add_136_4_n264 ),.A2(_add_1_root_add_136_4_n242 ), .ZN(_add_1_root_add_136_4_n263 ) );
NAND2_X4 _add_1_root_add_136_4_U133  ( .A1(_add_1_root_add_136_4_n181 ),.A2(_add_1_root_add_136_4_n182 ), .ZN(_add_1_root_add_136_4_n163 ) );
NOR3_X4 _add_1_root_add_136_4_U132  ( .A1(_add_1_root_add_136_4_n183 ), .A2(_add_1_root_add_136_4_n184 ), .A3(_add_1_root_add_136_4_n213 ), .ZN(_add_1_root_add_136_4_n177 ) );
INV_X4 _add_1_root_add_136_4_U131  ( .A(_add_1_root_add_136_4_n103 ), .ZN(_add_1_root_add_136_4_n40 ) );
NAND2_X1 _add_1_root_add_136_4_U130  ( .A1(_add_1_root_add_136_4_n364 ),.A2(_add_1_root_add_136_4_n348 ), .ZN(_add_1_root_add_136_4_n351 ) );
NOR2_X4 _add_1_root_add_136_4_U129  ( .A1(N74), .A2(Wt[10]), .ZN(_add_1_root_add_136_4_n377 ) );
NOR2_X4 _add_1_root_add_136_4_U128  ( .A1(_add_1_root_add_136_4_n262 ), .A2(_add_1_root_add_136_4_n298 ), .ZN(_add_1_root_add_136_4_n259 ) );
AND3_X4 _add_1_root_add_136_4_U127  ( .A1(_add_1_root_add_136_4_n59 ), .A2(_add_1_root_add_136_4_n84 ), .A3(_add_1_root_add_136_4_n85 ), .ZN(_add_1_root_add_136_4_n33 ) );
NAND2_X1 _add_1_root_add_136_4_U126  ( .A1(_add_1_root_add_136_4_n32 ), .A2(Wt[9]), .ZN(_add_1_root_add_136_4_n389 ) );
NAND2_X4 _add_1_root_add_136_4_U125  ( .A1(_add_1_root_add_136_4_n172 ),.A2(_add_1_root_add_136_4_n173 ), .ZN(_add_1_root_add_136_4_n165 ) );
NAND3_X4 _add_1_root_add_136_4_U124  ( .A1(_add_1_root_add_136_4_n163 ),.A2(_add_1_root_add_136_4_n164 ), .A3(_add_1_root_add_136_4_n165 ),.ZN(_add_1_root_add_136_4_n162 ) );
NOR2_X4 _add_1_root_add_136_4_U123  ( .A1(_add_1_root_add_136_4_n73 ), .A2(_add_1_root_add_136_4_n76 ), .ZN(_add_1_root_add_136_4_n396 ) );
NOR2_X4 _add_1_root_add_136_4_U122  ( .A1(_add_1_root_add_136_4_n396 ), .A2(_add_1_root_add_136_4_n75 ), .ZN(_add_1_root_add_136_4_n394 ) );
NOR2_X2 _add_1_root_add_136_4_U121  ( .A1(Wt[24]), .A2(N88), .ZN(_add_1_root_add_136_4_n183 ) );
NAND2_X4 _add_1_root_add_136_4_U120  ( .A1(_add_1_root_add_136_4_n190 ),.A2(_add_1_root_add_136_4_n191 ), .ZN(_add_1_root_add_136_4_n174 ) );
INV_X8 _add_1_root_add_136_4_U119  ( .A(_add_1_root_add_136_4_n174 ), .ZN(_add_1_root_add_136_4_n184 ) );
NAND2_X4 _add_1_root_add_136_4_U118  ( .A1(_add_1_root_add_136_4_n310 ),.A2(_add_1_root_add_136_4_n311 ), .ZN(_add_1_root_add_136_4_n309 ) );
NOR2_X2 _add_1_root_add_136_4_U117  ( .A1(_add_1_root_add_136_4_n252 ), .A2(_add_1_root_add_136_4_n253 ), .ZN(_add_1_root_add_136_4_n248 ) );
NAND2_X1 _add_1_root_add_136_4_U116  ( .A1(_add_1_root_add_136_4_n165 ),.A2(_add_1_root_add_136_4_n163 ), .ZN(_add_1_root_add_136_4_n171 ) );
NAND2_X1 _add_1_root_add_136_4_U115  ( .A1(_add_1_root_add_136_4_n137 ),.A2(_add_1_root_add_136_4_n153 ), .ZN(_add_1_root_add_136_4_n156 ) );
NOR2_X2 _add_1_root_add_136_4_U114  ( .A1(_add_1_root_add_136_4_n156 ), .A2(_add_1_root_add_136_4_n130 ), .ZN(_add_1_root_add_136_4_n149 ) );
NOR2_X2 _add_1_root_add_136_4_U113  ( .A1(_add_1_root_add_136_4_n72 ), .A2(_add_1_root_add_136_4_n139 ), .ZN(_add_1_root_add_136_4_n123 ) );
NAND3_X2 _add_1_root_add_136_4_U112  ( .A1(_add_1_root_add_136_4_n123 ),.A2(_add_1_root_add_136_4_n137 ), .A3(_add_1_root_add_136_4_n34 ),.ZN(_add_1_root_add_136_4_n136 ) );
NAND2_X1 _add_1_root_add_136_4_U111  ( .A1(_add_1_root_add_136_4_n124 ),.A2(_add_1_root_add_136_4_n123 ), .ZN(_add_1_root_add_136_4_n129 ) );
INV_X2 _add_1_root_add_136_4_U110  ( .A(_add_1_root_add_136_4_n195 ), .ZN(_add_1_root_add_136_4_n194 ) );
NOR2_X2 _add_1_root_add_136_4_U109  ( .A1(Wt[4]), .A2(N68), .ZN(_add_1_root_add_136_4_n31 ) );
NAND2_X4 _add_1_root_add_136_4_U108  ( .A1(_add_1_root_add_136_4_n30 ), .A2(_add_1_root_add_136_4_n162 ), .ZN(_add_1_root_add_136_4_n29 ) );
NAND3_X2 _add_1_root_add_136_4_U107  ( .A1(_add_1_root_add_136_4_n18 ), .A2(_add_1_root_add_136_4_n404 ), .A3(_add_1_root_add_136_4_n405 ), .ZN(_add_1_root_add_136_4_n44 ) );
NAND3_X2 _add_1_root_add_136_4_U106  ( .A1(_add_1_root_add_136_4_n18 ), .A2(_add_1_root_add_136_4_n404 ), .A3(_add_1_root_add_136_4_n405 ), .ZN(_add_1_root_add_136_4_n43 ) );
INV_X4 _add_1_root_add_136_4_U105  ( .A(N90), .ZN(_add_1_root_add_136_4_n181 ) );
NOR2_X2 _add_1_root_add_136_4_U104  ( .A1(_add_1_root_add_136_4_n321 ), .A2(_add_1_root_add_136_4_n17 ), .ZN(_add_1_root_add_136_4_n227 ) );
NAND2_X1 _add_1_root_add_136_4_U103  ( .A1(_add_1_root_add_136_4_n284 ),.A2(_add_1_root_add_136_4_n285 ), .ZN(_add_1_root_add_136_4_n283 ) );
NAND2_X1 _add_1_root_add_136_4_U102  ( .A1(_add_1_root_add_136_4_n42 ), .A2(Wt[5]), .ZN(_add_1_root_add_136_4_n91 ) );
OR2_X4 _add_1_root_add_136_4_U101  ( .A1(_add_1_root_add_136_4_n184 ), .A2(_add_1_root_add_136_4_n185 ), .ZN(_add_1_root_add_136_4_n27 ) );
INV_X4 _add_1_root_add_136_4_U100  ( .A(_add_1_root_add_136_4_n26 ), .ZN(_add_1_root_add_136_4_n178 ) );
NAND2_X2 _add_1_root_add_136_4_U99  ( .A1(_add_1_root_add_136_4_n27 ), .A2(_add_1_root_add_136_4_n28 ), .ZN(_add_1_root_add_136_4_n26 ) );
NOR2_X4 _add_1_root_add_136_4_U98  ( .A1(Wt[13]), .A2(N77), .ZN(_add_1_root_add_136_4_n25 ) );
INV_X2 _add_1_root_add_136_4_U97  ( .A(_add_1_root_add_136_4_n348 ), .ZN(_add_1_root_add_136_4_n347 ) );
NOR2_X4 _add_1_root_add_136_4_U96  ( .A1(_add_1_root_add_136_4_n346 ), .A2(_add_1_root_add_136_4_n347 ), .ZN(_add_1_root_add_136_4_n343 ) );
NOR2_X4 _add_1_root_add_136_4_U95  ( .A1(_add_1_root_add_136_4_n243 ), .A2(_add_1_root_add_136_4_n244 ), .ZN(_add_1_root_add_136_4_n24 ) );
INV_X4 _add_1_root_add_136_4_U94  ( .A(_add_1_root_add_136_4_n237 ), .ZN(_add_1_root_add_136_4_n303 ) );
INV_X2 _add_1_root_add_136_4_U93  ( .A(_add_1_root_add_136_4_n91 ), .ZN(_add_1_root_add_136_4_n100 ) );
NOR2_X1 _add_1_root_add_136_4_U92  ( .A1(Wt[14]), .A2(N78), .ZN(_add_1_root_add_136_4_n231 ) );
NAND2_X2 _add_1_root_add_136_4_U91  ( .A1(_add_1_root_add_136_4_n177 ), .A2(_add_1_root_add_136_4_n138 ), .ZN(_add_1_root_add_136_4_n28 ) );
NOR2_X2 _add_1_root_add_136_4_U90  ( .A1(_add_1_root_add_136_4_n282 ), .A2(_add_1_root_add_136_4_n283 ), .ZN(_add_1_root_add_136_4_n279 ) );
INV_X2 _add_1_root_add_136_4_U89  ( .A(_add_1_root_add_136_4_n206 ), .ZN(_add_1_root_add_136_4_n202 ) );
CLKBUF_X3 _add_1_root_add_136_4_U88  ( .A(_add_1_root_add_136_4_n323 ), .Z(_add_1_root_add_136_4_n47 ) );
INV_X8 _add_1_root_add_136_4_U87  ( .A(_add_1_root_add_136_4_n350 ), .ZN(_add_1_root_add_136_4_n349 ) );
INV_X4 _add_1_root_add_136_4_U86  ( .A(_add_1_root_add_136_4_n22 ), .ZN(_add_1_root_add_136_4_n204 ) );
NOR2_X2 _add_1_root_add_136_4_U85  ( .A1(_add_1_root_add_136_4_n242 ), .A2(_add_1_root_add_136_4_n229 ), .ZN(_add_1_root_add_136_4_n22 ) );
AND2_X2 _add_1_root_add_136_4_U84  ( .A1(_add_1_root_add_136_4_n256 ), .A2(_add_1_root_add_136_4_n258 ), .ZN(_add_1_root_add_136_4_n21 ) );
AND2_X2 _add_1_root_add_136_4_U83  ( .A1(_add_1_root_add_136_4_n59 ), .A2(_add_1_root_add_136_4_n13 ), .ZN(_add_1_root_add_136_4_n19 ) );
OR2_X2 _add_1_root_add_136_4_U82  ( .A1(Wt[4]), .A2(N68), .ZN(_add_1_root_add_136_4_n18 ) );
INV_X2 _add_1_root_add_136_4_U81  ( .A(_add_1_root_add_136_4_n333 ), .ZN(_add_1_root_add_136_4_n289 ) );
NOR2_X4 _add_1_root_add_136_4_U80  ( .A1(_add_1_root_add_136_4_n6 ), .A2(Wt[7]), .ZN(_add_1_root_add_136_4_n17 ) );
NOR2_X4 _add_1_root_add_136_4_U79  ( .A1(_add_1_root_add_136_4_n273 ), .A2(_add_1_root_add_136_4_n261 ), .ZN(_add_1_root_add_136_4_n269 ) );
NAND2_X2 _add_1_root_add_136_4_U78  ( .A1(_add_1_root_add_136_4_n13 ), .A2(_add_1_root_add_136_4_n40 ), .ZN(_add_1_root_add_136_4_n82 ) );
NOR2_X4 _add_1_root_add_136_4_U77  ( .A1(_add_1_root_add_136_4_n374 ), .A2(_add_1_root_add_136_4_n70 ), .ZN(_add_1_root_add_136_4_n373 ) );
NAND2_X4 _add_1_root_add_136_4_U76  ( .A1(N75), .A2(Wt[11]), .ZN(_add_1_root_add_136_4_n372 ) );
INV_X4 _add_1_root_add_136_4_U75  ( .A(_add_1_root_add_136_4_n107 ), .ZN(_add_1_root_add_136_4_n411 ) );
NAND2_X4 _add_1_root_add_136_4_U74  ( .A1(_add_1_root_add_136_4_n58 ), .A2(_add_1_root_add_136_4_n91 ), .ZN(_add_1_root_add_136_4_n89 ) );
INV_X4 _add_1_root_add_136_4_U73  ( .A(_add_1_root_add_136_4_n377 ), .ZN(_add_1_root_add_136_4_n378 ) );
NOR3_X4 _add_1_root_add_136_4_U72  ( .A1(_add_1_root_add_136_4_n376 ), .A2(_add_1_root_add_136_4_n375 ), .A3(_add_1_root_add_136_4_n377 ), .ZN(_add_1_root_add_136_4_n374 ) );
NOR2_X2 _add_1_root_add_136_4_U71  ( .A1(_add_1_root_add_136_4_n247 ), .A2(_add_1_root_add_136_4_n243 ), .ZN(_add_1_root_add_136_4_n253 ) );
NOR2_X2 _add_1_root_add_136_4_U70  ( .A1(_add_1_root_add_136_4_n215 ), .A2(_add_1_root_add_136_4_n246 ), .ZN(_add_1_root_add_136_4_n249 ) );
NAND2_X2 _add_1_root_add_136_4_U69  ( .A1(_add_1_root_add_136_4_n26 ), .A2(_add_1_root_add_136_4_n180 ), .ZN(_add_1_root_add_136_4_n49 ) );
NOR2_X2 _add_1_root_add_136_4_U68  ( .A1(_add_1_root_add_136_4_n161 ), .A2(_add_1_root_add_136_4_n29 ), .ZN(_add_1_root_add_136_4_n157 ) );
NOR2_X2 _add_1_root_add_136_4_U67  ( .A1(_add_1_root_add_136_4_n139 ), .A2(_add_1_root_add_136_4_n154 ), .ZN(_add_1_root_add_136_4_n158 ) );
NOR2_X2 _add_1_root_add_136_4_U66  ( .A1(_add_1_root_add_136_4_n107 ), .A2(_add_1_root_add_136_4_n330 ), .ZN(_add_1_root_add_136_4_n52 ) );
NOR2_X2 _add_1_root_add_136_4_U65  ( .A1(_add_1_root_add_136_4_n296 ), .A2(_add_1_root_add_136_4_n275 ), .ZN(_add_1_root_add_136_4_n295 ) );
INV_X4 _add_1_root_add_136_4_U64  ( .A(_add_1_root_add_136_4_n127 ), .ZN(_add_1_root_add_136_4_n30 ) );
NOR2_X4 _add_1_root_add_136_4_U63  ( .A1(N78), .A2(Wt[14]), .ZN(_add_1_root_add_136_4_n342 ) );
NOR2_X4 _add_1_root_add_136_4_U62  ( .A1(_add_1_root_add_136_4_n262 ), .A2(_add_1_root_add_136_4_n263 ), .ZN(_add_1_root_add_136_4_n296 ) );
NOR2_X2 _add_1_root_add_136_4_U61  ( .A1(_add_1_root_add_136_4_n262 ), .A2(_add_1_root_add_136_4_n263 ), .ZN(_add_1_root_add_136_4_n282 ) );
BUF_X8 _add_1_root_add_136_4_U60  ( .A(N73), .Z(_add_1_root_add_136_4_n32 ));
INV_X8 _add_1_root_add_136_4_U59  ( .A(_add_1_root_add_136_4_n342 ), .ZN(_add_1_root_add_136_4_n341 ) );
NOR3_X4 _add_1_root_add_136_4_U58  ( .A1(_add_1_root_add_136_4_n229 ), .A2(_add_1_root_add_136_4_n230 ), .A3(_add_1_root_add_136_4_n60 ), .ZN(_add_1_root_add_136_4_n221 ) );
NOR2_X4 _add_1_root_add_136_4_U57  ( .A1(Wt[23]), .A2(N87), .ZN(_add_1_root_add_136_4_n213 ) );
NAND2_X4 _add_1_root_add_136_4_U56  ( .A1(_add_1_root_add_136_4_n280 ), .A2(_add_1_root_add_136_4_n256 ), .ZN(_add_1_root_add_136_4_n271 ) );
NAND2_X1 _add_1_root_add_136_4_U55  ( .A1(_add_1_root_add_136_4_n163 ), .A2(_add_1_root_add_136_4_n176 ), .ZN(_add_1_root_add_136_4_n180 ) );
INV_X2 _add_1_root_add_136_4_U54  ( .A(_add_1_root_add_136_4_n180 ), .ZN(_add_1_root_add_136_4_n179 ) );
NAND2_X4 _add_1_root_add_136_4_U53  ( .A1(N72), .A2(Wt[8]), .ZN(_add_1_root_add_136_4_n375 ) );
NOR2_X2 _add_1_root_add_136_4_U52  ( .A1(Wt[9]), .A2(_add_1_root_add_136_4_n32 ), .ZN(_add_1_root_add_136_4_n76 ) );
AND2_X2 _add_1_root_add_136_4_U51  ( .A1(_add_1_root_add_136_4_n339 ), .A2(_add_1_root_add_136_4_n314 ), .ZN(_add_1_root_add_136_4_n16 ) );
NAND2_X4 _add_1_root_add_136_4_U50  ( .A1(N64), .A2(Wt[0]), .ZN(_add_1_root_add_136_4_n333 ) );
NAND2_X1 _add_1_root_add_136_4_U49  ( .A1(_add_1_root_add_136_4_n59 ), .A2(_add_1_root_add_136_4_n39 ), .ZN(_add_1_root_add_136_4_n15 ) );
NOR2_X2 _add_1_root_add_136_4_U48  ( .A1(_add_1_root_add_136_4_n80 ), .A2(_add_1_root_add_136_4_n382 ), .ZN(_add_1_root_add_136_4_n79 ) );
NAND2_X2 _add_1_root_add_136_4_U47  ( .A1(_add_1_root_add_136_4_n193 ), .A2(_add_1_root_add_136_4_n174 ), .ZN(_add_1_root_add_136_4_n173 ) );
NOR2_X2 _add_1_root_add_136_4_U46  ( .A1(_add_1_root_add_136_4_n275 ), .A2(_add_1_root_add_136_4_n8 ), .ZN(_add_1_root_add_136_4_n274 ) );
OR2_X1 _add_1_root_add_136_4_U45  ( .A1(Wt[6]), .A2(_add_1_root_add_136_4_n4 ), .ZN(_add_1_root_add_136_4_n14 ) );
OR3_X2 _add_1_root_add_136_4_U44  ( .A1(_add_1_root_add_136_4_n92 ), .A2(_add_1_root_add_136_4_n31 ), .A3(_add_1_root_add_136_4_n407 ), .ZN(_add_1_root_add_136_4_n58 ) );
NAND2_X4 _add_1_root_add_136_4_U43  ( .A1(_add_1_root_add_136_4_n369 ), .A2(_add_1_root_add_136_4_n338 ), .ZN(_add_1_root_add_136_4_n368 ) );
NAND2_X4 _add_1_root_add_136_4_U42  ( .A1(_add_1_root_add_136_4_n368 ), .A2(_add_1_root_add_136_4_n335 ), .ZN(_add_1_root_add_136_4_n365 ) );
INV_X2 _add_1_root_add_136_4_U41  ( .A(N69), .ZN(_add_1_root_add_136_4_n41 ));
NOR2_X4 _add_1_root_add_136_4_U40  ( .A1(N75), .A2(Wt[11]), .ZN(_add_1_root_add_136_4_n381 ) );
NOR2_X2 _add_1_root_add_136_4_U39  ( .A1(_add_1_root_add_136_4_n275 ), .A2(_add_1_root_add_136_4_n69 ), .ZN(_add_1_root_add_136_4_n297 ) );
INV_X2 _add_1_root_add_136_4_U38  ( .A(_add_1_root_add_136_4_n275 ), .ZN(_add_1_root_add_136_4_n284 ) );
INV_X4 _add_1_root_add_136_4_U37  ( .A(_add_1_root_add_136_4_n44 ), .ZN(_add_1_root_add_136_4_n334 ) );
CLKBUF_X2 _add_1_root_add_136_4_U36  ( .A(_add_1_root_add_136_4_n334 ), .Z(_add_1_root_add_136_4_n13 ) );
INV_X4 _add_1_root_add_136_4_U35  ( .A(_add_1_root_add_136_4_n12 ), .ZN(_add_1_root_add_136_4_n67 ) );
NAND2_X2 _add_1_root_add_136_4_U34  ( .A1(Wt[7]), .A2(N71), .ZN(_add_1_root_add_136_4_n12 ) );
OR2_X1 _add_1_root_add_136_4_U33  ( .A1(Wt[11]), .A2(N75), .ZN(_add_1_root_add_136_4_n11 ) );
AND2_X2 _add_1_root_add_136_4_U32  ( .A1(N85), .A2(Wt[21]), .ZN(_add_1_root_add_136_4_n10 ) );
NAND2_X4 _add_1_root_add_136_4_U31  ( .A1(_add_1_root_add_136_4_n71 ), .A2(_add_1_root_add_136_4_n272 ), .ZN(_add_1_root_add_136_4_n280 ) );
OR2_X4 _add_1_root_add_136_4_U30  ( .A1(_add_1_root_add_136_4_n17 ), .A2(_add_1_root_add_136_4_n67 ), .ZN(_add_1_root_add_136_4_n9 ) );
INV_X2 _add_1_root_add_136_4_U29  ( .A(_add_1_root_add_136_4_n111 ), .ZN(_add_1_root_add_136_4_n145 ) );
NAND2_X2 _add_1_root_add_136_4_U28  ( .A1(_add_1_root_add_136_4_n388 ), .A2(_add_1_root_add_136_4_n387 ), .ZN(_add_1_root_add_136_4_n385 ) );
INV_X2 _add_1_root_add_136_4_U27  ( .A(N83), .ZN(_add_1_root_add_136_4_n294 ) );
INV_X4 _add_1_root_add_136_4_U26  ( .A(_add_1_root_add_136_4_n8 ), .ZN(_add_1_root_add_136_4_n285 ) );
NOR2_X4 _add_1_root_add_136_4_U25  ( .A1(N83), .A2(Wt[19]), .ZN(_add_1_root_add_136_4_n8 ) );
INV_X4 _add_1_root_add_136_4_U24  ( .A(_add_1_root_add_136_4_n33 ), .ZN(_add_1_root_add_136_4_n356 ) );
INV_X1 _add_1_root_add_136_4_U23  ( .A(_add_1_root_add_136_4_n306 ), .ZN(_add_1_root_add_136_4_n7 ) );
NOR2_X1 _add_1_root_add_136_4_U22  ( .A1(_add_1_root_add_136_4_n76 ), .A2(_add_1_root_add_136_4_n393 ), .ZN(_add_1_root_add_136_4_n387 ) );
NAND2_X2 _add_1_root_add_136_4_U21  ( .A1(_add_1_root_add_136_4_n385 ), .A2(_add_1_root_add_136_4_n386 ), .ZN(_add_1_root_add_136_4_n383 ) );
NOR2_X2 _add_1_root_add_136_4_U20  ( .A1(_add_1_root_add_136_4_n257 ), .A2(_add_1_root_add_136_4_n10 ), .ZN(_add_1_root_add_136_4_n255 ) );
INV_X4 _add_1_root_add_136_4_U19  ( .A(_add_1_root_add_136_4_n5 ), .ZN(_add_1_root_add_136_4_n6 ) );
INV_X1 _add_1_root_add_136_4_U18  ( .A(N71), .ZN(_add_1_root_add_136_4_n5 ));
INV_X2 _add_1_root_add_136_4_U17  ( .A(_add_1_root_add_136_4_n379 ), .ZN(_add_1_root_add_136_4_n54 ) );
BUF_X16 _add_1_root_add_136_4_U16  ( .A(N70), .Z(_add_1_root_add_136_4_n4 ));
NOR2_X2 _add_1_root_add_136_4_U15  ( .A1(N69), .A2(Wt[5]), .ZN(_add_1_root_add_136_4_n400 ) );
NOR2_X2 _add_1_root_add_136_4_U14  ( .A1(N69), .A2(Wt[5]), .ZN(_add_1_root_add_136_4_n407 ) );
AND3_X2 _add_1_root_add_136_4_U13  ( .A1(_add_1_root_add_136_4_n302 ), .A2(_add_1_root_add_136_4_n364 ), .A3(_add_1_root_add_136_4_n234 ), .ZN(_add_1_root_add_136_4_n20 ) );
OR2_X4 _add_1_root_add_136_4_U12  ( .A1(N70), .A2(Wt[6]), .ZN(_add_1_root_add_136_4_n66 ) );
INV_X4 _add_1_root_add_136_4_U11  ( .A(_add_1_root_add_136_4_n301 ), .ZN(_add_1_root_add_136_4_n262 ) );
NAND3_X2 _add_1_root_add_136_4_U10  ( .A1(Wt[9]), .A2(_add_1_root_add_136_4_n378 ), .A3(N73), .ZN(_add_1_root_add_136_4_n371 ) );
NAND3_X1 _add_1_root_add_136_4_U9  ( .A1(_add_1_root_add_136_4_n373 ), .A2(_add_1_root_add_136_4_n372 ), .A3(_add_1_root_add_136_4_n371 ), .ZN(_add_1_root_add_136_4_n228 ) );
NAND3_X2 _add_1_root_add_136_4_U8  ( .A1(_add_1_root_add_136_4_n373 ), .A2(_add_1_root_add_136_4_n372 ), .A3(_add_1_root_add_136_4_n371 ), .ZN(_add_1_root_add_136_4_n3 ) );
NAND3_X1 _add_1_root_add_136_4_U7  ( .A1(_add_1_root_add_136_4_n373 ), .A2(_add_1_root_add_136_4_n372 ), .A3(_add_1_root_add_136_4_n371 ), .ZN(_add_1_root_add_136_4_n2 ) );
INV_X2 _add_1_root_add_136_4_U6  ( .A(_add_1_root_add_136_4_n341 ), .ZN(_add_1_root_add_136_4_n23 ) );
AND2_X4 _add_1_root_add_136_4_U5  ( .A1(N70), .A2(Wt[6]), .ZN(_add_1_root_add_136_4_n65 ) );
NAND2_X2 _add_1_root_add_136_4_U4  ( .A1(N82), .A2(Wt[18]), .ZN(_add_1_root_add_136_4_n281 ) );
INV_X4 _add_1_root_add_136_4_U3  ( .A(_add_1_root_add_136_4_n1 ), .ZN(_add_1_root_add_136_4_n311 ) );
NOR2_X4 _add_1_root_add_136_4_U2  ( .A1(N80), .A2(Wt[16]), .ZN(_add_1_root_add_136_4_n1 ) );
NAND2_X2 _add_512_U458  ( .A1(next_A[2]), .A2(H0[2]), .ZN(_add_512_n426 ) );
NAND2_X2 _add_512_U457  ( .A1(H0[3]), .A2(next_A[3]), .ZN(_add_512_n100 ) );
NAND2_X2 _add_512_U456  ( .A1(H0[0]), .A2(next_A[0]), .ZN(_add_512_n424 ) );
NAND2_X2 _add_512_U455  ( .A1(H0[1]), .A2(next_A[1]), .ZN(_add_512_n425 ) );
NAND2_X2 _add_512_U454  ( .A1(_add_512_n424 ), .A2(_add_512_n425 ), .ZN(_add_512_n422 ) );
NOR2_X4 _add_512_U453  ( .A1(next_A[8]), .A2(H0[8]), .ZN(_add_512_n78 ) );
NOR2_X4 _add_512_U452  ( .A1(next_A[9]), .A2(H0[9]), .ZN(_add_512_n73 ) );
INV_X4 _add_512_U451  ( .A(_add_512_n412 ), .ZN(_add_512_n417 ) );
NOR2_X4 _add_512_U450  ( .A1(next_A[5]), .A2(H0[5]), .ZN(_add_512_n105 ) );
INV_X4 _add_512_U449  ( .A(_add_512_n105 ), .ZN(_add_512_n418 ) );
INV_X4 _add_512_U448  ( .A(_add_512_n104 ), .ZN(_add_512_n419 ) );
INV_X4 _add_512_U447  ( .A(_add_512_n93 ), .ZN(_add_512_n337 ) );
INV_X4 _add_512_U446  ( .A(_add_512_n87 ), .ZN(_add_512_n336 ) );
NAND2_X2 _add_512_U445  ( .A1(H0[8]), .A2(next_A[8]), .ZN(_add_512_n84 ) );
NAND2_X2 _add_512_U444  ( .A1(H0[9]), .A2(next_A[9]), .ZN(_add_512_n74 ) );
NAND2_X2 _add_512_U443  ( .A1(H0[7]), .A2(next_A[7]), .ZN(_add_512_n90 ) );
NAND2_X2 _add_512_U442  ( .A1(H0[6]), .A2(next_A[6]), .ZN(_add_512_n92 ) );
NAND2_X2 _add_512_U441  ( .A1(H0[4]), .A2(next_A[4]), .ZN(_add_512_n416 ) );
NAND2_X2 _add_512_U440  ( .A1(_add_512_n416 ), .A2(_add_512_n94 ), .ZN(_add_512_n415 ) );
NAND2_X2 _add_512_U439  ( .A1(_add_512_n414 ), .A2(_add_512_n415 ), .ZN(_add_512_n413 ) );
NOR2_X4 _add_512_U438  ( .A1(next_A[10]), .A2(H0[10]), .ZN(_add_512_n334 ));
XNOR2_X2 _add_512_U437  ( .A(_add_512_n407 ), .B(_add_512_n408 ), .ZN(N862));
NAND2_X2 _add_512_U436  ( .A1(H0[11]), .A2(next_A[11]), .ZN(_add_512_n400 ));
INV_X4 _add_512_U435  ( .A(_add_512_n400 ), .ZN(_add_512_n405 ) );
XNOR2_X2 _add_512_U434  ( .A(_add_512_n403 ), .B(_add_512_n404 ), .ZN(N863));
INV_X4 _add_512_U433  ( .A(_add_512_n333 ), .ZN(_add_512_n401 ) );
NOR2_X4 _add_512_U432  ( .A1(_add_512_n78 ), .A2(_add_512_n334 ), .ZN(_add_512_n402 ) );
NAND2_X2 _add_512_U431  ( .A1(_add_512_n399 ), .A2(_add_512_n400 ), .ZN(_add_512_n395 ) );
NOR3_X4 _add_512_U430  ( .A1(_add_512_n397 ), .A2(_add_512_n396 ), .A3(_add_512_n395 ), .ZN(_add_512_n205 ) );
INV_X4 _add_512_U429  ( .A(_add_512_n86 ), .ZN(_add_512_n394 ) );
XNOR2_X2 _add_512_U428  ( .A(_add_512_n391 ), .B(_add_512_n392 ), .ZN(N864));
INV_X4 _add_512_U427  ( .A(_add_512_n375 ), .ZN(_add_512_n384 ) );
XNOR2_X2 _add_512_U426  ( .A(_add_512_n388 ), .B(_add_512_n389 ), .ZN(N865));
INV_X4 _add_512_U425  ( .A(H0[14]), .ZN(_add_512_n381 ) );
XNOR2_X2 _add_512_U424  ( .A(_add_512_n378 ), .B(_add_512_n379 ), .ZN(N866));
NAND2_X2 _add_512_U423  ( .A1(_add_512_n60 ), .A2(_add_512_n351 ), .ZN(_add_512_n374 ) );
INV_X4 _add_512_U422  ( .A(H0[15]), .ZN(_add_512_n371 ) );
INV_X4 _add_512_U421  ( .A(next_A[15]), .ZN(_add_512_n372 ) );
XNOR2_X2 _add_512_U420  ( .A(_add_512_n368 ), .B(_add_512_n369 ), .ZN(N867));
NAND2_X2 _add_512_U419  ( .A1(H0[16]), .A2(n13108), .ZN(_add_512_n327 ) );
NOR2_X4 _add_512_U418  ( .A1(n13108), .A2(H0[16]), .ZN(_add_512_n320 ) );
NAND2_X2 _add_512_U417  ( .A1(_add_512_n327 ), .A2(_add_512_n329 ), .ZN(_add_512_n330 ) );
NAND2_X2 _add_512_U416  ( .A1(_add_512_n364 ), .A2(_add_512_n365 ), .ZN(_add_512_n340 ) );
INV_X4 _add_512_U415  ( .A(_add_512_n334 ), .ZN(_add_512_n361 ) );
INV_X4 _add_512_U414  ( .A(_add_512_n78 ), .ZN(_add_512_n362 ) );
NOR3_X4 _add_512_U413  ( .A1(_add_512_n360 ), .A2(_add_512_n335 ), .A3(_add_512_n336 ), .ZN(_add_512_n355 ) );
NAND4_X2 _add_512_U412  ( .A1(H0[4]), .A2(next_A[4]), .A3(_add_512_n418 ),.A4(_add_512_n93 ), .ZN(_add_512_n358 ) );
NAND3_X4 _add_512_U411  ( .A1(_add_512_n354 ), .A2(_add_512_n355 ), .A3(_add_512_n356 ), .ZN(_add_512_n200 ) );
INV_X4 _add_512_U410  ( .A(_add_512_n165 ), .ZN(_add_512_n347 ) );
NAND4_X2 _add_512_U409  ( .A1(H0[0]), .A2(next_A[0]), .A3(_add_512_n347 ),.A4(_add_512_n166 ), .ZN(_add_512_n343 ) );
INV_X4 _add_512_U408  ( .A(_add_512_n100 ), .ZN(_add_512_n114 ) );
NOR2_X4 _add_512_U407  ( .A1(_add_512_n335 ), .A2(_add_512_n332 ), .ZN(_add_512_n213 ) );
NAND2_X2 _add_512_U406  ( .A1(_add_512_n213 ), .A2(_add_512_n385 ), .ZN(_add_512_n342 ) );
XNOR2_X2 _add_512_U405  ( .A(_add_512_n330 ), .B(_add_512_n53 ), .ZN(N868));
NAND2_X2 _add_512_U404  ( .A1(_add_512_n53 ), .A2(_add_512_n329 ), .ZN(_add_512_n328 ) );
INV_X4 _add_512_U403  ( .A(H0[17]), .ZN(_add_512_n325 ) );
XNOR2_X2 _add_512_U402  ( .A(_add_512_n323 ), .B(_add_512_n324 ), .ZN(N869));
INV_X4 _add_512_U401  ( .A(_add_512_n68 ), .ZN(_add_512_n319 ) );
NOR2_X4 _add_512_U400  ( .A1(_add_512_n319 ), .A2(_add_512_n320 ), .ZN(_add_512_n312 ) );
NAND2_X2 _add_512_U399  ( .A1(_add_512_n53 ), .A2(_add_512_n23 ), .ZN(_add_512_n318 ) );
INV_X4 _add_512_U398  ( .A(H0[18]), .ZN(_add_512_n315 ) );
NAND2_X2 _add_512_U397  ( .A1(H0[18]), .A2(next_A[18]), .ZN(_add_512_n192 ));
NAND4_X2 _add_512_U396  ( .A1(_add_512_n307 ), .A2(_add_512_n31 ), .A3(_add_512_n271 ), .A4(_add_512_n308 ), .ZN(_add_512_n306 ) );
NOR2_X4 _add_512_U395  ( .A1(_add_512_n304 ), .A2(_add_512_n303 ), .ZN(_add_512_n285 ) );
INV_X4 _add_512_U394  ( .A(_add_512_n425 ), .ZN(_add_512_n301 ) );
XNOR2_X2 _add_512_U393  ( .A(_add_512_n424 ), .B(_add_512_n300 ), .ZN(N853));
NAND2_X2 _add_512_U392  ( .A1(next_A[20]), .A2(H0[20]), .ZN(_add_512_n295 ));
INV_X4 _add_512_U391  ( .A(_add_512_n295 ), .ZN(_add_512_n258 ) );
XNOR2_X2 _add_512_U390  ( .A(_add_512_n297 ), .B(_add_512_n298 ), .ZN(N872));
NOR2_X4 _add_512_U389  ( .A1(_add_512_n8 ), .A2(_add_512_n296 ), .ZN(_add_512_n257 ) );
INV_X4 _add_512_U388  ( .A(H0[21]), .ZN(_add_512_n290 ) );
XNOR2_X2 _add_512_U387  ( .A(_add_512_n288 ), .B(_add_512_n289 ), .ZN(N873));
INV_X4 _add_512_U386  ( .A(_add_512_n282 ), .ZN(_add_512_n280 ) );
INV_X4 _add_512_U385  ( .A(_add_512_n191 ), .ZN(_add_512_n254 ) );
INV_X4 _add_512_U384  ( .A(H0[22]), .ZN(_add_512_n276 ) );
INV_X4 _add_512_U383  ( .A(_add_512_n256 ), .ZN(_add_512_n275 ) );
XNOR2_X2 _add_512_U382  ( .A(_add_512_n273 ), .B(_add_512_n274 ), .ZN(N874));
INV_X4 _add_512_U381  ( .A(_add_512_n192 ), .ZN(_add_512_n267 ) );
NAND2_X2 _add_512_U380  ( .A1(_add_512_n203 ), .A2(_add_512_n200 ), .ZN(_add_512_n269 ) );
NOR4_X4 _add_512_U379  ( .A1(_add_512_n268 ), .A2(_add_512_n269 ), .A3(_add_512_n189 ), .A4(_add_512_n310 ), .ZN(_add_512_n259 ) );
INV_X4 _add_512_U378  ( .A(_add_512_n264 ), .ZN(_add_512_n263 ) );
INV_X4 _add_512_U377  ( .A(_add_512_n218 ), .ZN(_add_512_n262 ) );
NOR2_X4 _add_512_U376  ( .A1(_add_512_n259 ), .A2(_add_512_n260 ), .ZN(_add_512_n253 ) );
NAND3_X4 _add_512_U375  ( .A1(_add_512_n37 ), .A2(_add_512_n256 ), .A3(_add_512_n66 ), .ZN(_add_512_n219 ) );
NOR2_X4 _add_512_U374  ( .A1(_add_512_n253 ), .A2(_add_512_n51 ), .ZN(_add_512_n229 ) );
NOR2_X4 _add_512_U373  ( .A1(next_A[23]), .A2(H0[23]), .ZN(_add_512_n240 ));
INV_X4 _add_512_U372  ( .A(H0[24]), .ZN(_add_512_n247 ) );
INV_X4 _add_512_U371  ( .A(next_A[24]), .ZN(_add_512_n248 ) );
NAND2_X2 _add_512_U370  ( .A1(H0[25]), .A2(next_A[25]), .ZN(_add_512_n228 ));
XNOR2_X2 _add_512_U369  ( .A(_add_512_n242 ), .B(_add_512_n243 ), .ZN(N877));
NOR3_X4 _add_512_U368  ( .A1(_add_512_n240 ), .A2(_add_512_n69 ), .A3(_add_512_n241 ), .ZN(_add_512_n230 ) );
INV_X4 _add_512_U367  ( .A(H0[26]), .ZN(_add_512_n231 ) );
INV_X4 _add_512_U366  ( .A(H0[27]), .ZN(_add_512_n221 ) );
XNOR2_X2 _add_512_U365  ( .A(_add_512_n220 ), .B(_add_512_n10 ), .ZN(N879));
NAND2_X2 _add_512_U364  ( .A1(_add_512_n214 ), .A2(_add_512_n215 ), .ZN(_add_512_n207 ) );
NAND2_X2 _add_512_U363  ( .A1(_add_512_n209 ), .A2(_add_512_n210 ), .ZN(_add_512_n208 ) );
NOR2_X4 _add_512_U362  ( .A1(_add_512_n52 ), .A2(_add_512_n184 ), .ZN(_add_512_n180 ) );
INV_X4 _add_512_U361  ( .A(H0[28]), .ZN(_add_512_n182 ) );
INV_X4 _add_512_U360  ( .A(next_A[28]), .ZN(_add_512_n183 ) );
NAND2_X2 _add_512_U359  ( .A1(H0[28]), .A2(next_A[28]), .ZN(_add_512_n159 ));
INV_X4 _add_512_U358  ( .A(_add_512_n159 ), .ZN(_add_512_n174 ) );
XNOR2_X2 _add_512_U357  ( .A(_add_512_n180 ), .B(_add_512_n181 ), .ZN(N880));
NAND2_X2 _add_512_U356  ( .A1(_add_512_n176 ), .A2(_add_512_n136 ), .ZN(_add_512_n172 ) );
XNOR2_X2 _add_512_U355  ( .A(_add_512_n167 ), .B(_add_512_n168 ), .ZN(N881));
INV_X4 _add_512_U354  ( .A(_add_512_n346 ), .ZN(_add_512_n166 ) );
NAND2_X2 _add_512_U353  ( .A1(H0[2]), .A2(next_A[2]), .ZN(_add_512_n118 ) );
NAND2_X2 _add_512_U352  ( .A1(_add_512_n166 ), .A2(_add_512_n118 ), .ZN(_add_512_n164 ) );
NAND2_X2 _add_512_U351  ( .A1(_add_512_n54 ), .A2(_add_512_n425 ), .ZN(_add_512_n120 ) );
XNOR2_X2 _add_512_U350  ( .A(_add_512_n164 ), .B(_add_512_n120 ), .ZN(N854));
NAND2_X2 _add_512_U349  ( .A1(_add_512_n145 ), .A2(_add_512_n142 ), .ZN(_add_512_n162 ) );
NAND2_X2 _add_512_U348  ( .A1(_add_512_n160 ), .A2(_add_512_n136 ), .ZN(_add_512_n152 ) );
NAND2_X2 _add_512_U347  ( .A1(_add_512_n159 ), .A2(_add_512_n158 ), .ZN(_add_512_n156 ) );
NAND2_X2 _add_512_U346  ( .A1(_add_512_n156 ), .A2(_add_512_n157 ), .ZN(_add_512_n134 ) );
INV_X4 _add_512_U345  ( .A(_add_512_n130 ), .ZN(_add_512_n149 ) );
XNOR2_X2 _add_512_U344  ( .A(_add_512_n147 ), .B(_add_512_n148 ), .ZN(N882));
NAND2_X2 _add_512_U343  ( .A1(_add_512_n135 ), .A2(_add_512_n136 ), .ZN(_add_512_n125 ) );
NAND2_X2 _add_512_U342  ( .A1(_add_512_n131 ), .A2(_add_512_n132 ), .ZN(_add_512_n129 ) );
NAND2_X2 _add_512_U341  ( .A1(_add_512_n125 ), .A2(_add_512_n126 ), .ZN(_add_512_n124 ) );
XNOR2_X2 _add_512_U340  ( .A(_add_512_n121 ), .B(_add_512_n122 ), .ZN(N883));
INV_X4 _add_512_U339  ( .A(_add_512_n120 ), .ZN(_add_512_n119 ) );
INV_X4 _add_512_U338  ( .A(_add_512_n118 ), .ZN(_add_512_n117 ) );
XNOR2_X2 _add_512_U337  ( .A(_add_512_n112 ), .B(_add_512_n113 ), .ZN(N855));
INV_X4 _add_512_U336  ( .A(_add_512_n416 ), .ZN(_add_512_n110 ) );
XNOR2_X2 _add_512_U335  ( .A(_add_512_n80 ), .B(_add_512_n111 ), .ZN(N856));
NAND2_X2 _add_512_U334  ( .A1(H0[5]), .A2(next_A[5]), .ZN(_add_512_n94 ) );
INV_X4 _add_512_U333  ( .A(_add_512_n94 ), .ZN(_add_512_n108 ) );
XNOR2_X2 _add_512_U332  ( .A(_add_512_n106 ), .B(_add_512_n107 ), .ZN(N857));
INV_X4 _add_512_U331  ( .A(_add_512_n103 ), .ZN(_add_512_n102 ) );
NAND2_X2 _add_512_U330  ( .A1(_add_512_n95 ), .A2(_add_512_n99 ), .ZN(_add_512_n98 ) );
NAND2_X2 _add_512_U329  ( .A1(_add_512_n93 ), .A2(_add_512_n92 ), .ZN(_add_512_n97 ) );
XNOR2_X2 _add_512_U328  ( .A(_add_512_n96 ), .B(_add_512_n97 ), .ZN(N858) );
NAND2_X2 _add_512_U327  ( .A1(_add_512_n96 ), .A2(_add_512_n93 ), .ZN(_add_512_n91 ) );
NAND2_X2 _add_512_U326  ( .A1(_add_512_n91 ), .A2(_add_512_n92 ), .ZN(_add_512_n88 ) );
NAND2_X2 _add_512_U325  ( .A1(_add_512_n90 ), .A2(_add_512_n87 ), .ZN(_add_512_n89 ) );
XNOR2_X2 _add_512_U324  ( .A(_add_512_n88 ), .B(_add_512_n89 ), .ZN(N859) );
INV_X4 _add_512_U323  ( .A(_add_512_n84 ), .ZN(_add_512_n75 ) );
XNOR2_X2 _add_512_U322  ( .A(_add_512_n82 ), .B(_add_512_n83 ), .ZN(N860) );
INV_X4 _add_512_U321  ( .A(_add_512_n74 ), .ZN(_add_512_n72 ) );
XNOR2_X2 _add_512_U320  ( .A(_add_512_n70 ), .B(_add_512_n71 ), .ZN(N861) );
INV_X8 _add_512_U319  ( .A(_add_512_n353 ), .ZN(_add_512_n332 ) );
NOR3_X1 _add_512_U318  ( .A1(_add_512_n332 ), .A2(_add_512_n61 ), .A3(_add_512_n363 ), .ZN(_add_512_n377 ) );
NOR2_X1 _add_512_U317  ( .A1(_add_512_n380 ), .A2(_add_512_n332 ), .ZN(_add_512_n379 ) );
NAND2_X4 _add_512_U316  ( .A1(_add_512_n372 ), .A2(_add_512_n371 ), .ZN(_add_512_n349 ) );
NAND2_X4 _add_512_U315  ( .A1(_add_512_n286 ), .A2(_add_512_n255 ), .ZN(_add_512_n264 ) );
NAND3_X2 _add_512_U314  ( .A1(_add_512_n350 ), .A2(_add_512_n351 ), .A3(_add_512_n352 ), .ZN(_add_512_n348 ) );
NAND2_X4 _add_512_U313  ( .A1(_add_512_n382 ), .A2(_add_512_n381 ), .ZN(_add_512_n353 ) );
NAND2_X4 _add_512_U312  ( .A1(_add_512_n248 ), .A2(_add_512_n247 ), .ZN(_add_512_n246 ) );
NAND3_X2 _add_512_U311  ( .A1(_add_512_n218 ), .A2(_add_512_n219 ), .A3(_add_512_n191 ), .ZN(_add_512_n142 ) );
NOR2_X2 _add_512_U310  ( .A1(_add_512_n138 ), .A2(_add_512_n137 ), .ZN(_add_512_n160 ) );
NOR3_X2 _add_512_U309  ( .A1(_add_512_n137 ), .A2(_add_512_n1 ), .A3(_add_512_n138 ), .ZN(_add_512_n135 ) );
NOR2_X2 _add_512_U308  ( .A1(_add_512_n25 ), .A2(_add_512_n169 ), .ZN(_add_512_n168 ) );
INV_X4 _add_512_U307  ( .A(_add_512_n69 ), .ZN(_add_512_n236 ) );
NOR2_X4 _add_512_U306  ( .A1(next_A[25]), .A2(H0[25]), .ZN(_add_512_n69 ) );
NOR2_X2 _add_512_U305  ( .A1(_add_512_n137 ), .A2(_add_512_n133 ), .ZN(_add_512_n155 ) );
INV_X1 _add_512_U304  ( .A(_add_512_n236 ), .ZN(_add_512_n67 ) );
NOR3_X2 _add_512_U303  ( .A1(_add_512_n285 ), .A2(_add_512_n9 ), .A3(_add_512_n287 ), .ZN(_add_512_n292 ) );
NOR2_X1 _add_512_U302  ( .A1(_add_512_n9 ), .A2(_add_512_n258 ), .ZN(_add_512_n298 ) );
NAND3_X2 _add_512_U301  ( .A1(_add_512_n33 ), .A2(_add_512_n361 ), .A3(_add_512_n362 ), .ZN(_add_512_n360 ) );
NOR2_X1 _add_512_U300  ( .A1(_add_512_n4 ), .A2(_add_512_n229 ), .ZN(_add_512_n223 ) );
NAND2_X1 _add_512_U299  ( .A1(H0[30]), .A2(next_A[30]), .ZN(_add_512_n130 ));
NOR2_X2 _add_512_U298  ( .A1(_add_512_n194 ), .A2(_add_512_n193 ), .ZN(_add_512_n187 ) );
NAND2_X4 _add_512_U297  ( .A1(_add_512_n276 ), .A2(_add_512_n277 ), .ZN(_add_512_n256 ) );
INV_X2 _add_512_U296  ( .A(_add_512_n205 ), .ZN(_add_512_n365 ) );
NAND2_X4 _add_512_U295  ( .A1(_add_512_n216 ), .A2(_add_512_n177 ), .ZN(_add_512_n146 ) );
NAND2_X2 _add_512_U294  ( .A1(_add_512_n270 ), .A2(_add_512_n271 ), .ZN(_add_512_n268 ) );
NAND2_X2 _add_512_U293  ( .A1(_add_512_n100 ), .A2(_add_512_n101 ), .ZN(_add_512_n421 ) );
XOR2_X2 _add_512_U292  ( .A(next_A[31]), .B(H0[31]), .Z(_add_512_n122 ) );
AND2_X2 _add_512_U291  ( .A1(H0[19]), .A2(_add_512_n39 ), .ZN(_add_512_n65 ));
AND2_X2 _add_512_U290  ( .A1(H0[10]), .A2(_add_512_n35 ), .ZN(_add_512_n64 ));
OR2_X2 _add_512_U289  ( .A1(next_A[0]), .A2(H0[0]), .ZN(_add_512_n63 ) );
NAND3_X2 _add_512_U288  ( .A1(_add_512_n246 ), .A2(H0[23]), .A3(next_A[23]),.ZN(_add_512_n237 ) );
NOR2_X2 _add_512_U287  ( .A1(_add_512_n114 ), .A2(_add_512_n103 ), .ZN(_add_512_n345 ) );
NAND3_X2 _add_512_U286  ( .A1(next_A[1]), .A2(H0[1]), .A3(_add_512_n166 ),.ZN(_add_512_n344 ) );
NAND3_X2 _add_512_U285  ( .A1(_add_512_n343 ), .A2(_add_512_n344 ), .A3(_add_512_n345 ), .ZN(_add_512_n215 ) );
NAND3_X1 _add_512_U284  ( .A1(next_A[5]), .A2(H0[5]), .A3(_add_512_n93 ),.ZN(_add_512_n359 ) );
AND2_X2 _add_512_U283  ( .A1(_add_512_n359 ), .A2(_add_512_n90 ), .ZN(_add_512_n357 ) );
AND2_X2 _add_512_U282  ( .A1(H0[12]), .A2(next_A[12]), .ZN(_add_512_n62 ) );
NOR2_X2 _add_512_U281  ( .A1(next_A[2]), .A2(H0[2]), .ZN(_add_512_n346 ) );
NOR2_X2 _add_512_U280  ( .A1(_add_512_n115 ), .A2(_add_512_n426 ), .ZN(_add_512_n103 ) );
NOR2_X4 _add_512_U279  ( .A1(H0[12]), .A2(next_A[12]), .ZN(_add_512_n61 ) );
NOR2_X2 _add_512_U278  ( .A1(next_A[1]), .A2(H0[1]), .ZN(_add_512_n165 ) );
NOR2_X2 _add_512_U277  ( .A1(next_A[4]), .A2(H0[4]), .ZN(_add_512_n104 ) );
OR2_X2 _add_512_U276  ( .A1(next_A[7]), .A2(H0[7]), .ZN(_add_512_n87 ) );
INV_X8 _add_512_U275  ( .A(_add_512_n349 ), .ZN(_add_512_n335 ) );
INV_X4 _add_512_U274  ( .A(_add_512_n255 ), .ZN(_add_512_n283 ) );
INV_X4 _add_512_U273  ( .A(_add_512_n283 ), .ZN(_add_512_n66 ) );
NAND3_X2 _add_512_U272  ( .A1(_add_512_n214 ), .A2(_add_512_n341 ), .A3(_add_512_n215 ), .ZN(_add_512_n271 ) );
NOR2_X2 _add_512_U271  ( .A1(_add_512_n383 ), .A2(_add_512_n384 ), .ZN(_add_512_n378 ) );
NOR2_X1 _add_512_U270  ( .A1(_add_512_n163 ), .A2(_add_512_n174 ), .ZN(_add_512_n181 ) );
NOR2_X1 _add_512_U269  ( .A1(_add_512_n254 ), .A2(_add_512_n275 ), .ZN(_add_512_n274 ) );
NOR2_X2 _add_512_U268  ( .A1(_add_512_n115 ), .A2(_add_512_n346 ), .ZN(_add_512_n423 ) );
NAND3_X2 _add_512_U267  ( .A1(_add_512_n347 ), .A2(_add_512_n422 ), .A3(_add_512_n423 ), .ZN(_add_512_n101 ) );
AND2_X2 _add_512_U266  ( .A1(_add_512_n86 ), .A2(_add_512_n87 ), .ZN(_add_512_n58 ) );
NOR2_X1 _add_512_U265  ( .A1(_add_512_n283 ), .A2(_add_512_n43 ), .ZN(_add_512_n289 ) );
NOR2_X2 _add_512_U264  ( .A1(_add_512_n61 ), .A2(_add_512_n391 ), .ZN(_add_512_n390 ) );
NOR2_X2 _add_512_U263  ( .A1(_add_512_n62 ), .A2(_add_512_n390 ), .ZN(_add_512_n388 ) );
NOR2_X1 _add_512_U262  ( .A1(_add_512_n384 ), .A2(_add_512_n16 ), .ZN(_add_512_n389 ) );
NAND3_X2 _add_512_U261  ( .A1(_add_512_n62 ), .A2(_add_512_n338 ), .A3(_add_512_n339 ), .ZN(_add_512_n201 ) );
NOR2_X1 _add_512_U260  ( .A1(_add_512_n80 ), .A2(_add_512_n81 ), .ZN(_add_512_n79 ) );
NOR2_X2 _add_512_U259  ( .A1(_add_512_n79 ), .A2(_add_512_n58 ), .ZN(_add_512_n77 ) );
NOR2_X1 _add_512_U258  ( .A1(_add_512_n77 ), .A2(_add_512_n78 ), .ZN(_add_512_n76 ) );
NOR2_X2 _add_512_U257  ( .A1(_add_512_n346 ), .A2(_add_512_n119 ), .ZN(_add_512_n116 ) );
NAND3_X2 _add_512_U256  ( .A1(_add_512_n357 ), .A2(_add_512_n92 ), .A3(_add_512_n358 ), .ZN(_add_512_n356 ) );
NOR2_X2 _add_512_U255  ( .A1(_add_512_n387 ), .A2(_add_512_n57 ), .ZN(_add_512_n56 ) );
NOR2_X1 _add_512_U254  ( .A1(_add_512_n104 ), .A2(_add_512_n105 ), .ZN(_add_512_n95 ) );
NOR2_X2 _add_512_U253  ( .A1(_add_512_n174 ), .A2(_add_512_n175 ), .ZN(_add_512_n173 ) );
NOR2_X1 _add_512_U252  ( .A1(_add_512_n258 ), .A2(_add_512_n257 ), .ZN(_add_512_n284 ) );
NOR2_X2 _add_512_U251  ( .A1(_add_512_n284 ), .A2(_add_512_n283 ), .ZN(_add_512_n282 ) );
NAND3_X2 _add_512_U250  ( .A1(_add_512_n11 ), .A2(_add_512_n401 ), .A3(_add_512_n402 ), .ZN(_add_512_n211 ) );
NOR2_X1 _add_512_U249  ( .A1(_add_512_n337 ), .A2(_add_512_n105 ), .ZN(_add_512_n414 ) );
NAND3_X2 _add_512_U248  ( .A1(_add_512_n90 ), .A2(_add_512_n92 ), .A3(_add_512_n413 ), .ZN(_add_512_n86 ) );
NOR3_X1 _add_512_U247  ( .A1(_add_512_n80 ), .A2(_add_512_n417 ), .A3(_add_512_n81 ), .ZN(_add_512_n409 ) );
NAND3_X2 _add_512_U246  ( .A1(_add_512_n12 ), .A2(_add_512_n74 ), .A3(_add_512_n411 ), .ZN(_add_512_n410 ) );
NOR2_X2 _add_512_U245  ( .A1(_add_512_n409 ), .A2(_add_512_n410 ), .ZN(_add_512_n407 ) );
NOR2_X1 _add_512_U244  ( .A1(_add_512_n65 ), .A2(_add_512_n287 ), .ZN(_add_512_n302 ) );
NOR2_X1 _add_512_U243  ( .A1(_add_512_n252 ), .A2(_add_512_n240 ), .ZN(_add_512_n251 ) );
NOR2_X2 _add_512_U242  ( .A1(_add_512_n67 ), .A2(_add_512_n244 ), .ZN(_add_512_n243 ) );
NOR2_X2 _add_512_U241  ( .A1(_add_512_n75 ), .A2(_add_512_n76 ), .ZN(_add_512_n70 ) );
NOR2_X1 _add_512_U240  ( .A1(_add_512_n72 ), .A2(_add_512_n73 ), .ZN(_add_512_n71 ) );
NOR2_X1 _add_512_U239  ( .A1(_add_512_n80 ), .A2(_add_512_n81 ), .ZN(_add_512_n85 ) );
NOR2_X2 _add_512_U238  ( .A1(_add_512_n85 ), .A2(_add_512_n58 ), .ZN(_add_512_n82 ) );
NOR2_X1 _add_512_U237  ( .A1(_add_512_n78 ), .A2(_add_512_n75 ), .ZN(_add_512_n83 ) );
NOR2_X2 _add_512_U236  ( .A1(_add_512_n406 ), .A2(_add_512_n64 ), .ZN(_add_512_n403 ) );
NOR2_X1 _add_512_U235  ( .A1(_add_512_n80 ), .A2(_add_512_n104 ), .ZN(_add_512_n109 ) );
NOR2_X1 _add_512_U234  ( .A1(_add_512_n108 ), .A2(_add_512_n105 ), .ZN(_add_512_n107 ) );
NOR2_X2 _add_512_U233  ( .A1(_add_512_n109 ), .A2(_add_512_n110 ), .ZN(_add_512_n106 ) );
NOR2_X2 _add_512_U232  ( .A1(_add_512_n301 ), .A2(_add_512_n165 ), .ZN(_add_512_n300 ) );
NOR2_X2 _add_512_U231  ( .A1(_add_512_n116 ), .A2(_add_512_n117 ), .ZN(_add_512_n112 ) );
NOR2_X1 _add_512_U230  ( .A1(_add_512_n78 ), .A2(_add_512_n73 ), .ZN(_add_512_n412 ) );
OR2_X2 _add_512_U229  ( .A1(_add_512_n165 ), .A2(_add_512_n424 ), .ZN(_add_512_n54 ) );
NOR3_X2 _add_512_U228  ( .A1(_add_512_n387 ), .A2(_add_512_n393 ), .A3(_add_512_n386 ), .ZN(_add_512_n391 ) );
NOR2_X2 _add_512_U227  ( .A1(_add_512_n103 ), .A2(_add_512_n421 ), .ZN(_add_512_n80 ) );
AND4_X2 _add_512_U226  ( .A1(_add_512_n179 ), .A2(_add_512_n186 ), .A3(_add_512_n145 ), .A4(_add_512_n142 ), .ZN(_add_512_n52 ) );
AND2_X2 _add_512_U225  ( .A1(_add_512_n385 ), .A2(_add_512_n213 ), .ZN(_add_512_n209 ) );
NOR2_X1 _add_512_U224  ( .A1(_add_512_n163 ), .A2(_add_512_n138 ), .ZN(_add_512_n176 ) );
NOR2_X2 _add_512_U223  ( .A1(_add_512_n198 ), .A2(_add_512_n199 ), .ZN(_add_512_n197 ) );
NAND3_X2 _add_512_U222  ( .A1(_add_512_n196 ), .A2(_add_512_n195 ), .A3(_add_512_n197 ), .ZN(_add_512_n179 ) );
INV_X4 _add_512_U221  ( .A(next_A[17]), .ZN(_add_512_n326 ) );
OR2_X4 _add_512_U220  ( .A1(H0[6]), .A2(next_A[6]), .ZN(_add_512_n93 ) );
AND3_X4 _add_512_U219  ( .A1(_add_512_n101 ), .A2(_add_512_n102 ), .A3(_add_512_n100 ), .ZN(_add_512_n59 ) );
NOR2_X1 _add_512_U218  ( .A1(_add_512_n163 ), .A2(_add_512_n133 ), .ZN(_add_512_n175 ) );
NAND3_X1 _add_512_U217  ( .A1(_add_512_n412 ), .A2(_add_512_n87 ), .A3(_add_512_n86 ), .ZN(_add_512_n411 ) );
INV_X1 _add_512_U216  ( .A(_add_512_n351 ), .ZN(_add_512_n380 ) );
NOR2_X1 _add_512_U215  ( .A1(_add_512_n114 ), .A2(_add_512_n115 ), .ZN(_add_512_n113 ) );
INV_X2 _add_512_U214  ( .A(_add_512_n249 ), .ZN(_add_512_n252 ) );
NOR2_X1 _add_512_U213  ( .A1(_add_512_n64 ), .A2(_add_512_n334 ), .ZN(_add_512_n408 ) );
NOR2_X1 _add_512_U212  ( .A1(_add_512_n104 ), .A2(_add_512_n110 ), .ZN(_add_512_n111 ) );
NOR2_X1 _add_512_U211  ( .A1(_add_512_n62 ), .A2(_add_512_n61 ), .ZN(_add_512_n392 ) );
NAND3_X4 _add_512_U210  ( .A1(_add_512_n418 ), .A2(_add_512_n419 ), .A3(_add_512_n420 ), .ZN(_add_512_n81 ) );
NAND2_X1 _add_512_U209  ( .A1(_add_512_n186 ), .A2(_add_512_n132 ), .ZN(_add_512_n161 ) );
NOR2_X1 _add_512_U208  ( .A1(_add_512_n334 ), .A2(_add_512_n407 ), .ZN(_add_512_n406 ) );
NOR2_X2 _add_512_U207  ( .A1(_add_512_n204 ), .A2(_add_512_n310 ), .ZN(_add_512_n195 ) );
NOR3_X1 _add_512_U206  ( .A1(_add_512_n80 ), .A2(_add_512_n15 ), .A3(_add_512_n81 ), .ZN(_add_512_n387 ) );
NOR3_X4 _add_512_U205  ( .A1(_add_512_n140 ), .A2(_add_512_n139 ), .A3(_add_512_n141 ), .ZN(_add_512_n123 ) );
NOR2_X4 _add_512_U204  ( .A1(_add_512_n337 ), .A2(_add_512_n336 ), .ZN(_add_512_n420 ) );
NAND3_X2 _add_512_U203  ( .A1(_add_512_n366 ), .A2(_add_512_n367 ), .A3(_add_512_n33 ), .ZN(_add_512_n206 ) );
OR3_X2 _add_512_U202  ( .A1(_add_512_n393 ), .A2(_add_512_n62 ), .A3(_add_512_n386 ), .ZN(_add_512_n57 ) );
NOR3_X2 _add_512_U201  ( .A1(_add_512_n194 ), .A2(_add_512_n202 ), .A3(_add_512_n189 ), .ZN(_add_512_n196 ) );
NOR2_X4 _add_512_U200  ( .A1(next_A[11]), .A2(H0[11]), .ZN(_add_512_n333 ));
INV_X4 _add_512_U199  ( .A(_add_512_n36 ), .ZN(_add_512_n138 ) );
NOR2_X4 _add_512_U198  ( .A1(next_A[13]), .A2(H0[13]), .ZN(_add_512_n363 ));
NAND2_X1 _add_512_U197  ( .A1(H0[10]), .A2(_add_512_n35 ), .ZN(_add_512_n399 ) );
NOR2_X4 _add_512_U196  ( .A1(_add_512_n25 ), .A2(_add_512_n163 ), .ZN(_add_512_n132 ) );
INV_X8 _add_512_U195  ( .A(_add_512_n132 ), .ZN(_add_512_n137 ) );
NAND2_X4 _add_512_U194  ( .A1(_add_512_n314 ), .A2(_add_512_n313 ), .ZN(_add_512_n266 ) );
NOR3_X2 _add_512_U193  ( .A1(_add_512_n334 ), .A2(_add_512_n84 ), .A3(_add_512_n73 ), .ZN(_add_512_n397 ) );
NAND2_X4 _add_512_U192  ( .A1(_add_512_n224 ), .A2(_add_512_n225 ), .ZN(_add_512_n136 ) );
INV_X2 _add_512_U191  ( .A(_add_512_n15 ), .ZN(_add_512_n210 ) );
NOR2_X4 _add_512_U190  ( .A1(_add_512_n124 ), .A2(_add_512_n123 ), .ZN(_add_512_n121 ) );
INV_X1 _add_512_U189  ( .A(_add_512_n65 ), .ZN(_add_512_n46 ) );
AND2_X2 _add_512_U188  ( .A1(_add_512_n46 ), .A2(_add_512_n287 ), .ZN(_add_512_n45 ) );
INV_X8 _add_512_U187  ( .A(_add_512_n219 ), .ZN(_add_512_n194 ) );
NAND2_X4 _add_512_U186  ( .A1(_add_512_n232 ), .A2(_add_512_n231 ), .ZN(_add_512_n226 ) );
NAND2_X4 _add_512_U185  ( .A1(_add_512_n234 ), .A2(_add_512_n30 ), .ZN(_add_512_n224 ) );
NAND2_X4 _add_512_U184  ( .A1(_add_512_n230 ), .A2(_add_512_n226 ), .ZN(_add_512_n217 ) );
NAND2_X4 _add_512_U183  ( .A1(_add_512_n183 ), .A2(_add_512_n182 ), .ZN(_add_512_n178 ) );
INV_X8 _add_512_U182  ( .A(_add_512_n178 ), .ZN(_add_512_n163 ) );
NAND2_X1 _add_512_U181  ( .A1(H0[15]), .A2(_add_512_n28 ), .ZN(_add_512_n350 ) );
NAND2_X4 _add_512_U180  ( .A1(_add_512_n321 ), .A2(_add_512_n322 ), .ZN(_add_512_n314 ) );
NAND2_X1 _add_512_U179  ( .A1(_add_512_n27 ), .A2(_add_512_n322 ), .ZN(_add_512_n324 ) );
NAND2_X1 _add_512_U178  ( .A1(_add_512_n280 ), .A2(_add_512_n281 ), .ZN(_add_512_n279 ) );
NAND2_X2 _add_512_U177  ( .A1(_add_512_n185 ), .A2(_add_512_n133 ), .ZN(_add_512_n184 ) );
NOR2_X2 _add_512_U176  ( .A1(_add_512_n285 ), .A2(_add_512_n264 ), .ZN(_add_512_n278 ) );
NOR2_X4 _add_512_U175  ( .A1(_add_512_n292 ), .A2(_add_512_n293 ), .ZN(_add_512_n288 ) );
NAND2_X4 _add_512_U174  ( .A1(_add_512_n326 ), .A2(_add_512_n325 ), .ZN(_add_512_n68 ) );
NOR2_X4 _add_512_U173  ( .A1(_add_512_n150 ), .A2(_add_512_n151 ), .ZN(_add_512_n147 ) );
INV_X2 _add_512_U172  ( .A(_add_512_n272 ), .ZN(_add_512_n308 ) );
NOR2_X4 _add_512_U171  ( .A1(_add_512_n128 ), .A2(_add_512_n127 ), .ZN(_add_512_n126 ) );
NOR2_X1 _add_512_U170  ( .A1(_add_512_n205 ), .A2(_add_512_n333 ), .ZN(_add_512_n393 ) );
NOR3_X2 _add_512_U169  ( .A1(_add_512_n139 ), .A2(_add_512_n161 ), .A3(_add_512_n162 ), .ZN(_add_512_n150 ) );
NAND2_X2 _add_512_U168  ( .A1(_add_512_n129 ), .A2(_add_512_n130 ), .ZN(_add_512_n128 ) );
INV_X2 _add_512_U167  ( .A(_add_512_n41 ), .ZN(_add_512_n42 ) );
INV_X2 _add_512_U166  ( .A(_add_512_n134 ), .ZN(_add_512_n154 ) );
NOR2_X2 _add_512_U165  ( .A1(_add_512_n334 ), .A2(_add_512_n398 ), .ZN(_add_512_n396 ) );
OR2_X2 _add_512_U164  ( .A1(_add_512_n241 ), .A2(_add_512_n240 ), .ZN(_add_512_n55 ) );
NOR2_X4 _add_512_U163  ( .A1(_add_512_n278 ), .A2(_add_512_n279 ), .ZN(_add_512_n273 ) );
NAND2_X1 _add_512_U162  ( .A1(H0[14]), .A2(next_A[14]), .ZN(_add_512_n351 ));
NOR2_X1 _add_512_U161  ( .A1(_add_512_n229 ), .A2(_add_512_n55 ), .ZN(_add_512_n245 ) );
INV_X4 _add_512_U160  ( .A(next_A[14]), .ZN(_add_512_n382 ) );
OR2_X4 _add_512_U159  ( .A1(_add_512_n331 ), .A2(_add_512_n272 ), .ZN(_add_512_n53 ) );
NAND2_X4 _add_512_U158  ( .A1(_add_512_n305 ), .A2(_add_512_n192 ), .ZN(_add_512_n304 ) );
AND2_X2 _add_512_U157  ( .A1(_add_512_n142 ), .A2(_add_512_n21 ), .ZN(_add_512_n40 ) );
NAND2_X2 _add_512_U156  ( .A1(_add_512_n179 ), .A2(_add_512_n40 ), .ZN(_add_512_n49 ) );
NOR2_X2 _add_512_U155  ( .A1(_add_512_n14 ), .A2(_add_512_n133 ), .ZN(_add_512_n131 ) );
INV_X4 _add_512_U154  ( .A(next_A[27]), .ZN(_add_512_n222 ) );
NOR2_X2 _add_512_U153  ( .A1(_add_512_n223 ), .A2(_add_512_n20 ), .ZN(_add_512_n220 ) );
NAND2_X2 _add_512_U152  ( .A1(_add_512_n290 ), .A2(_add_512_n291 ), .ZN(_add_512_n255 ) );
NAND2_X4 _add_512_U151  ( .A1(_add_512_n187 ), .A2(_add_512_n188 ), .ZN(_add_512_n145 ) );
NOR2_X2 _add_512_U150  ( .A1(_add_512_n335 ), .A2(_add_512_n363 ), .ZN(_add_512_n367 ) );
NAND2_X2 _add_512_U149  ( .A1(_add_512_n144 ), .A2(_add_512_n145 ), .ZN(_add_512_n140 ) );
NOR2_X2 _add_512_U148  ( .A1(_add_512_n137 ), .A2(_add_512_n146 ), .ZN(_add_512_n144 ) );
NAND2_X1 _add_512_U147  ( .A1(_add_512_n186 ), .A2(_add_512_n145 ), .ZN(_add_512_n48 ) );
NOR2_X4 _add_512_U146  ( .A1(_add_512_n206 ), .A2(_add_512_n205 ), .ZN(_add_512_n310 ) );
NAND2_X1 _add_512_U145  ( .A1(_add_512_n142 ), .A2(_add_512_n143 ), .ZN(_add_512_n141 ) );
INV_X1 _add_512_U144  ( .A(_add_512_n350 ), .ZN(_add_512_n370 ) );
NOR2_X2 _add_512_U143  ( .A1(_add_512_n267 ), .A2(_add_512_n272 ), .ZN(_add_512_n270 ) );
INV_X4 _add_512_U142  ( .A(_add_512_n201 ), .ZN(_add_512_n272 ) );
NAND2_X1 _add_512_U141  ( .A1(_add_512_n200 ), .A2(_add_512_n201 ), .ZN(_add_512_n198 ) );
INV_X4 _add_512_U140  ( .A(_add_512_n43 ), .ZN(_add_512_n281 ) );
NOR2_X2 _add_512_U139  ( .A1(_add_512_n291 ), .A2(_add_512_n290 ), .ZN(_add_512_n43 ) );
NAND3_X4 _add_512_U138  ( .A1(_add_512_n294 ), .A2(_add_512_n38 ), .A3(_add_512_n281 ), .ZN(_add_512_n37 ) );
NAND2_X4 _add_512_U137  ( .A1(next_A[22]), .A2(H0[22]), .ZN(_add_512_n191 ));
NOR2_X4 _add_512_U136  ( .A1(_add_512_n170 ), .A2(_add_512_n171 ), .ZN(_add_512_n167 ) );
NAND2_X4 _add_512_U135  ( .A1(_add_512_n235 ), .A2(_add_512_n236 ), .ZN(_add_512_n227 ) );
NAND2_X2 _add_512_U134  ( .A1(_add_512_n222 ), .A2(_add_512_n221 ), .ZN(_add_512_n177 ) );
NAND2_X4 _add_512_U133  ( .A1(_add_512_n221 ), .A2(_add_512_n222 ), .ZN(_add_512_n36 ) );
NAND2_X4 _add_512_U132  ( .A1(_add_512_n312 ), .A2(_add_512_n313 ), .ZN(_add_512_n311 ) );
INV_X8 _add_512_U131  ( .A(_add_512_n311 ), .ZN(_add_512_n193 ) );
INV_X2 _add_512_U130  ( .A(_add_512_n377 ), .ZN(_add_512_n376 ) );
INV_X1 _add_512_U129  ( .A(_add_512_n363 ), .ZN(_add_512_n338 ) );
NOR2_X4 _add_512_U128  ( .A1(_add_512_n363 ), .A2(_add_512_n61 ), .ZN(_add_512_n385 ) );
INV_X8 _add_512_U127  ( .A(_add_512_n266 ), .ZN(_add_512_n189 ) );
INV_X2 _add_512_U126  ( .A(_add_512_n34 ), .ZN(_add_512_n35 ) );
INV_X1 _add_512_U125  ( .A(next_A[13]), .ZN(_add_512_n41 ) );
OR2_X2 _add_512_U124  ( .A1(_add_512_n303 ), .A2(_add_512_n65 ), .ZN(_add_512_n47 ) );
INV_X4 _add_512_U123  ( .A(_add_512_n258 ), .ZN(_add_512_n38 ) );
NAND2_X1 _add_512_U122  ( .A1(next_A[9]), .A2(H0[9]), .ZN(_add_512_n398 ) );
INV_X8 _add_512_U121  ( .A(_add_512_n203 ), .ZN(_add_512_n202 ) );
INV_X4 _add_512_U120  ( .A(_add_512_n202 ), .ZN(_add_512_n31 ) );
NOR2_X1 _add_512_U119  ( .A1(_add_512_n335 ), .A2(_add_512_n370 ), .ZN(_add_512_n369 ) );
INV_X2 _add_512_U118  ( .A(_add_512_n206 ), .ZN(_add_512_n364 ) );
INV_X4 _add_512_U117  ( .A(_add_512_n29 ), .ZN(_add_512_n30 ) );
INV_X2 _add_512_U116  ( .A(_add_512_n226 ), .ZN(_add_512_n29 ) );
INV_X1 _add_512_U115  ( .A(_add_512_n372 ), .ZN(_add_512_n28 ) );
NAND2_X2 _add_512_U114  ( .A1(H0[17]), .A2(next_A[17]), .ZN(_add_512_n322 ));
INV_X1 _add_512_U113  ( .A(_add_512_n230 ), .ZN(_add_512_n239 ) );
INV_X1 _add_512_U112  ( .A(_add_512_n228 ), .ZN(_add_512_n244 ) );
INV_X1 _add_512_U111  ( .A(_add_512_n319 ), .ZN(_add_512_n27 ) );
XNOR2_X1 _add_512_U110  ( .A(_add_512_n285 ), .B(_add_512_n302 ), .ZN(N871));
INV_X1 _add_512_U109  ( .A(_add_512_n314 ), .ZN(_add_512_n317 ) );
INV_X4 _add_512_U108  ( .A(_add_512_n25 ), .ZN(_add_512_n157 ) );
INV_X1 _add_512_U107  ( .A(_add_512_n335 ), .ZN(_add_512_n24 ) );
NOR2_X4 _add_512_U106  ( .A1(_add_512_n155 ), .A2(_add_512_n154 ), .ZN(_add_512_n153 ) );
INV_X2 _add_512_U105  ( .A(_add_512_n22 ), .ZN(_add_512_n23 ) );
INV_X1 _add_512_U104  ( .A(_add_512_n312 ), .ZN(_add_512_n22 ) );
NAND2_X1 _add_512_U103  ( .A1(H0[23]), .A2(next_A[23]), .ZN(_add_512_n249 ));
INV_X1 _add_512_U102  ( .A(_add_512_n163 ), .ZN(_add_512_n21 ) );
INV_X2 _add_512_U101  ( .A(_add_512_n19 ), .ZN(_add_512_n20 ) );
INV_X1 _add_512_U100  ( .A(_add_512_n136 ), .ZN(_add_512_n19 ) );
NAND2_X4 _add_512_U99  ( .A1(_add_512_n262 ), .A2(_add_512_n261 ), .ZN(_add_512_n260 ) );
AND2_X2 _add_512_U98  ( .A1(_add_512_n238 ), .A2(_add_512_n3 ), .ZN(_add_512_n18 ) );
XNOR2_X2 _add_512_U97  ( .A(_add_512_n17 ), .B(_add_512_n18 ), .ZN(N876) );
AND3_X4 _add_512_U96  ( .A1(_add_512_n385 ), .A2(_add_512_n11 ), .A3(_add_512_n401 ), .ZN(_add_512_n354 ) );
NAND2_X1 _add_512_U95  ( .A1(_add_512_n192 ), .A2(_add_512_n191 ), .ZN(_add_512_n199 ) );
NAND2_X1 _add_512_U94  ( .A1(_add_512_n191 ), .A2(_add_512_n192 ), .ZN(_add_512_n190 ) );
NOR2_X4 _add_512_U93  ( .A1(_add_512_n207 ), .A2(_add_512_n208 ), .ZN(_add_512_n204 ) );
NOR2_X1 _add_512_U92  ( .A1(_add_512_n229 ), .A2(_add_512_n240 ), .ZN(_add_512_n250 ) );
NOR2_X2 _add_512_U91  ( .A1(_add_512_n189 ), .A2(_add_512_n190 ), .ZN(_add_512_n188 ) );
INV_X1 _add_512_U90  ( .A(_add_512_n338 ), .ZN(_add_512_n16 ) );
NAND2_X4 _add_512_U89  ( .A1(_add_512_n348 ), .A2(_add_512_n24 ), .ZN(_add_512_n203 ) );
NOR3_X2 _add_512_U88  ( .A1(_add_512_n394 ), .A2(_add_512_n336 ), .A3(_add_512_n211 ), .ZN(_add_512_n386 ) );
NOR2_X4 _add_512_U87  ( .A1(_add_512_n211 ), .A2(_add_512_n342 ), .ZN(_add_512_n341 ) );
NAND2_X4 _add_512_U86  ( .A1(_add_512_n153 ), .A2(_add_512_n152 ), .ZN(_add_512_n151 ) );
NAND3_X2 _add_512_U85  ( .A1(_add_512_n11 ), .A2(_add_512_n401 ), .A3(_add_512_n402 ), .ZN(_add_512_n15 ) );
INV_X2 _add_512_U84  ( .A(next_A[18]), .ZN(_add_512_n316 ) );
NAND2_X4 _add_512_U83  ( .A1(_add_512_n315 ), .A2(_add_512_n316 ), .ZN(_add_512_n313 ) );
INV_X4 _add_512_U82  ( .A(next_A[22]), .ZN(_add_512_n277 ) );
INV_X8 _add_512_U81  ( .A(_add_512_n146 ), .ZN(_add_512_n186 ) );
INV_X4 _add_512_U80  ( .A(_add_512_n179 ), .ZN(_add_512_n139 ) );
NAND2_X4 _add_512_U79  ( .A1(_add_512_n263 ), .A2(_add_512_n256 ), .ZN(_add_512_n218 ) );
NOR2_X2 _add_512_U78  ( .A1(_add_512_n134 ), .A2(_add_512_n1 ), .ZN(_add_512_n127 ) );
INV_X4 _add_512_U77  ( .A(_add_512_n14 ), .ZN(_add_512_n143 ) );
NOR2_X4 _add_512_U76  ( .A1(next_A[30]), .A2(H0[30]), .ZN(_add_512_n14 ) );
NOR2_X2 _add_512_U75  ( .A1(_add_512_n304 ), .A2(_add_512_n47 ), .ZN(_add_512_n44 ) );
OR2_X2 _add_512_U74  ( .A1(_add_512_n44 ), .A2(_add_512_n45 ), .ZN(_add_512_n297 ) );
NAND2_X2 _add_512_U73  ( .A1(_add_512_n136 ), .A2(_add_512_n36 ), .ZN(_add_512_n185 ) );
NAND2_X2 _add_512_U72  ( .A1(_add_512_n306 ), .A2(_add_512_n193 ), .ZN(_add_512_n305 ) );
XNOR2_X2 _add_512_U71  ( .A(_add_512_n26 ), .B(_add_512_n251 ), .ZN(N875) );
INV_X2 _add_512_U70  ( .A(_add_512_n200 ), .ZN(_add_512_n309 ) );
NOR2_X2 _add_512_U69  ( .A1(_add_512_n310 ), .A2(_add_512_n309 ), .ZN(_add_512_n307 ) );
OR2_X2 _add_512_U68  ( .A1(_add_512_n332 ), .A2(_add_512_n375 ), .ZN(_add_512_n60 ) );
NOR2_X2 _add_512_U67  ( .A1(_add_512_n335 ), .A2(_add_512_n332 ), .ZN(_add_512_n339 ) );
NOR2_X1 _add_512_U66  ( .A1(_add_512_n56 ), .A2(_add_512_n212 ), .ZN(_add_512_n383 ) );
NOR2_X2 _add_512_U65  ( .A1(_add_512_n56 ), .A2(_add_512_n376 ), .ZN(_add_512_n373 ) );
NOR2_X4 _add_512_U64  ( .A1(_add_512_n373 ), .A2(_add_512_n374 ), .ZN(_add_512_n368 ) );
NAND2_X4 _add_512_U63  ( .A1(_add_512_n328 ), .A2(_add_512_n327 ), .ZN(_add_512_n323 ) );
BUF_X8 _add_512_U62  ( .A(_add_512_n229 ), .Z(_add_512_n26 ) );
AND2_X4 _add_512_U61  ( .A1(_add_512_n424 ), .A2(_add_512_n63 ), .ZN(N852));
INV_X1 _add_512_U60  ( .A(_add_512_n320 ), .ZN(_add_512_n329 ) );
OR2_X4 _add_512_U59  ( .A1(_add_512_n73 ), .A2(_add_512_n84 ), .ZN(_add_512_n12 ) );
INV_X1 _add_512_U58  ( .A(_add_512_n385 ), .ZN(_add_512_n212 ) );
OR2_X2 _add_512_U57  ( .A1(next_A[9]), .A2(H0[9]), .ZN(_add_512_n11 ) );
NAND3_X4 _add_512_U56  ( .A1(_add_512_n68 ), .A2(H0[16]), .A3(n13108), .ZN(_add_512_n321 ) );
NOR2_X4 _add_512_U55  ( .A1(_add_512_n267 ), .A2(_add_512_n193 ), .ZN(_add_512_n265 ) );
NAND2_X4 _add_512_U54  ( .A1(_add_512_n314 ), .A2(_add_512_n313 ), .ZN(_add_512_n32 ) );
NAND2_X4 _add_512_U53  ( .A1(_add_512_n265 ), .A2(_add_512_n32 ), .ZN(_add_512_n261 ) );
BUF_X16 _add_512_U52  ( .A(next_A[19]), .Z(_add_512_n39 ) );
NAND2_X2 _add_512_U51  ( .A1(next_A[27]), .A2(H0[27]), .ZN(_add_512_n133 ));
NAND2_X2 _add_512_U50  ( .A1(next_A[19]), .A2(H0[19]), .ZN(_add_512_n296 ));
NOR2_X2 _add_512_U49  ( .A1(next_A[19]), .A2(H0[19]), .ZN(_add_512_n287 ) );
OR2_X2 _add_512_U48  ( .A1(_add_512_n194 ), .A2(_add_512_n254 ), .ZN(_add_512_n51 ) );
INV_X8 _add_512_U47  ( .A(_add_512_n217 ), .ZN(_add_512_n216 ) );
NOR2_X2 _add_512_U46  ( .A1(_add_512_n1 ), .A2(_add_512_n149 ), .ZN(_add_512_n148 ) );
NAND2_X2 _add_512_U45  ( .A1(_add_512_n172 ), .A2(_add_512_n173 ), .ZN(_add_512_n171 ) );
NOR2_X2 _add_512_U44  ( .A1(_add_512_n287 ), .A2(_add_512_n8 ), .ZN(_add_512_n286 ) );
INV_X4 _add_512_U43  ( .A(_add_512_n332 ), .ZN(_add_512_n33 ) );
NOR2_X4 _add_512_U42  ( .A1(_add_512_n49 ), .A2(_add_512_n48 ), .ZN(_add_512_n170 ) );
INV_X8 _add_512_U41  ( .A(next_A[21]), .ZN(_add_512_n291 ) );
NOR2_X2 _add_512_U40  ( .A1(_add_512_n250 ), .A2(_add_512_n252 ), .ZN(_add_512_n17 ) );
INV_X4 _add_512_U39  ( .A(next_A[10]), .ZN(_add_512_n34 ) );
NOR2_X2 _add_512_U38  ( .A1(_add_512_n245 ), .A2(_add_512_n2 ), .ZN(_add_512_n242 ) );
INV_X4 _add_512_U37  ( .A(_add_512_n257 ), .ZN(_add_512_n294 ) );
AND2_X2 _add_512_U36  ( .A1(_add_512_n133 ), .A2(_add_512_n36 ), .ZN(_add_512_n10 ) );
NAND2_X4 _add_512_U35  ( .A1(_add_512_n227 ), .A2(_add_512_n228 ), .ZN(_add_512_n234 ) );
NAND2_X1 _add_512_U34  ( .A1(_add_512_n59 ), .A2(_add_512_n416 ), .ZN(_add_512_n99 ) );
NOR2_X4 _add_512_U33  ( .A1(next_A[3]), .A2(H0[3]), .ZN(_add_512_n115 ) );
INV_X4 _add_512_U32  ( .A(_add_512_n246 ), .ZN(_add_512_n241 ) );
INV_X4 _add_512_U31  ( .A(_add_512_n32 ), .ZN(_add_512_n303 ) );
NOR2_X4 _add_512_U30  ( .A1(next_A[29]), .A2(H0[29]), .ZN(_add_512_n25 ) );
INV_X1 _add_512_U29  ( .A(_add_512_n299 ), .ZN(_add_512_n9 ) );
NOR2_X4 _add_512_U28  ( .A1(_add_512_n81 ), .A2(_add_512_n115 ), .ZN(_add_512_n214 ) );
NAND2_X1 _add_512_U27  ( .A1(_add_512_n98 ), .A2(_add_512_n94 ), .ZN(_add_512_n96 ) );
INV_X4 _add_512_U26  ( .A(_add_512_n8 ), .ZN(_add_512_n299 ) );
NOR2_X4 _add_512_U25  ( .A1(next_A[20]), .A2(H0[20]), .ZN(_add_512_n8 ) );
NOR2_X1 _add_512_U24  ( .A1(_add_512_n333 ), .A2(_add_512_n405 ), .ZN(_add_512_n404 ) );
NOR2_X1 _add_512_U23  ( .A1(_add_512_n61 ), .A2(_add_512_n333 ), .ZN(_add_512_n366 ) );
AND2_X4 _add_512_U22  ( .A1(_add_512_n225 ), .A2(_add_512_n30 ), .ZN(_add_512_n7 ) );
XNOR2_X2 _add_512_U21  ( .A(_add_512_n50 ), .B(_add_512_n7 ), .ZN(N878) );
AND2_X2 _add_512_U20  ( .A1(_add_512_n313 ), .A2(_add_512_n192 ), .ZN(_add_512_n6 ) );
AND2_X2 _add_512_U19  ( .A1(_add_512_n318 ), .A2(_add_512_n317 ), .ZN(_add_512_n5 ) );
XNOR2_X2 _add_512_U18  ( .A(_add_512_n5 ), .B(_add_512_n6 ), .ZN(N870) );
INV_X1 _add_512_U17  ( .A(_add_512_n216 ), .ZN(_add_512_n4 ) );
NOR2_X2 _add_512_U16  ( .A1(_add_512_n233 ), .A2(_add_512_n234 ), .ZN(_add_512_n50 ) );
NAND2_X1 _add_512_U15  ( .A1(_add_512_n294 ), .A2(_add_512_n295 ), .ZN(_add_512_n293 ) );
INV_X4 _add_512_U14  ( .A(next_A[26]), .ZN(_add_512_n232 ) );
NAND2_X1 _add_512_U13  ( .A1(H0[26]), .A2(next_A[26]), .ZN(_add_512_n225 ));
INV_X2 _add_512_U12  ( .A(_add_512_n241 ), .ZN(_add_512_n3 ) );
OR2_X2 _add_512_U11  ( .A1(_add_512_n247 ), .A2(_add_512_n248 ), .ZN(_add_512_n238 ) );
NAND2_X2 _add_512_U10  ( .A1(_add_512_n237 ), .A2(_add_512_n238 ), .ZN(_add_512_n235 ) );
BUF_X16 _add_512_U9  ( .A(_add_512_n235 ), .Z(_add_512_n2 ) );
NAND2_X4 _add_512_U8  ( .A1(H0[29]), .A2(next_A[29]), .ZN(_add_512_n158 ) );
INV_X4 _add_512_U7  ( .A(_add_512_n158 ), .ZN(_add_512_n169 ) );
NOR2_X1 _add_512_U6  ( .A1(_add_512_n229 ), .A2(_add_512_n239 ), .ZN(_add_512_n233 ) );
INV_X4 _add_512_U5  ( .A(_add_512_n143 ), .ZN(_add_512_n1 ) );
NAND4_X1 _add_512_U4  ( .A1(_add_512_n31 ), .A2(_add_512_n271 ), .A3(_add_512_n340 ), .A4(_add_512_n200 ), .ZN(_add_512_n331 ) );
NAND3_X1 _add_512_U3  ( .A1(_add_512_n42 ), .A2(H0[13]), .A3(_add_512_n353 ),.ZN(_add_512_n352 ) );
NAND2_X1 _add_512_U2  ( .A1(H0[13]), .A2(_add_512_n42 ), .ZN(_add_512_n375 ));
NOR2_X4 _add_0_root_add_136_4_U458  ( .A1(N104), .A2(N136), .ZN(_add_0_root_add_136_4_n100 ) );
NOR2_X4 _add_0_root_add_136_4_U457  ( .A1(N137), .A2(N105), .ZN(_add_0_root_add_136_4_n95 ) );
NAND2_X2 _add_0_root_add_136_4_U456  ( .A1(_add_0_root_add_136_4_n433 ),.A2(_add_0_root_add_136_4_n434 ), .ZN(_add_0_root_add_136_4_n429 ) );
NAND2_X2 _add_0_root_add_136_4_U455  ( .A1(N101), .A2(N133), .ZN(_add_0_root_add_136_4_n432 ) );
NAND2_X2 _add_0_root_add_136_4_U454  ( .A1(_add_0_root_add_136_4_n29 ), .A2(N99), .ZN(_add_0_root_add_136_4_n120 ) );
NAND2_X2 _add_0_root_add_136_4_U453  ( .A1(_add_0_root_add_136_4_n258 ),.A2(_add_0_root_add_136_4_n428 ), .ZN(_add_0_root_add_136_4_n427 ) );
NOR2_X4 _add_0_root_add_136_4_U452  ( .A1(_add_0_root_add_136_4_n133 ), .A2(_add_0_root_add_136_4_n425 ), .ZN(_add_0_root_add_136_4_n121 ) );
INV_X4 _add_0_root_add_136_4_U451  ( .A(_add_0_root_add_136_4_n131 ), .ZN(_add_0_root_add_136_4_n424 ) );
INV_X4 _add_0_root_add_136_4_U450  ( .A(_add_0_root_add_136_4_n119 ), .ZN(_add_0_root_add_136_4_n256 ) );
INV_X4 _add_0_root_add_136_4_U449  ( .A(_add_0_root_add_136_4_n126 ), .ZN(_add_0_root_add_136_4_n103 ) );
INV_X4 _add_0_root_add_136_4_U448  ( .A(_add_0_root_add_136_4_n435 ), .ZN(_add_0_root_add_136_4_n421 ) );
INV_X4 _add_0_root_add_136_4_U447  ( .A(_add_0_root_add_136_4_n125 ), .ZN(_add_0_root_add_136_4_n116 ) );
NOR2_X4 _add_0_root_add_136_4_U446  ( .A1(_add_0_root_add_136_4_n34 ), .A2(_add_0_root_add_136_4_n431 ), .ZN(_add_0_root_add_136_4_n422 ) );
NAND3_X4 _add_0_root_add_136_4_U445  ( .A1(_add_0_root_add_136_4_n422 ),.A2(_add_0_root_add_136_4_n116 ), .A3(_add_0_root_add_136_4_n421 ),.ZN(_add_0_root_add_136_4_n104 ) );
NAND2_X2 _add_0_root_add_136_4_U444  ( .A1(N137), .A2(N105), .ZN(_add_0_root_add_136_4_n96 ) );
NAND2_X2 _add_0_root_add_136_4_U443  ( .A1(N139), .A2(N107), .ZN(_add_0_root_add_136_4_n395 ) );
INV_X4 _add_0_root_add_136_4_U442  ( .A(_add_0_root_add_136_4_n416 ), .ZN(_add_0_root_add_136_4_n415 ) );
NAND2_X2 _add_0_root_add_136_4_U441  ( .A1(_add_0_root_add_136_4_n415 ),.A2(_add_0_root_add_136_4_n96 ), .ZN(_add_0_root_add_136_4_n412 ) );
NAND2_X2 _add_0_root_add_136_4_U440  ( .A1(_add_0_root_add_136_4_n412 ),.A2(_add_0_root_add_136_4_n413 ), .ZN(_add_0_root_add_136_4_n411 ) );
XNOR2_X2 _add_0_root_add_136_4_U439  ( .A(_add_0_root_add_136_4_n406 ), .B(_add_0_root_add_136_4_n407 ), .ZN(_add_0_root_add_136_4_n405 ) );
INV_X4 _add_0_root_add_136_4_U438  ( .A(_add_0_root_add_136_4_n405 ), .ZN(next_A[11]) );
INV_X4 _add_0_root_add_136_4_U437  ( .A(_add_0_root_add_136_4_n100 ), .ZN(_add_0_root_add_136_4_n404 ) );
NOR2_X4 _add_0_root_add_136_4_U436  ( .A1(_add_0_root_add_136_4_n402 ), .A2(_add_0_root_add_136_4_n95 ), .ZN(_add_0_root_add_136_4_n360 ) );
NAND2_X2 _add_0_root_add_136_4_U435  ( .A1(N105), .A2(N137), .ZN(_add_0_root_add_136_4_n398 ) );
NOR2_X4 _add_0_root_add_136_4_U434  ( .A1(_add_0_root_add_136_4_n391 ), .A2(_add_0_root_add_136_4_n390 ), .ZN(_add_0_root_add_136_4_n389 ) );
INV_X4 _add_0_root_add_136_4_U433  ( .A(_add_0_root_add_136_4_n104 ), .ZN(_add_0_root_add_136_4_n370 ) );
NAND2_X2 _add_0_root_add_136_4_U432  ( .A1(N140), .A2(N108), .ZN(_add_0_root_add_136_4_n377 ) );
INV_X4 _add_0_root_add_136_4_U431  ( .A(_add_0_root_add_136_4_n377 ), .ZN(_add_0_root_add_136_4_n175 ) );
INV_X4 _add_0_root_add_136_4_U430  ( .A(_add_0_root_add_136_4_n355 ), .ZN(_add_0_root_add_136_4_n380 ) );
XNOR2_X2 _add_0_root_add_136_4_U429  ( .A(_add_0_root_add_136_4_n383 ), .B(_add_0_root_add_136_4_n384 ), .ZN(next_A[13]) );
NAND2_X2 _add_0_root_add_136_4_U428  ( .A1(N142), .A2(N110), .ZN(_add_0_root_add_136_4_n344 ) );
INV_X4 _add_0_root_add_136_4_U427  ( .A(N142), .ZN(_add_0_root_add_136_4_n381 ) );
INV_X4 _add_0_root_add_136_4_U426  ( .A(N110), .ZN(_add_0_root_add_136_4_n382 ) );
NAND2_X2 _add_0_root_add_136_4_U425  ( .A1(_add_0_root_add_136_4_n378 ),.A2(_add_0_root_add_136_4_n377 ), .ZN(_add_0_root_add_136_4_n375 ) );
INV_X4 _add_0_root_add_136_4_U424  ( .A(_add_0_root_add_136_4_n376 ), .ZN(_add_0_root_add_136_4_n356 ) );
NAND2_X2 _add_0_root_add_136_4_U423  ( .A1(N144), .A2(N112), .ZN(_add_0_root_add_136_4_n337 ) );
INV_X4 _add_0_root_add_136_4_U422  ( .A(_add_0_root_add_136_4_n346 ), .ZN(_add_0_root_add_136_4_n358 ) );
NAND2_X2 _add_0_root_add_136_4_U421  ( .A1(_add_0_root_add_136_4_n182 ),.A2(_add_0_root_add_136_4_n120 ), .ZN(_add_0_root_add_136_4_n354 ) );
NAND2_X2 _add_0_root_add_136_4_U420  ( .A1(_add_0_root_add_136_4_n258 ),.A2(_add_0_root_add_136_4_n428 ), .ZN(_add_0_root_add_136_4_n353 ) );
INV_X4 _add_0_root_add_136_4_U419  ( .A(_add_0_root_add_136_4_n120 ), .ZN(_add_0_root_add_136_4_n130 ) );
NAND2_X2 _add_0_root_add_136_4_U418  ( .A1(_add_0_root_add_136_4_n12 ), .A2(_add_0_root_add_136_4_n351 ), .ZN(_add_0_root_add_136_4_n348 ) );
NAND3_X4 _add_0_root_add_136_4_U417  ( .A1(_add_0_root_add_136_4_n347 ),.A2(_add_0_root_add_136_4_n108 ), .A3(_add_0_root_add_136_4_n72 ),.ZN(_add_0_root_add_136_4_n234 ) );
INV_X4 _add_0_root_add_136_4_U416  ( .A(_add_0_root_add_136_4_n330 ), .ZN(_add_0_root_add_136_4_n321 ) );
INV_X4 _add_0_root_add_136_4_U415  ( .A(_add_0_root_add_136_4_n318 ), .ZN(_add_0_root_add_136_4_n339 ) );
NAND2_X2 _add_0_root_add_136_4_U414  ( .A1(_add_0_root_add_136_4_n54 ), .A2(N113), .ZN(_add_0_root_add_136_4_n315 ) );
INV_X4 _add_0_root_add_136_4_U413  ( .A(N145), .ZN(_add_0_root_add_136_4_n335 ) );
INV_X4 _add_0_root_add_136_4_U412  ( .A(N113), .ZN(_add_0_root_add_136_4_n336 ) );
NAND2_X2 _add_0_root_add_136_4_U411  ( .A1(_add_0_root_add_136_4_n328 ),.A2(_add_0_root_add_136_4_n329 ), .ZN(_add_0_root_add_136_4_n327 ) );
NAND2_X2 _add_0_root_add_136_4_U410  ( .A1(_add_0_root_add_136_4_n326 ),.A2(_add_0_root_add_136_4_n327 ), .ZN(_add_0_root_add_136_4_n324 ) );
NAND2_X2 _add_0_root_add_136_4_U409  ( .A1(_add_0_root_add_136_4_n314 ),.A2(_add_0_root_add_136_4_n307 ), .ZN(_add_0_root_add_136_4_n325 ) );
INV_X4 _add_0_root_add_136_4_U408  ( .A(N147), .ZN(_add_0_root_add_136_4_n322 ) );
INV_X4 _add_0_root_add_136_4_U407  ( .A(N115), .ZN(_add_0_root_add_136_4_n323 ) );
NOR2_X4 _add_0_root_add_136_4_U406  ( .A1(_add_0_root_add_136_4_n319 ), .A2(_add_0_root_add_136_4_n318 ), .ZN(_add_0_root_add_136_4_n317 ) );
XNOR2_X2 _add_0_root_add_136_4_U405  ( .A(_add_0_root_add_136_4_n258 ), .B(_add_0_root_add_136_4_n310 ), .ZN(next_A[1]) );
NOR2_X4 _add_0_root_add_136_4_U404  ( .A1(_add_0_root_add_136_4_n144 ), .A2(_add_0_root_add_136_4_n30 ), .ZN(_add_0_root_add_136_4_n308 ) );
NAND2_X2 _add_0_root_add_136_4_U403  ( .A1(_add_0_root_add_136_4_n307 ),.A2(_add_0_root_add_136_4_n184 ), .ZN(_add_0_root_add_136_4_n306 ) );
NOR2_X4 _add_0_root_add_136_4_U402  ( .A1(N148), .A2(N116), .ZN(_add_0_root_add_136_4_n282 ) );
XNOR2_X2 _add_0_root_add_136_4_U401  ( .A(_add_0_root_add_136_4_n299 ), .B(_add_0_root_add_136_4_n300 ), .ZN(next_A[20]) );
NOR2_X4 _add_0_root_add_136_4_U400  ( .A1(_add_0_root_add_136_4_n299 ), .A2(_add_0_root_add_136_4_n282 ), .ZN(_add_0_root_add_136_4_n298 ) );
NOR2_X4 _add_0_root_add_136_4_U399  ( .A1(_add_0_root_add_136_4_n291 ), .A2(_add_0_root_add_136_4_n88 ), .ZN(_add_0_root_add_136_4_n269 ) );
INV_X4 _add_0_root_add_136_4_U398  ( .A(N118), .ZN(_add_0_root_add_136_4_n289 ) );
INV_X4 _add_0_root_add_136_4_U397  ( .A(_add_0_root_add_136_4_n277 ), .ZN(_add_0_root_add_136_4_n270 ) );
XNOR2_X2 _add_0_root_add_136_4_U396  ( .A(_add_0_root_add_136_4_n286 ), .B(_add_0_root_add_136_4_n287 ), .ZN(next_A[22]) );
NAND2_X2 _add_0_root_add_136_4_U395  ( .A1(_add_0_root_add_136_4_n283 ),.A2(_add_0_root_add_136_4_n281 ), .ZN(_add_0_root_add_136_4_n276 ) );
NAND2_X2 _add_0_root_add_136_4_U394  ( .A1(_add_0_root_add_136_4_n70 ), .A2(_add_0_root_add_136_4_n8 ), .ZN(_add_0_root_add_136_4_n279 ) );
NAND2_X2 _add_0_root_add_136_4_U393  ( .A1(_add_0_root_add_136_4_n265 ),.A2(_add_0_root_add_136_4_n58 ), .ZN(_add_0_root_add_136_4_n275 ) );
XNOR2_X2 _add_0_root_add_136_4_U392  ( .A(_add_0_root_add_136_4_n261 ), .B(_add_0_root_add_136_4_n262 ), .ZN(next_A[24]) );
NAND3_X2 _add_0_root_add_136_4_U391  ( .A1(_add_0_root_add_136_4_n258 ),.A2(_add_0_root_add_136_4_n428 ), .A3(_add_0_root_add_136_4_n120 ),.ZN(_add_0_root_add_136_4_n257 ) );
NAND2_X2 _add_0_root_add_136_4_U390  ( .A1(_add_0_root_add_136_4_n252 ),.A2(_add_0_root_add_136_4_n253 ), .ZN(_add_0_root_add_136_4_n251 ) );
INV_X4 _add_0_root_add_136_4_U389  ( .A(_add_0_root_add_136_4_n232 ), .ZN(_add_0_root_add_136_4_n170 ) );
NAND3_X4 _add_0_root_add_136_4_U388  ( .A1(_add_0_root_add_136_4_n58 ), .A2(_add_0_root_add_136_4_n239 ), .A3(_add_0_root_add_136_4_n250 ), .ZN(_add_0_root_add_136_4_n142 ) );
NAND2_X2 _add_0_root_add_136_4_U387  ( .A1(_add_0_root_add_136_4_n247 ),.A2(_add_0_root_add_136_4_n246 ), .ZN(_add_0_root_add_136_4_n235 ) );
NAND2_X2 _add_0_root_add_136_4_U386  ( .A1(_add_0_root_add_136_4_n242 ),.A2(_add_0_root_add_136_4_n243 ), .ZN(_add_0_root_add_136_4_n241 ) );
INV_X4 _add_0_root_add_136_4_U385  ( .A(_add_0_root_add_136_4_n204 ), .ZN(_add_0_root_add_136_4_n225 ) );
XNOR2_X2 _add_0_root_add_136_4_U384  ( .A(_add_0_root_add_136_4_n193 ), .B(_add_0_root_add_136_4_n11 ), .ZN(next_A[25]) );
NAND2_X2 _add_0_root_add_136_4_U383  ( .A1(_add_0_root_add_136_4_n228 ),.A2(_add_0_root_add_136_4_n229 ), .ZN(_add_0_root_add_136_4_n227 ) );
NAND2_X2 _add_0_root_add_136_4_U382  ( .A1(N154), .A2(N122), .ZN(_add_0_root_add_136_4_n203 ) );
NAND2_X2 _add_0_root_add_136_4_U381  ( .A1(N155), .A2(N123), .ZN(_add_0_root_add_136_4_n200 ) );
INV_X4 _add_0_root_add_136_4_U380  ( .A(_add_0_root_add_136_4_n214 ), .ZN(_add_0_root_add_136_4_n205 ) );
NAND2_X2 _add_0_root_add_136_4_U379  ( .A1(_add_0_root_add_136_4_n209 ),.A2(_add_0_root_add_136_4_n48 ), .ZN(_add_0_root_add_136_4_n208 ) );
NAND2_X2 _add_0_root_add_136_4_U378  ( .A1(_add_0_root_add_136_4_n203 ),.A2(_add_0_root_add_136_4_n204 ), .ZN(_add_0_root_add_136_4_n202 ) );
NAND2_X2 _add_0_root_add_136_4_U377  ( .A1(_add_0_root_add_136_4_n201 ),.A2(_add_0_root_add_136_4_n202 ), .ZN(_add_0_root_add_136_4_n199 ) );
XNOR2_X2 _add_0_root_add_136_4_U376  ( .A(_add_0_root_add_136_4_n134 ), .B(_add_0_root_add_136_4_n187 ), .ZN(next_A[2]) );
INV_X4 _add_0_root_add_136_4_U375  ( .A(_add_0_root_add_136_4_n162 ), .ZN(_add_0_root_add_136_4_n141 ) );
INV_X4 _add_0_root_add_136_4_U374  ( .A(_add_0_root_add_136_4_n182 ), .ZN(_add_0_root_add_136_4_n181 ) );
NAND4_X2 _add_0_root_add_136_4_U373  ( .A1(N128), .A2(N96), .A3(_add_0_root_add_136_4_n180 ), .A4(_add_0_root_add_136_4_n181 ), .ZN(_add_0_root_add_136_4_n178 ) );
NAND4_X2 _add_0_root_add_136_4_U372  ( .A1(_add_0_root_add_136_4_n178 ),.A2(_add_0_root_add_136_4_n179 ), .A3(_add_0_root_add_136_4_n119 ),.A4(_add_0_root_add_136_4_n120 ), .ZN(_add_0_root_add_136_4_n177 ) );
NAND2_X2 _add_0_root_add_136_4_U371  ( .A1(_add_0_root_add_136_4_n176 ),.A2(_add_0_root_add_136_4_n177 ), .ZN(_add_0_root_add_136_4_n173 ) );
NAND2_X2 _add_0_root_add_136_4_U370  ( .A1(_add_0_root_add_136_4_n168 ),.A2(_add_0_root_add_136_4_n169 ), .ZN(_add_0_root_add_136_4_n167 ) );
NAND2_X2 _add_0_root_add_136_4_U369  ( .A1(_add_0_root_add_136_4_n161 ),.A2(_add_0_root_add_136_4_n26 ), .ZN(_add_0_root_add_136_4_n153 ) );
NAND2_X2 _add_0_root_add_136_4_U368  ( .A1(_add_0_root_add_136_4_n150 ),.A2(_add_0_root_add_136_4_n149 ), .ZN(_add_0_root_add_136_4_n159 ) );
NAND2_X2 _add_0_root_add_136_4_U367  ( .A1(_add_0_root_add_136_4_n160 ),.A2(_add_0_root_add_136_4_n141 ), .ZN(_add_0_root_add_136_4_n155 ) );
NAND4_X2 _add_0_root_add_136_4_U366  ( .A1(_add_0_root_add_136_4_n153 ),.A2(_add_0_root_add_136_4_n159 ), .A3(_add_0_root_add_136_4_n155 ),.A4(_add_0_root_add_136_4_n145 ), .ZN(_add_0_root_add_136_4_n158 ) );
NAND2_X2 _add_0_root_add_136_4_U365  ( .A1(N158), .A2(N126), .ZN(_add_0_root_add_136_4_n147 ) );
XNOR2_X2 _add_0_root_add_136_4_U364  ( .A(_add_0_root_add_136_4_n156 ), .B(_add_0_root_add_136_4_n13 ), .ZN(next_A[30]) );
INV_X4 _add_0_root_add_136_4_U363  ( .A(_add_0_root_add_136_4_n146 ), .ZN(_add_0_root_add_136_4_n154 ) );
XNOR2_X2 _add_0_root_add_136_4_U362  ( .A(N127), .B(N159), .ZN(_add_0_root_add_136_4_n136 ) );
XNOR2_X2 _add_0_root_add_136_4_U361  ( .A(_add_0_root_add_136_4_n135 ), .B(_add_0_root_add_136_4_n136 ), .ZN(next_A[31]) );
XNOR2_X2 _add_0_root_add_136_4_U360  ( .A(_add_0_root_add_136_4_n128 ), .B(_add_0_root_add_136_4_n129 ), .ZN(next_A[3]) );
XNOR2_X2 _add_0_root_add_136_4_U359  ( .A(_add_0_root_add_136_4_n122 ), .B(_add_0_root_add_136_4_n123 ), .ZN(next_A[5]) );
NAND2_X2 _add_0_root_add_136_4_U358  ( .A1(_add_0_root_add_136_4_n116 ),.A2(_add_0_root_add_136_4_n117 ), .ZN(_add_0_root_add_136_4_n115 ) );
XNOR2_X2 _add_0_root_add_136_4_U357  ( .A(_add_0_root_add_136_4_n113 ), .B(_add_0_root_add_136_4_n114 ), .ZN(next_A[6]) );
XNOR2_X2 _add_0_root_add_136_4_U356  ( .A(_add_0_root_add_136_4_n109 ), .B(_add_0_root_add_136_4_n110 ), .ZN(next_A[7]) );
INV_X4 _add_0_root_add_136_4_U355  ( .A(_add_0_root_add_136_4_n107 ), .ZN(_add_0_root_add_136_4_n97 ) );
XNOR2_X2 _add_0_root_add_136_4_U354  ( .A(_add_0_root_add_136_4_n105 ), .B(_add_0_root_add_136_4_n106 ), .ZN(next_A[8]) );
INV_X4 _add_0_root_add_136_4_U353  ( .A(_add_0_root_add_136_4_n96 ), .ZN(_add_0_root_add_136_4_n94 ) );
XNOR2_X2 _add_0_root_add_136_4_U352  ( .A(_add_0_root_add_136_4_n92 ), .B(_add_0_root_add_136_4_n93 ), .ZN(next_A[9]) );
NOR2_X1 _add_0_root_add_136_4_U351  ( .A1(_add_0_root_add_136_4_n360 ), .A2(_add_0_root_add_136_4_n175 ), .ZN(_add_0_root_add_136_4_n359 ) );
NAND3_X1 _add_0_root_add_136_4_U350  ( .A1(_add_0_root_add_136_4_n370 ),.A2(_add_0_root_add_136_4_n360 ), .A3(_add_0_root_add_136_4_n126 ),.ZN(_add_0_root_add_136_4_n369 ) );
NOR2_X1 _add_0_root_add_136_4_U349  ( .A1(_add_0_root_add_136_4_n175 ), .A2(_add_0_root_add_136_4_n91 ), .ZN(_add_0_root_add_136_4_n174 ) );
NOR2_X2 _add_0_root_add_136_4_U348  ( .A1(_add_0_root_add_136_4_n371 ), .A2(_add_0_root_add_136_4_n91 ), .ZN(_add_0_root_add_136_4_n367 ) );
NAND3_X2 _add_0_root_add_136_4_U347  ( .A1(_add_0_root_add_136_4_n232 ),.A2(_add_0_root_add_136_4_n233 ), .A3(_add_0_root_add_136_4_n234 ),.ZN(_add_0_root_add_136_4_n296 ) );
NAND3_X2 _add_0_root_add_136_4_U346  ( .A1(_add_0_root_add_136_4_n366 ),.A2(_add_0_root_add_136_4_n3 ), .A3(_add_0_root_add_136_4_n365 ), .ZN(_add_0_root_add_136_4_n364 ) );
INV_X2 _add_0_root_add_136_4_U345  ( .A(_add_0_root_add_136_4_n296 ), .ZN(_add_0_root_add_136_4_n272 ) );
INV_X1 _add_0_root_add_136_4_U344  ( .A(_add_0_root_add_136_4_n281 ), .ZN(_add_0_root_add_136_4_n268 ) );
NAND2_X4 _add_0_root_add_136_4_U343  ( .A1(_add_0_root_add_136_4_n288 ),.A2(_add_0_root_add_136_4_n289 ), .ZN(_add_0_root_add_136_4_n281 ) );
NAND2_X4 _add_0_root_add_136_4_U342  ( .A1(_add_0_root_add_136_4_n317 ),.A2(_add_0_root_add_136_4_n307 ), .ZN(_add_0_root_add_136_4_n171 ) );
NAND2_X4 _add_0_root_add_136_4_U341  ( .A1(_add_0_root_add_136_4_n335 ),.A2(_add_0_root_add_136_4_n336 ), .ZN(_add_0_root_add_136_4_n332 ) );
NAND4_X1 _add_0_root_add_136_4_U340  ( .A1(_add_0_root_add_136_4_n211 ),.A2(_add_0_root_add_136_4_n216 ), .A3(_add_0_root_add_136_4_n19 ),.A4(_add_0_root_add_136_4_n210 ), .ZN(_add_0_root_add_136_4_n230 ) );
NOR2_X2 _add_0_root_add_136_4_U339  ( .A1(_add_0_root_add_136_4_n230 ), .A2(_add_0_root_add_136_4_n70 ), .ZN(_add_0_root_add_136_4_n226 ) );
INV_X2 _add_0_root_add_136_4_U338  ( .A(_add_0_root_add_136_4_n206 ), .ZN(_add_0_root_add_136_4_n220 ) );
NAND2_X1 _add_0_root_add_136_4_U337  ( .A1(N111), .A2(N143), .ZN(_add_0_root_add_136_4_n343 ) );
INV_X8 _add_0_root_add_136_4_U336  ( .A(_add_0_root_add_136_4_n171 ), .ZN(_add_0_root_add_136_4_n304 ) );
NAND2_X4 _add_0_root_add_136_4_U335  ( .A1(_add_0_root_add_136_4_n231 ),.A2(_add_0_root_add_136_4_n244 ), .ZN(_add_0_root_add_136_4_n273 ) );
INV_X1 _add_0_root_add_136_4_U334  ( .A(_add_0_root_add_136_4_n150 ), .ZN(_add_0_root_add_136_4_n191 ) );
NAND3_X1 _add_0_root_add_136_4_U333  ( .A1(_add_0_root_add_136_4_n149 ),.A2(_add_0_root_add_136_4_n146 ), .A3(_add_0_root_add_136_4_n150 ),.ZN(_add_0_root_add_136_4_n148 ) );
NAND2_X1 _add_0_root_add_136_4_U332  ( .A1(_add_0_root_add_136_4_n342 ),.A2(_add_0_root_add_136_4_n343 ), .ZN(_add_0_root_add_136_4_n363 ) );
NOR3_X4 _add_0_root_add_136_4_U331  ( .A1(_add_0_root_add_136_4_n392 ), .A2(_add_0_root_add_136_4_n393 ), .A3(_add_0_root_add_136_4_n394 ), .ZN(_add_0_root_add_136_4_n391 ) );
NAND3_X1 _add_0_root_add_136_4_U330  ( .A1(_add_0_root_add_136_4_n360 ),.A2(_add_0_root_add_136_4_n126 ), .A3(_add_0_root_add_136_4_n370 ),.ZN(_add_0_root_add_136_4_n388 ) );
NAND3_X2 _add_0_root_add_136_4_U329  ( .A1(_add_0_root_add_136_4_n185 ),.A2(_add_0_root_add_136_4_n149 ), .A3(_add_0_root_add_136_4_n186 ),.ZN(_add_0_root_add_136_4_n162 ) );
NAND3_X2 _add_0_root_add_136_4_U328  ( .A1(_add_0_root_add_136_4_n193 ),.A2(_add_0_root_add_136_4_n185 ), .A3(_add_0_root_add_136_4_n48 ),.ZN(_add_0_root_add_136_4_n192 ) );
NAND3_X2 _add_0_root_add_136_4_U327  ( .A1(_add_0_root_add_136_4_n193 ),.A2(_add_0_root_add_136_4_n229 ), .A3(_add_0_root_add_136_4_n220 ),.ZN(_add_0_root_add_136_4_n219 ) );
NAND2_X1 _add_0_root_add_136_4_U326  ( .A1(_add_0_root_add_136_4_n250 ),.A2(_add_0_root_add_136_4_n58 ), .ZN(_add_0_root_add_136_4_n271 ) );
NAND2_X4 _add_0_root_add_136_4_U325  ( .A1(N115), .A2(_add_0_root_add_136_4_n90 ), .ZN(_add_0_root_add_136_4_n164 ) );
NAND2_X2 _add_0_root_add_136_4_U324  ( .A1(_add_0_root_add_136_4_n120 ),.A2(_add_0_root_add_136_4_n423 ), .ZN(_add_0_root_add_136_4_n126 ) );
AND2_X2 _add_0_root_add_136_4_U323  ( .A1(_add_0_root_add_136_4_n258 ), .A2(_add_0_root_add_136_4_n89 ), .ZN(next_A[0]) );
NAND3_X1 _add_0_root_add_136_4_U322  ( .A1(N97), .A2(N129), .A3(_add_0_root_add_136_4_n180 ), .ZN(_add_0_root_add_136_4_n179 ) );
NAND3_X2 _add_0_root_add_136_4_U321  ( .A1(_add_0_root_add_136_4_n137 ),.A2(_add_0_root_add_136_4_n138 ), .A3(_add_0_root_add_136_4_n139 ),.ZN(_add_0_root_add_136_4_n135 ) );
AND2_X2 _add_0_root_add_136_4_U320  ( .A1(N100), .A2(N132), .ZN(_add_0_root_add_136_4_n433 ) );
NOR2_X2 _add_0_root_add_136_4_U319  ( .A1(_add_0_root_add_136_4_n353 ), .A2(_add_0_root_add_136_4_n130 ), .ZN(_add_0_root_add_136_4_n352 ) );
NOR2_X2 _add_0_root_add_136_4_U318  ( .A1(_add_0_root_add_136_4_n431 ), .A2(_add_0_root_add_136_4_n435 ), .ZN(_add_0_root_add_136_4_n434 ) );
AND2_X2 _add_0_root_add_136_4_U317  ( .A1(N148), .A2(N116), .ZN(_add_0_root_add_136_4_n87 ) );
AND2_X2 _add_0_root_add_136_4_U316  ( .A1(N130), .A2(N98), .ZN(_add_0_root_add_136_4_n86 ) );
NOR2_X1 _add_0_root_add_136_4_U315  ( .A1(_add_0_root_add_136_4_n256 ), .A2(_add_0_root_add_136_4_n257 ), .ZN(_add_0_root_add_136_4_n254 ) );
NAND3_X1 _add_0_root_add_136_4_U314  ( .A1(_add_0_root_add_136_4_n174 ),.A2(_add_0_root_add_136_4_n108 ), .A3(_add_0_root_add_136_4_n173 ),.ZN(_add_0_root_add_136_4_n168 ) );
NOR2_X1 _add_0_root_add_136_4_U313  ( .A1(_add_0_root_add_136_4_n255 ), .A2(_add_0_root_add_136_4_n133 ), .ZN(_add_0_root_add_136_4_n350 ) );
NAND2_X2 _add_0_root_add_136_4_U312  ( .A1(N138), .A2(N106), .ZN(_add_0_root_add_136_4_n396 ) );
AND2_X2 _add_0_root_add_136_4_U311  ( .A1(N133), .A2(N101), .ZN(_add_0_root_add_136_4_n84 ) );
NAND3_X2 _add_0_root_add_136_4_U310  ( .A1(_add_0_root_add_136_4_n343 ),.A2(_add_0_root_add_136_4_n344 ), .A3(_add_0_root_add_136_4_n345 ),.ZN(_add_0_root_add_136_4_n309 ) );
AND2_X2 _add_0_root_add_136_4_U309  ( .A1(N134), .A2(N102), .ZN(_add_0_root_add_136_4_n83 ) );
NAND3_X2 _add_0_root_add_136_4_U308  ( .A1(N112), .A2(N144), .A3(_add_0_root_add_136_4_n332 ), .ZN(_add_0_root_add_136_4_n316 ) );
NOR2_X1 _add_0_root_add_136_4_U307  ( .A1(N99), .A2(_add_0_root_add_136_4_n29 ), .ZN(_add_0_root_add_136_4_n255 ) );
NOR2_X1 _add_0_root_add_136_4_U306  ( .A1(_add_0_root_add_136_4_n259 ), .A2(_add_0_root_add_136_4_n104 ), .ZN(_add_0_root_add_136_4_n252 ) );
NOR2_X2 _add_0_root_add_136_4_U305  ( .A1(_add_0_root_add_136_4_n254 ), .A2(_add_0_root_add_136_4_n255 ), .ZN(_add_0_root_add_136_4_n253 ) );
NAND3_X2 _add_0_root_add_136_4_U304  ( .A1(N98), .A2(N130), .A3(_add_0_root_add_136_4_n424 ), .ZN(_add_0_root_add_136_4_n119 ) );
AND2_X2 _add_0_root_add_136_4_U303  ( .A1(_add_0_root_add_136_4_n315 ), .A2(_add_0_root_add_136_4_n316 ), .ZN(_add_0_root_add_136_4_n326 ) );
NOR2_X2 _add_0_root_add_136_4_U302  ( .A1(_add_0_root_add_136_4_n85 ), .A2(_add_0_root_add_136_4_n83 ), .ZN(_add_0_root_add_136_4_n430 ) );
NAND3_X2 _add_0_root_add_136_4_U301  ( .A1(_add_0_root_add_136_4_n429 ),.A2(_add_0_root_add_136_4_n14 ), .A3(_add_0_root_add_136_4_n430 ),.ZN(_add_0_root_add_136_4_n401 ) );
NAND3_X2 _add_0_root_add_136_4_U300  ( .A1(_add_0_root_add_136_4_n316 ),.A2(_add_0_root_add_136_4_n315 ), .A3(_add_0_root_add_136_4_n314 ),.ZN(_add_0_root_add_136_4_n313 ) );
XNOR2_X2 _add_0_root_add_136_4_U299  ( .A(_add_0_root_add_136_4_n362 ), .B(_add_0_root_add_136_4_n363 ), .ZN(next_A[15]) );
NOR2_X1 _add_0_root_add_136_4_U298  ( .A1(_add_0_root_add_136_4_n104 ), .A2(_add_0_root_add_136_4_n183 ), .ZN(_add_0_root_add_136_4_n176 ) );
NOR2_X2 _add_0_root_add_136_4_U297  ( .A1(_add_0_root_add_136_4_n292 ), .A2(_add_0_root_add_136_4_n293 ), .ZN(_add_0_root_add_136_4_n290 ) );
NOR2_X2 _add_0_root_add_136_4_U296  ( .A1(_add_0_root_add_136_4_n410 ), .A2(_add_0_root_add_136_4_n411 ), .ZN(_add_0_root_add_136_4_n408 ) );
NOR2_X2 _add_0_root_add_136_4_U295  ( .A1(_add_0_root_add_136_4_n101 ), .A2(_add_0_root_add_136_4_n102 ), .ZN(_add_0_root_add_136_4_n99 ) );
NOR2_X2 _add_0_root_add_136_4_U294  ( .A1(_add_0_root_add_136_4_n99 ), .A2(_add_0_root_add_136_4_n100 ), .ZN(_add_0_root_add_136_4_n98 ) );
XNOR2_X2 _add_0_root_add_136_4_U293  ( .A(_add_0_root_add_136_4_n217 ), .B(_add_0_root_add_136_4_n218 ), .ZN(next_A[27]) );
XNOR2_X2 _add_0_root_add_136_4_U292  ( .A(_add_0_root_add_136_4_n333 ), .B(_add_0_root_add_136_4_n334 ), .ZN(next_A[17]) );
NOR2_X1 _add_0_root_add_136_4_U291  ( .A1(_add_0_root_add_136_4_n154 ), .A2(_add_0_root_add_136_4_n153 ), .ZN(_add_0_root_add_136_4_n152 ) );
NOR2_X1 _add_0_root_add_136_4_U290  ( .A1(_add_0_root_add_136_4_n154 ), .A2(_add_0_root_add_136_4_n155 ), .ZN(_add_0_root_add_136_4_n151 ) );
XNOR2_X2 _add_0_root_add_136_4_U289  ( .A(_add_0_root_add_136_4_n418 ), .B(_add_0_root_add_136_4_n77 ), .ZN(next_A[10]) );
NOR2_X1 _add_0_root_add_136_4_U288  ( .A1(_add_0_root_add_136_4_n100 ), .A2(_add_0_root_add_136_4_n95 ), .ZN(_add_0_root_add_136_4_n416 ) );
NAND3_X1 _add_0_root_add_136_4_U287  ( .A1(_add_0_root_add_136_4_n174 ),.A2(_add_0_root_add_136_4_n108 ), .A3(_add_0_root_add_136_4_n251 ),.ZN(_add_0_root_add_136_4_n246 ) );
NOR2_X2 _add_0_root_add_136_4_U286  ( .A1(_add_0_root_add_136_4_n115 ), .A2(_add_0_root_add_136_4_n435 ), .ZN(_add_0_root_add_136_4_n112 ) );
NOR2_X1 _add_0_root_add_136_4_U285  ( .A1(_add_0_root_add_136_4_n133 ), .A2(_add_0_root_add_136_4_n182 ), .ZN(_add_0_root_add_136_4_n260 ) );
NOR3_X1 _add_0_root_add_136_4_U284  ( .A1(_add_0_root_add_136_4_n256 ), .A2(_add_0_root_add_136_4_n130 ), .A3(_add_0_root_add_136_4_n260 ), .ZN(_add_0_root_add_136_4_n259 ) );
NOR2_X2 _add_0_root_add_136_4_U283  ( .A1(_add_0_root_add_136_4_n182 ), .A2(_add_0_root_add_136_4_n258 ), .ZN(_add_0_root_add_136_4_n188 ) );
NOR2_X2 _add_0_root_add_136_4_U282  ( .A1(_add_0_root_add_136_4_n9 ), .A2(_add_0_root_add_136_4_n188 ), .ZN(_add_0_root_add_136_4_n134 ) );
NAND3_X2 _add_0_root_add_136_4_U281  ( .A1(_add_0_root_add_136_4_n399 ),.A2(_add_0_root_add_136_4_n403 ), .A3(_add_0_root_add_136_4_n404 ),.ZN(_add_0_root_add_136_4_n402 ) );
AND2_X2 _add_0_root_add_136_4_U280  ( .A1(_add_0_root_add_136_4_n75 ), .A2(_add_0_root_add_136_4_n167 ), .ZN(_add_0_root_add_136_4_n143 ) );
XNOR2_X2 _add_0_root_add_136_4_U279  ( .A(_add_0_root_add_136_4_n274 ), .B(_add_0_root_add_136_4_n275 ), .ZN(next_A[23]) );
OR2_X4 _add_0_root_add_136_4_U278  ( .A1(_add_0_root_add_136_4_n154 ), .A2(_add_0_root_add_136_4_n145 ), .ZN(_add_0_root_add_136_4_n73 ) );
AND3_X2 _add_0_root_add_136_4_U277  ( .A1(_add_0_root_add_136_4_n148 ), .A2(_add_0_root_add_136_4_n147 ), .A3(_add_0_root_add_136_4_n73 ), .ZN(_add_0_root_add_136_4_n138 ) );
NOR2_X2 _add_0_root_add_136_4_U276  ( .A1(_add_0_root_add_136_4_n121 ), .A2(_add_0_root_add_136_4_n256 ), .ZN(_add_0_root_add_136_4_n423 ) );
NOR2_X1 _add_0_root_add_136_4_U275  ( .A1(_add_0_root_add_136_4_n83 ), .A2(_add_0_root_add_136_4_n431 ), .ZN(_add_0_root_add_136_4_n114 ) );
NOR2_X1 _add_0_root_add_136_4_U274  ( .A1(_add_0_root_add_136_4_n431 ), .A2(_add_0_root_add_136_4_n113 ), .ZN(_add_0_root_add_136_4_n111 ) );
NOR2_X2 _add_0_root_add_136_4_U273  ( .A1(_add_0_root_add_136_4_n111 ), .A2(_add_0_root_add_136_4_n83 ), .ZN(_add_0_root_add_136_4_n109 ) );
NOR2_X1 _add_0_root_add_136_4_U272  ( .A1(_add_0_root_add_136_4_n15 ), .A2(_add_0_root_add_136_4_n85 ), .ZN(_add_0_root_add_136_4_n110 ) );
NOR2_X1 _add_0_root_add_136_4_U271  ( .A1(_add_0_root_add_136_4_n100 ), .A2(_add_0_root_add_136_4_n97 ), .ZN(_add_0_root_add_136_4_n106 ) );
NOR2_X2 _add_0_root_add_136_4_U270  ( .A1(_add_0_root_add_136_4_n133 ), .A2(_add_0_root_add_136_4_n134 ), .ZN(_add_0_root_add_136_4_n132 ) );
NOR2_X1 _add_0_root_add_136_4_U269  ( .A1(_add_0_root_add_136_4_n130 ), .A2(_add_0_root_add_136_4_n131 ), .ZN(_add_0_root_add_136_4_n129 ) );
NOR2_X2 _add_0_root_add_136_4_U268  ( .A1(_add_0_root_add_136_4_n132 ), .A2(_add_0_root_add_136_4_n86 ), .ZN(_add_0_root_add_136_4_n128 ) );
NOR2_X2 _add_0_root_add_136_4_U267  ( .A1(_add_0_root_add_136_4_n86 ), .A2(_add_0_root_add_136_4_n133 ), .ZN(_add_0_root_add_136_4_n187 ) );
NOR2_X2 _add_0_root_add_136_4_U266  ( .A1(_add_0_root_add_136_4_n97 ), .A2(_add_0_root_add_136_4_n98 ), .ZN(_add_0_root_add_136_4_n92 ) );
NOR2_X1 _add_0_root_add_136_4_U265  ( .A1(_add_0_root_add_136_4_n94 ), .A2(_add_0_root_add_136_4_n95 ), .ZN(_add_0_root_add_136_4_n93 ) );
NOR2_X1 _add_0_root_add_136_4_U264  ( .A1(_add_0_root_add_136_4_n103 ), .A2(_add_0_root_add_136_4_n125 ), .ZN(_add_0_root_add_136_4_n124 ) );
NOR2_X2 _add_0_root_add_136_4_U263  ( .A1(_add_0_root_add_136_4_n124 ), .A2(_add_0_root_add_136_4_n10 ), .ZN(_add_0_root_add_136_4_n122 ) );
XNOR2_X2 _add_0_root_add_136_4_U262  ( .A(_add_0_root_add_136_4_n324 ), .B(_add_0_root_add_136_4_n325 ), .ZN(next_A[18]) );
NAND3_X2 _add_0_root_add_136_4_U261  ( .A1(_add_0_root_add_136_4_n232 ),.A2(_add_0_root_add_136_4_n234 ), .A3(_add_0_root_add_136_4_n303 ),.ZN(_add_0_root_add_136_4_n331 ) );
NOR2_X1 _add_0_root_add_136_4_U260  ( .A1(_add_0_root_add_136_4_n154 ), .A2(_add_0_root_add_136_4_n2 ), .ZN(_add_0_root_add_136_4_n140 ) );
NOR2_X1 _add_0_root_add_136_4_U259  ( .A1(_add_0_root_add_136_4_n175 ), .A2(_add_0_root_add_136_4_n380 ), .ZN(_add_0_root_add_136_4_n387 ) );
INV_X1 _add_0_root_add_136_4_U258  ( .A(_add_0_root_add_136_4_n133 ), .ZN(_add_0_root_add_136_4_n180 ) );
OR2_X1 _add_0_root_add_136_4_U257  ( .A1(N96), .A2(N128), .ZN(_add_0_root_add_136_4_n89 ) );
OR2_X4 _add_0_root_add_136_4_U256  ( .A1(N140), .A2(N108), .ZN(_add_0_root_add_136_4_n355 ) );
OR2_X4 _add_0_root_add_136_4_U255  ( .A1(N155), .A2(N123), .ZN(_add_0_root_add_136_4_n214 ) );
NOR2_X1 _add_0_root_add_136_4_U254  ( .A1(N100), .A2(N132), .ZN(_add_0_root_add_136_4_n125 ) );
OR2_X4 _add_0_root_add_136_4_U253  ( .A1(N158), .A2(N126), .ZN(_add_0_root_add_136_4_n146 ) );
NOR2_X4 _add_0_root_add_136_4_U252  ( .A1(N112), .A2(N144), .ZN(_add_0_root_add_136_4_n318 ) );
NAND2_X1 _add_0_root_add_136_4_U251  ( .A1(_add_0_root_add_136_4_n352 ),.A2(_add_0_root_add_136_4_n119 ), .ZN(_add_0_root_add_136_4_n351 ) );
NAND2_X1 _add_0_root_add_136_4_U250  ( .A1(_add_0_root_add_136_4_n399 ),.A2(_add_0_root_add_136_4_n395 ), .ZN(_add_0_root_add_136_4_n406 ) );
INV_X2 _add_0_root_add_136_4_U249  ( .A(_add_0_root_add_136_4_n212 ), .ZN(_add_0_root_add_136_4_n229 ) );
NOR2_X1 _add_0_root_add_136_4_U248  ( .A1(_add_0_root_add_136_4_n151 ), .A2(_add_0_root_add_136_4_n152 ), .ZN(_add_0_root_add_136_4_n137 ) );
OR3_X4 _add_0_root_add_136_4_U247  ( .A1(_add_0_root_add_136_4_n348 ), .A2(_add_0_root_add_136_4_n349 ), .A3(_add_0_root_add_136_4_n104 ), .ZN(_add_0_root_add_136_4_n72 ) );
NOR2_X2 _add_0_root_add_136_4_U246  ( .A1(_add_0_root_add_136_4_n417 ), .A2(_add_0_root_add_136_4_n101 ), .ZN(_add_0_root_add_136_4_n410 ) );
OR2_X4 _add_0_root_add_136_4_U245  ( .A1(_add_0_root_add_136_4_n206 ), .A2(_add_0_root_add_136_4_n204 ), .ZN(_add_0_root_add_136_4_n82 ) );
XOR2_X1 _add_0_root_add_136_4_U244  ( .A(_add_0_root_add_136_4_n126 ), .B(_add_0_root_add_136_4_n127 ), .Z(next_A[4]) );
INV_X1 _add_0_root_add_136_4_U243  ( .A(_add_0_root_add_136_4_n203 ), .ZN(_add_0_root_add_136_4_n223 ) );
NAND3_X2 _add_0_root_add_136_4_U242  ( .A1(_add_0_root_add_136_4_n357 ),.A2(_add_0_root_add_136_4_n356 ), .A3(_add_0_root_add_136_4_n355 ),.ZN(_add_0_root_add_136_4_n172 ) );
NOR2_X2 _add_0_root_add_136_4_U241  ( .A1(_add_0_root_add_136_4_n24 ), .A2(_add_0_root_add_136_4_n245 ), .ZN(_add_0_root_add_136_4_n166 ) );
NOR2_X1 _add_0_root_add_136_4_U240  ( .A1(_add_0_root_add_136_4_n101 ), .A2(_add_0_root_add_136_4_n102 ), .ZN(_add_0_root_add_136_4_n105 ) );
NOR2_X1 _add_0_root_add_136_4_U239  ( .A1(_add_0_root_add_136_4_n9 ), .A2(_add_0_root_add_136_4_n182 ), .ZN(_add_0_root_add_136_4_n310 ) );
NOR2_X1 _add_0_root_add_136_4_U238  ( .A1(_add_0_root_add_136_4_n84 ), .A2(_add_0_root_add_136_4_n435 ), .ZN(_add_0_root_add_136_4_n123 ) );
INV_X2 _add_0_root_add_136_4_U237  ( .A(_add_0_root_add_136_4_n337 ), .ZN(_add_0_root_add_136_4_n361 ) );
NOR2_X4 _add_0_root_add_136_4_U236  ( .A1(_add_0_root_add_136_4_n65 ), .A2(_add_0_root_add_136_4_n66 ), .ZN(_add_0_root_add_136_4_n379 ) );
NOR2_X1 _add_0_root_add_136_4_U235  ( .A1(_add_0_root_add_136_4_n121 ), .A2(_add_0_root_add_136_4_n10 ), .ZN(_add_0_root_add_136_4_n118 ) );
NAND3_X1 _add_0_root_add_136_4_U234  ( .A1(_add_0_root_add_136_4_n119 ),.A2(_add_0_root_add_136_4_n120 ), .A3(_add_0_root_add_136_4_n118 ),.ZN(_add_0_root_add_136_4_n117 ) );
NOR2_X4 _add_0_root_add_136_4_U233  ( .A1(_add_0_root_add_136_4_n224 ), .A2(_add_0_root_add_136_4_n225 ), .ZN(_add_0_root_add_136_4_n221 ) );
NOR2_X1 _add_0_root_add_136_4_U232  ( .A1(_add_0_root_add_136_4_n125 ), .A2(_add_0_root_add_136_4_n10 ), .ZN(_add_0_root_add_136_4_n127 ) );
NAND2_X4 _add_0_root_add_136_4_U231  ( .A1(_add_0_root_add_136_4_n61 ), .A2(_add_0_root_add_136_4_n62 ), .ZN(next_A[26]) );
NAND2_X1 _add_0_root_add_136_4_U230  ( .A1(_add_0_root_add_136_4_n149 ),.A2(_add_0_root_add_136_4_n145 ), .ZN(_add_0_root_add_136_4_n190 ) );
NOR2_X4 _add_0_root_add_136_4_U229  ( .A1(_add_0_root_add_136_4_n91 ), .A2(_add_0_root_add_136_4_n175 ), .ZN(_add_0_root_add_136_4_n347 ) );
OR2_X4 _add_0_root_add_136_4_U228  ( .A1(_add_0_root_add_136_4_n45 ), .A2(N119), .ZN(_add_0_root_add_136_4_n58 ) );
INV_X2 _add_0_root_add_136_4_U227  ( .A(_add_0_root_add_136_4_n222 ), .ZN(_add_0_root_add_136_4_n60 ) );
NOR2_X1 _add_0_root_add_136_4_U226  ( .A1(_add_0_root_add_136_4_n51 ), .A2(_add_0_root_add_136_4_n88 ), .ZN(_add_0_root_add_136_4_n297 ) );
INV_X1 _add_0_root_add_136_4_U225  ( .A(_add_0_root_add_136_4_n297 ), .ZN(_add_0_root_add_136_4_n55 ) );
NAND2_X4 _add_0_root_add_136_4_U224  ( .A1(_add_0_root_add_136_4_n57 ), .A2(_add_0_root_add_136_4_n56 ), .ZN(next_A[21]) );
NAND2_X4 _add_0_root_add_136_4_U223  ( .A1(_add_0_root_add_136_4_n43 ), .A2(_add_0_root_add_136_4_n55 ), .ZN(_add_0_root_add_136_4_n57 ) );
NAND2_X4 _add_0_root_add_136_4_U222  ( .A1(_add_0_root_add_136_4_n236 ),.A2(_add_0_root_add_136_4_n235 ), .ZN(_add_0_root_add_136_4_n193 ) );
NOR2_X2 _add_0_root_add_136_4_U221  ( .A1(N99), .A2(N131), .ZN(_add_0_root_add_136_4_n183 ) );
NOR2_X2 _add_0_root_add_136_4_U220  ( .A1(_add_0_root_add_136_4_n5 ), .A2(_add_0_root_add_136_4_n162 ), .ZN(_add_0_root_add_136_4_n161 ) );
NOR2_X4 _add_0_root_add_136_4_U219  ( .A1(N149), .A2(N117), .ZN(_add_0_root_add_136_4_n88 ) );
NAND3_X2 _add_0_root_add_136_4_U218  ( .A1(_add_0_root_add_136_4_n219 ),.A2(_add_0_root_add_136_4_n203 ), .A3(_add_0_root_add_136_4_n82 ),.ZN(_add_0_root_add_136_4_n217 ) );
NAND2_X4 _add_0_root_add_136_4_U217  ( .A1(_add_0_root_add_136_4_n322 ),.A2(_add_0_root_add_136_4_n323 ), .ZN(_add_0_root_add_136_4_n184 ) );
NAND3_X4 _add_0_root_add_136_4_U216  ( .A1(_add_0_root_add_136_4_n303 ),.A2(_add_0_root_add_136_4_n23 ), .A3(_add_0_root_add_136_4_n304 ),.ZN(_add_0_root_add_136_4_n248 ) );
NAND3_X1 _add_0_root_add_136_4_U215  ( .A1(_add_0_root_add_136_4_n360 ),.A2(_add_0_root_add_136_4_n400 ), .A3(_add_0_root_add_136_4_n401 ),.ZN(_add_0_root_add_136_4_n368 ) );
NAND2_X4 _add_0_root_add_136_4_U214  ( .A1(_add_0_root_add_136_4_n401 ),.A2(_add_0_root_add_136_4_n400 ), .ZN(_add_0_root_add_136_4_n108 ) );
NAND2_X1 _add_0_root_add_136_4_U213  ( .A1(N156), .A2(N124), .ZN(_add_0_root_add_136_4_n195 ) );
NAND2_X1 _add_0_root_add_136_4_U212  ( .A1(N157), .A2(N125), .ZN(_add_0_root_add_136_4_n145 ) );
NAND2_X4 _add_0_root_add_136_4_U211  ( .A1(_add_0_root_add_136_4_n194 ),.A2(_add_0_root_add_136_4_n195 ), .ZN(_add_0_root_add_136_4_n150 ) );
NAND2_X2 _add_0_root_add_136_4_U210  ( .A1(_add_0_root_add_136_4_n17 ), .A2(_add_0_root_add_136_4_n388 ), .ZN(_add_0_root_add_136_4_n66 ) );
NOR3_X4 _add_0_root_add_136_4_U209  ( .A1(_add_0_root_add_136_4_n213 ), .A2(_add_0_root_add_136_4_n212 ), .A3(_add_0_root_add_136_4_n205 ), .ZN(_add_0_root_add_136_4_n186 ) );
NAND2_X1 _add_0_root_add_136_4_U208  ( .A1(_add_0_root_add_136_4_n141 ),.A2(_add_0_root_add_136_4_n23 ), .ZN(_add_0_root_add_136_4_n163 ) );
NOR3_X2 _add_0_root_add_136_4_U207  ( .A1(_add_0_root_add_136_4_n163 ), .A2(_add_0_root_add_136_4_n143 ), .A3(_add_0_root_add_136_4_n21 ), .ZN(_add_0_root_add_136_4_n157 ) );
NAND3_X1 _add_0_root_add_136_4_U206  ( .A1(_add_0_root_add_136_4_n367 ),.A2(_add_0_root_add_136_4_n368 ), .A3(_add_0_root_add_136_4_n369 ),.ZN(_add_0_root_add_136_4_n366 ) );
INV_X2 _add_0_root_add_136_4_U205  ( .A(_add_0_root_add_136_4_n368 ), .ZN(_add_0_root_add_136_4_n65 ) );
NAND3_X2 _add_0_root_add_136_4_U204  ( .A1(_add_0_root_add_136_4_n243 ),.A2(_add_0_root_add_136_4_n231 ), .A3(_add_0_root_add_136_4_n244 ),.ZN(_add_0_root_add_136_4_n240 ) );
NOR3_X1 _add_0_root_add_136_4_U203  ( .A1(_add_0_root_add_136_4_n170 ), .A2(_add_0_root_add_136_4_n16 ), .A3(_add_0_root_add_136_4_n4 ), .ZN(_add_0_root_add_136_4_n169 ) );
NAND2_X2 _add_0_root_add_136_4_U202  ( .A1(_add_0_root_add_136_4_n330 ),.A2(_add_0_root_add_136_4_n331 ), .ZN(_add_0_root_add_136_4_n329 ) );
NOR2_X4 _add_0_root_add_136_4_U201  ( .A1(N154), .A2(N122), .ZN(_add_0_root_add_136_4_n206 ) );
NOR2_X2 _add_0_root_add_136_4_U200  ( .A1(_add_0_root_add_136_4_n223 ), .A2(_add_0_root_add_136_4_n206 ), .ZN(_add_0_root_add_136_4_n222 ) );
OR2_X4 _add_0_root_add_136_4_U199  ( .A1(N139), .A2(N107), .ZN(_add_0_root_add_136_4_n399 ) );
INV_X1 _add_0_root_add_136_4_U198  ( .A(_add_0_root_add_136_4_n335 ), .ZN(_add_0_root_add_136_4_n54 ) );
AND2_X2 _add_0_root_add_136_4_U197  ( .A1(_add_0_root_add_136_4_n185 ), .A2(_add_0_root_add_136_4_n195 ), .ZN(_add_0_root_add_136_4_n53 ) );
XNOR2_X2 _add_0_root_add_136_4_U196  ( .A(_add_0_root_add_136_4_n197 ), .B(_add_0_root_add_136_4_n53 ), .ZN(next_A[28]) );
NOR2_X4 _add_0_root_add_136_4_U195  ( .A1(_add_0_root_add_136_4_n226 ), .A2(_add_0_root_add_136_4_n227 ), .ZN(_add_0_root_add_136_4_n224 ) );
NOR3_X4 _add_0_root_add_136_4_U194  ( .A1(_add_0_root_add_136_4_n269 ), .A2(_add_0_root_add_136_4_n51 ), .A3(_add_0_root_add_136_4_n270 ), .ZN(_add_0_root_add_136_4_n267 ) );
NAND2_X4 _add_0_root_add_136_4_U193  ( .A1(_add_0_root_add_136_4_n17 ), .A2(_add_0_root_add_136_4_n359 ), .ZN(_add_0_root_add_136_4_n232 ) );
INV_X8 _add_0_root_add_136_4_U192  ( .A(_add_0_root_add_136_4_n280 ), .ZN(_add_0_root_add_136_4_n250 ) );
INV_X2 _add_0_root_add_136_4_U191  ( .A(_add_0_root_add_136_4_n378 ), .ZN(_add_0_root_add_136_4_n386 ) );
NOR2_X4 _add_0_root_add_136_4_U190  ( .A1(_add_0_root_add_136_4_n47 ), .A2(_add_0_root_add_136_4_n267 ), .ZN(_add_0_root_add_136_4_n266 ) );
NAND2_X2 _add_0_root_add_136_4_U189  ( .A1(_add_0_root_add_136_4_n416 ),.A2(_add_0_root_add_136_4_n420 ), .ZN(_add_0_root_add_136_4_n419 ) );
INV_X2 _add_0_root_add_136_4_U188  ( .A(_add_0_root_add_136_4_n331 ), .ZN(_add_0_root_add_136_4_n320 ) );
NAND4_X1 _add_0_root_add_136_4_U187  ( .A1(_add_0_root_add_136_4_n276 ),.A2(_add_0_root_add_136_4_n277 ), .A3(_add_0_root_add_136_4_n278 ),.A4(_add_0_root_add_136_4_n279 ), .ZN(_add_0_root_add_136_4_n274 ) );
NAND2_X2 _add_0_root_add_136_4_U186  ( .A1(_add_0_root_add_136_4_n167 ),.A2(_add_0_root_add_136_4_n75 ), .ZN(_add_0_root_add_136_4_n50 ) );
OR2_X2 _add_0_root_add_136_4_U185  ( .A1(_add_0_root_add_136_4_n24 ), .A2(_add_0_root_add_136_4_n245 ), .ZN(_add_0_root_add_136_4_n49 ) );
NAND2_X4 _add_0_root_add_136_4_U184  ( .A1(_add_0_root_add_136_4_n306 ),.A2(_add_0_root_add_136_4_n164 ), .ZN(_add_0_root_add_136_4_n231 ) );
INV_X4 _add_0_root_add_136_4_U183  ( .A(_add_0_root_add_136_4_n266 ), .ZN(_add_0_root_add_136_4_n264 ) );
NAND2_X4 _add_0_root_add_136_4_U182  ( .A1(_add_0_root_add_136_4_n199 ),.A2(_add_0_root_add_136_4_n200 ), .ZN(_add_0_root_add_136_4_n196 ) );
NAND2_X4 _add_0_root_add_136_4_U181  ( .A1(_add_0_root_add_136_4_n196 ),.A2(_add_0_root_add_136_4_n185 ), .ZN(_add_0_root_add_136_4_n194 ) );
OR2_X2 _add_0_root_add_136_4_U180  ( .A1(_add_0_root_add_136_4_n379 ), .A2(_add_0_root_add_136_4_n380 ), .ZN(_add_0_root_add_136_4_n71 ) );
NAND2_X2 _add_0_root_add_136_4_U179  ( .A1(_add_0_root_add_136_4_n338 ),.A2(_add_0_root_add_136_4_n337 ), .ZN(_add_0_root_add_136_4_n333 ) );
NOR3_X2 _add_0_root_add_136_4_U178  ( .A1(_add_0_root_add_136_4_n170 ), .A2(_add_0_root_add_136_4_n22 ), .A3(_add_0_root_add_136_4_n142 ), .ZN(_add_0_root_add_136_4_n247 ) );
INV_X2 _add_0_root_add_136_4_U177  ( .A(_add_0_root_add_136_4_n322 ), .ZN(_add_0_root_add_136_4_n90 ) );
NAND2_X4 _add_0_root_add_136_4_U176  ( .A1(_add_0_root_add_136_4_n63 ), .A2(_add_0_root_add_136_4_n64 ), .ZN(next_A[29]) );
NAND2_X4 _add_0_root_add_136_4_U175  ( .A1(_add_0_root_add_136_4_n189 ),.A2(_add_0_root_add_136_4_n190 ), .ZN(_add_0_root_add_136_4_n63 ) );
INV_X8 _add_0_root_add_136_4_U174  ( .A(_add_0_root_add_136_4_n248 ), .ZN(_add_0_root_add_136_4_n233 ) );
NOR2_X1 _add_0_root_add_136_4_U173  ( .A1(_add_0_root_add_136_4_n150 ), .A2(_add_0_root_add_136_4_n190 ), .ZN(_add_0_root_add_136_4_n46 ) );
NOR2_X4 _add_0_root_add_136_4_U172  ( .A1(_add_0_root_add_136_4_n312 ), .A2(_add_0_root_add_136_4_n166 ), .ZN(_add_0_root_add_136_4_n311 ) );
NAND2_X2 _add_0_root_add_136_4_U171  ( .A1(_add_0_root_add_136_4_n192 ),.A2(_add_0_root_add_136_4_n46 ), .ZN(_add_0_root_add_136_4_n64 ) );
NOR2_X2 _add_0_root_add_136_4_U170  ( .A1(N122), .A2(N154), .ZN(_add_0_root_add_136_4_n213 ) );
NAND2_X4 _add_0_root_add_136_4_U169  ( .A1(_add_0_root_add_136_4_n40 ), .A2(_add_0_root_add_136_4_n41 ), .ZN(_add_0_root_add_136_4_n43 ) );
INV_X4 _add_0_root_add_136_4_U168  ( .A(_add_0_root_add_136_4_n298 ), .ZN(_add_0_root_add_136_4_n40 ) );
AND2_X2 _add_0_root_add_136_4_U167  ( .A1(_add_0_root_add_136_4_n297 ), .A2(_add_0_root_add_136_4_n41 ), .ZN(_add_0_root_add_136_4_n42 ) );
OR2_X4 _add_0_root_add_136_4_U166  ( .A1(N156), .A2(N124), .ZN(_add_0_root_add_136_4_n185 ) );
OR2_X4 _add_0_root_add_136_4_U165  ( .A1(N157), .A2(N125), .ZN(_add_0_root_add_136_4_n149 ) );
NOR2_X2 _add_0_root_add_136_4_U164  ( .A1(_add_0_root_add_136_4_n397 ), .A2(_add_0_root_add_136_4_n398 ), .ZN(_add_0_root_add_136_4_n393 ) );
NOR3_X2 _add_0_root_add_136_4_U163  ( .A1(_add_0_root_add_136_4_n397 ), .A2(_add_0_root_add_136_4_n107 ), .A3(_add_0_root_add_136_4_n95 ), .ZN(_add_0_root_add_136_4_n392 ) );
NOR2_X4 _add_0_root_add_136_4_U162  ( .A1(N138), .A2(N106), .ZN(_add_0_root_add_136_4_n397 ) );
INV_X8 _add_0_root_add_136_4_U161  ( .A(_add_0_root_add_136_4_n210 ), .ZN(_add_0_root_add_136_4_n160 ) );
NAND2_X4 _add_0_root_add_136_4_U160  ( .A1(_add_0_root_add_136_4_n52 ), .A2(N120), .ZN(_add_0_root_add_136_4_n210 ) );
NOR2_X2 _add_0_root_add_136_4_U159  ( .A1(_add_0_root_add_136_4_n215 ), .A2(_add_0_root_add_136_4_n160 ), .ZN(_add_0_root_add_136_4_n39 ) );
AND2_X2 _add_0_root_add_136_4_U158  ( .A1(_add_0_root_add_136_4_n211 ), .A2(_add_0_root_add_136_4_n39 ), .ZN(_add_0_root_add_136_4_n207 ) );
AND3_X4 _add_0_root_add_136_4_U157  ( .A1(_add_0_root_add_136_4_n232 ), .A2(_add_0_root_add_136_4_n233 ), .A3(_add_0_root_add_136_4_n234 ), .ZN(_add_0_root_add_136_4_n70 ) );
NAND2_X4 _add_0_root_add_136_4_U156  ( .A1(_add_0_root_add_136_4_n240 ),.A2(_add_0_root_add_136_4_n241 ), .ZN(_add_0_root_add_136_4_n237 ) );
NOR3_X4 _add_0_root_add_136_4_U155  ( .A1(_add_0_root_add_136_4_n237 ), .A2(_add_0_root_add_136_4_n160 ), .A3(_add_0_root_add_136_4_n238 ), .ZN(_add_0_root_add_136_4_n236 ) );
NAND2_X1 _add_0_root_add_136_4_U154  ( .A1(_add_0_root_add_136_4_n315 ),.A2(_add_0_root_add_136_4_n332 ), .ZN(_add_0_root_add_136_4_n334 ) );
INV_X4 _add_0_root_add_136_4_U153  ( .A(_add_0_root_add_136_4_n221 ), .ZN(_add_0_root_add_136_4_n59 ) );
BUF_X16 _add_0_root_add_136_4_U152  ( .A(N138), .Z(_add_0_root_add_136_4_n37 ) );
AND2_X2 _add_0_root_add_136_4_U151  ( .A1(_add_0_root_add_136_4_n344 ), .A2(_add_0_root_add_136_4_n346 ), .ZN(_add_0_root_add_136_4_n36 ) );
XNOR2_X2 _add_0_root_add_136_4_U150  ( .A(_add_0_root_add_136_4_n373 ), .B(_add_0_root_add_136_4_n36 ), .ZN(next_A[14]) );
NAND2_X4 _add_0_root_add_136_4_U149  ( .A1(N153), .A2(N121), .ZN(_add_0_root_add_136_4_n204 ) );
NOR2_X2 _add_0_root_add_136_4_U148  ( .A1(_add_0_root_add_136_4_n379 ), .A2(_add_0_root_add_136_4_n81 ), .ZN(_add_0_root_add_136_4_n374 ) );
INV_X2 _add_0_root_add_136_4_U147  ( .A(_add_0_root_add_136_4_n397 ), .ZN(_add_0_root_add_136_4_n403 ) );
INV_X1 _add_0_root_add_136_4_U146  ( .A(_add_0_root_add_136_4_n304 ), .ZN(_add_0_root_add_136_4_n33 ) );
AND2_X2 _add_0_root_add_136_4_U145  ( .A1(_add_0_root_add_136_4_n164 ), .A2(_add_0_root_add_136_4_n23 ), .ZN(_add_0_root_add_136_4_n32 ) );
XNOR2_X2 _add_0_root_add_136_4_U144  ( .A(_add_0_root_add_136_4_n311 ), .B(_add_0_root_add_136_4_n32 ), .ZN(next_A[19]) );
INV_X2 _add_0_root_add_136_4_U143  ( .A(_add_0_root_add_136_4_n38 ), .ZN(_add_0_root_add_136_4_n342 ) );
INV_X4 _add_0_root_add_136_4_U142  ( .A(_add_0_root_add_136_4_n332 ), .ZN(_add_0_root_add_136_4_n319 ) );
NOR2_X2 _add_0_root_add_136_4_U141  ( .A1(_add_0_root_add_136_4_n319 ), .A2(_add_0_root_add_136_4_n318 ), .ZN(_add_0_root_add_136_4_n328 ) );
NAND2_X2 _add_0_root_add_136_4_U140  ( .A1(_add_0_root_add_136_4_n192 ),.A2(_add_0_root_add_136_4_n191 ), .ZN(_add_0_root_add_136_4_n189 ) );
INV_X2 _add_0_root_add_136_4_U139  ( .A(_add_0_root_add_136_4_n87 ), .ZN(_add_0_root_add_136_4_n41 ) );
INV_X2 _add_0_root_add_136_4_U138  ( .A(_add_0_root_add_136_4_n28 ), .ZN(_add_0_root_add_136_4_n29 ) );
INV_X1 _add_0_root_add_136_4_U137  ( .A(N131), .ZN(_add_0_root_add_136_4_n28 ) );
INV_X4 _add_0_root_add_136_4_U136  ( .A(_add_0_root_add_136_4_n27 ), .ZN(_add_0_root_add_136_4_n101 ) );
OR2_X2 _add_0_root_add_136_4_U135  ( .A1(_add_0_root_add_136_4_n103 ), .A2(_add_0_root_add_136_4_n104 ), .ZN(_add_0_root_add_136_4_n27 ) );
NOR2_X4 _add_0_root_add_136_4_U134  ( .A1(_add_0_root_add_136_4_n320 ), .A2(_add_0_root_add_136_4_n321 ), .ZN(_add_0_root_add_136_4_n341 ) );
XNOR2_X1 _add_0_root_add_136_4_U133  ( .A(_add_0_root_add_136_4_n341 ), .B(_add_0_root_add_136_4_n340 ), .ZN(next_A[16]) );
NAND3_X1 _add_0_root_add_136_4_U132  ( .A1(_add_0_root_add_136_4_n216 ),.A2(_add_0_root_add_136_4_n19 ), .A3(_add_0_root_add_136_4_n296 ),.ZN(_add_0_root_add_136_4_n215 ) );
NAND2_X2 _add_0_root_add_136_4_U131  ( .A1(_add_0_root_add_136_4_n216 ),.A2(_add_0_root_add_136_4_n6 ), .ZN(_add_0_root_add_136_4_n295 ) );
NAND2_X2 _add_0_root_add_136_4_U130  ( .A1(N116), .A2(N148), .ZN(_add_0_root_add_136_4_n291 ) );
NAND2_X2 _add_0_root_add_136_4_U129  ( .A1(_add_0_root_add_136_4_n249 ),.A2(_add_0_root_add_136_4_n281 ), .ZN(_add_0_root_add_136_4_n47 ) );
INV_X2 _add_0_root_add_136_4_U128  ( .A(_add_0_root_add_136_4_n414 ), .ZN(_add_0_root_add_136_4_n413 ) );
OR2_X2 _add_0_root_add_136_4_U127  ( .A1(_add_0_root_add_136_4_n409 ), .A2(_add_0_root_add_136_4_n414 ), .ZN(_add_0_root_add_136_4_n77 ) );
INV_X1 _add_0_root_add_136_4_U126  ( .A(_add_0_root_add_136_4_n396 ), .ZN(_add_0_root_add_136_4_n409 ) );
NOR2_X4 _add_0_root_add_136_4_U125  ( .A1(N143), .A2(N111), .ZN(_add_0_root_add_136_4_n38 ) );
NOR2_X4 _add_0_root_add_136_4_U124  ( .A1(_add_0_root_add_136_4_n38 ), .A2(_add_0_root_add_136_4_n358 ), .ZN(_add_0_root_add_136_4_n357 ) );
NAND3_X1 _add_0_root_add_136_4_U123  ( .A1(_add_0_root_add_136_4_n346 ),.A2(N109), .A3(N141), .ZN(_add_0_root_add_136_4_n345 ) );
NAND3_X1 _add_0_root_add_136_4_U122  ( .A1(_add_0_root_add_136_4_n107 ),.A2(_add_0_root_add_136_4_n108 ), .A3(_add_0_root_add_136_4_n27 ),.ZN(_add_0_root_add_136_4_n420 ) );
INV_X1 _add_0_root_add_136_4_U121  ( .A(_add_0_root_add_136_4_n34 ), .ZN(_add_0_root_add_136_4_n400 ) );
OR2_X2 _add_0_root_add_136_4_U120  ( .A1(N151), .A2(N119), .ZN(_add_0_root_add_136_4_n249 ) );
INV_X4 _add_0_root_add_136_4_U119  ( .A(N151), .ZN(_add_0_root_add_136_4_n44 ) );
NOR2_X2 _add_0_root_add_136_4_U118  ( .A1(_add_0_root_add_136_4_n157 ), .A2(_add_0_root_add_136_4_n158 ), .ZN(_add_0_root_add_136_4_n156 ) );
NOR2_X4 _add_0_root_add_136_4_U117  ( .A1(_add_0_root_add_136_4_n282 ), .A2(_add_0_root_add_136_4_n88 ), .ZN(_add_0_root_add_136_4_n294 ) );
INV_X2 _add_0_root_add_136_4_U116  ( .A(_add_0_root_add_136_4_n108 ), .ZN(_add_0_root_add_136_4_n102 ) );
INV_X2 _add_0_root_add_136_4_U115  ( .A(_add_0_root_add_136_4_n399 ), .ZN(_add_0_root_add_136_4_n390 ) );
INV_X4 _add_0_root_add_136_4_U114  ( .A(_add_0_root_add_136_4_n269 ), .ZN(_add_0_root_add_136_4_n284 ) );
INV_X2 _add_0_root_add_136_4_U113  ( .A(_add_0_root_add_136_4_n25 ), .ZN(_add_0_root_add_136_4_n26 ) );
INV_X1 _add_0_root_add_136_4_U112  ( .A(_add_0_root_add_136_4_n18 ), .ZN(_add_0_root_add_136_4_n25 ) );
INV_X4 _add_0_root_add_136_4_U111  ( .A(_add_0_root_add_136_4_n24 ), .ZN(_add_0_root_add_136_4_n307 ) );
NOR2_X4 _add_0_root_add_136_4_U110  ( .A1(N146), .A2(N114), .ZN(_add_0_root_add_136_4_n24 ) );
NAND2_X1 _add_0_root_add_136_4_U109  ( .A1(_add_0_root_add_136_4_n81 ), .A2(_add_0_root_add_136_4_n372 ), .ZN(_add_0_root_add_136_4_n365 ) );
NOR2_X1 _add_0_root_add_136_4_U108  ( .A1(_add_0_root_add_136_4_n282 ), .A2(_add_0_root_add_136_4_n87 ), .ZN(_add_0_root_add_136_4_n300 ) );
NAND2_X2 _add_0_root_add_136_4_U107  ( .A1(_add_0_root_add_136_4_n329 ),.A2(_add_0_root_add_136_4_n339 ), .ZN(_add_0_root_add_136_4_n338 ) );
NAND2_X2 _add_0_root_add_136_4_U106  ( .A1(_add_0_root_add_136_4_n419 ),.A2(_add_0_root_add_136_4_n96 ), .ZN(_add_0_root_add_136_4_n418 ) );
INV_X8 _add_0_root_add_136_4_U105  ( .A(_add_0_root_add_136_4_n144 ), .ZN(_add_0_root_add_136_4_n23 ) );
NAND2_X2 _add_0_root_add_136_4_U104  ( .A1(_add_0_root_add_136_4_n40 ), .A2(_add_0_root_add_136_4_n42 ), .ZN(_add_0_root_add_136_4_n56 ) );
INV_X1 _add_0_root_add_136_4_U103  ( .A(_add_0_root_add_136_4_n294 ), .ZN(_add_0_root_add_136_4_n293 ) );
NAND2_X2 _add_0_root_add_136_4_U102  ( .A1(N146), .A2(N114), .ZN(_add_0_root_add_136_4_n314 ) );
NOR2_X2 _add_0_root_add_136_4_U101  ( .A1(N141), .A2(N109), .ZN(_add_0_root_add_136_4_n376 ) );
NAND2_X2 _add_0_root_add_136_4_U100  ( .A1(N141), .A2(N109), .ZN(_add_0_root_add_136_4_n378 ) );
XNOR2_X1 _add_0_root_add_136_4_U99  ( .A(_add_0_root_add_136_4_n379 ), .B(_add_0_root_add_136_4_n387 ), .ZN(next_A[12]) );
INV_X1 _add_0_root_add_136_4_U98  ( .A(_add_0_root_add_136_4_n233 ), .ZN(_add_0_root_add_136_4_n22 ) );
INV_X4 _add_0_root_add_136_4_U97  ( .A(_add_0_root_add_136_4_n243 ), .ZN(_add_0_root_add_136_4_n21 ) );
INV_X4 _add_0_root_add_136_4_U96  ( .A(_add_0_root_add_136_4_n342 ), .ZN(_add_0_root_add_136_4_n30 ) );
INV_X1 _add_0_root_add_136_4_U95  ( .A(_add_0_root_add_136_4_n30 ), .ZN(_add_0_root_add_136_4_n20 ) );
NAND2_X2 _add_0_root_add_136_4_U94  ( .A1(_add_0_root_add_136_4_n309 ), .A2(_add_0_root_add_136_4_n20 ), .ZN(_add_0_root_add_136_4_n330 ) );
NOR2_X2 _add_0_root_add_136_4_U93  ( .A1(N131), .A2(N99), .ZN(_add_0_root_add_136_4_n131 ) );
NOR2_X4 _add_0_root_add_136_4_U92  ( .A1(_add_0_root_add_136_4_n263 ), .A2(_add_0_root_add_136_4_n26 ), .ZN(_add_0_root_add_136_4_n261 ) );
INV_X2 _add_0_root_add_136_4_U91  ( .A(_add_0_root_add_136_4_n385 ), .ZN(_add_0_root_add_136_4_n384 ) );
NAND3_X2 _add_0_root_add_136_4_U90  ( .A1(_add_0_root_add_136_4_n308 ), .A2(_add_0_root_add_136_4_n309 ), .A3(_add_0_root_add_136_4_n304 ), .ZN(_add_0_root_add_136_4_n165 ) );
INV_X4 _add_0_root_add_136_4_U89  ( .A(_add_0_root_add_136_4_n242 ), .ZN(_add_0_root_add_136_4_n19 ) );
CLKBUF_X2 _add_0_root_add_136_4_U88  ( .A(_add_0_root_add_136_4_n186 ), .Z(_add_0_root_add_136_4_n48 ) );
NAND2_X4 _add_0_root_add_136_4_U87  ( .A1(_add_0_root_add_136_4_n45 ), .A2(N119), .ZN(_add_0_root_add_136_4_n265 ) );
NAND2_X4 _add_0_root_add_136_4_U86  ( .A1(_add_0_root_add_136_4_n264 ), .A2(_add_0_root_add_136_4_n265 ), .ZN(_add_0_root_add_136_4_n18 ) );
INV_X1 _add_0_root_add_136_4_U85  ( .A(_add_0_root_add_136_4_n304 ), .ZN(_add_0_root_add_136_4_n16 ) );
NOR2_X2 _add_0_root_add_136_4_U84  ( .A1(_add_0_root_add_136_4_n374 ), .A2(_add_0_root_add_136_4_n371 ), .ZN(_add_0_root_add_136_4_n373 ) );
INV_X1 _add_0_root_add_136_4_U83  ( .A(_add_0_root_add_136_4_n51 ), .ZN(_add_0_root_add_136_4_n285 ) );
NAND3_X2 _add_0_root_add_136_4_U82  ( .A1(_add_0_root_add_136_4_n211 ), .A2(_add_0_root_add_136_4_n210 ), .A3(_add_0_root_add_136_4_n21 ), .ZN(_add_0_root_add_136_4_n228 ) );
CLKBUF_X2 _add_0_root_add_136_4_U81  ( .A(_add_0_root_add_136_4_n34 ), .Z(_add_0_root_add_136_4_n15 ) );
NOR2_X2 _add_0_root_add_136_4_U80  ( .A1(_add_0_root_add_136_4_n205 ), .A2(_add_0_root_add_136_4_n206 ), .ZN(_add_0_root_add_136_4_n201 ) );
NAND2_X1 _add_0_root_add_136_4_U79  ( .A1(_add_0_root_add_136_4_n200 ), .A2(_add_0_root_add_136_4_n214 ), .ZN(_add_0_root_add_136_4_n218 ) );
NAND2_X2 _add_0_root_add_136_4_U78  ( .A1(_add_0_root_add_136_4_n395 ), .A2(_add_0_root_add_136_4_n396 ), .ZN(_add_0_root_add_136_4_n394 ) );
NAND2_X4 _add_0_root_add_136_4_U77  ( .A1(_add_0_root_add_136_4_n294 ), .A2(_add_0_root_add_136_4_n281 ), .ZN(_add_0_root_add_136_4_n280 ) );
OR2_X2 _add_0_root_add_136_4_U76  ( .A1(_add_0_root_add_136_4_n431 ), .A2(_add_0_root_add_136_4_n432 ), .ZN(_add_0_root_add_136_4_n14 ) );
AND2_X2 _add_0_root_add_136_4_U75  ( .A1(_add_0_root_add_136_4_n147 ), .A2(_add_0_root_add_136_4_n146 ), .ZN(_add_0_root_add_136_4_n13 ) );
OR2_X4 _add_0_root_add_136_4_U74  ( .A1(_add_0_root_add_136_4_n256 ), .A2(_add_0_root_add_136_4_n354 ), .ZN(_add_0_root_add_136_4_n12 ) );
OR2_X4 _add_0_root_add_136_4_U73  ( .A1(_add_0_root_add_136_4_n212 ), .A2(_add_0_root_add_136_4_n225 ), .ZN(_add_0_root_add_136_4_n11 ) );
AND2_X2 _add_0_root_add_136_4_U72  ( .A1(N132), .A2(N100), .ZN(_add_0_root_add_136_4_n10 ) );
AND2_X2 _add_0_root_add_136_4_U71  ( .A1(N129), .A2(N97), .ZN(_add_0_root_add_136_4_n9 ) );
INV_X2 _add_0_root_add_136_4_U70  ( .A(N150), .ZN(_add_0_root_add_136_4_n288 ) );
NAND2_X4 _add_0_root_add_136_4_U69  ( .A1(N150), .A2(N118), .ZN(_add_0_root_add_136_4_n277 ) );
NAND3_X2 _add_0_root_add_136_4_U68  ( .A1(_add_0_root_add_136_4_n21 ), .A2(_add_0_root_add_136_4_n210 ), .A3(_add_0_root_add_136_4_n211 ), .ZN(_add_0_root_add_136_4_n209 ) );
NOR2_X4 _add_0_root_add_136_4_U67  ( .A1(_add_0_root_add_136_4_n341 ), .A2(_add_0_root_add_136_4_n33 ), .ZN(_add_0_root_add_136_4_n312 ) );
NAND2_X4 _add_0_root_add_136_4_U66  ( .A1(_add_0_root_add_136_4_n221 ), .A2(_add_0_root_add_136_4_n222 ), .ZN(_add_0_root_add_136_4_n61 ) );
INV_X8 _add_0_root_add_136_4_U65  ( .A(_add_0_root_add_136_4_n7 ), .ZN(_add_0_root_add_136_4_n91 ) );
INV_X4 _add_0_root_add_136_4_U64  ( .A(_add_0_root_add_136_4_n211 ), .ZN(_add_0_root_add_136_4_n238 ) );
NAND2_X1 _add_0_root_add_136_4_U63  ( .A1(_add_0_root_add_136_4_n295 ), .A2(_add_0_root_add_136_4_n8 ), .ZN(_add_0_root_add_136_4_n278 ) );
NAND2_X4 _add_0_root_add_136_4_U62  ( .A1(_add_0_root_add_136_4_n59 ), .A2(_add_0_root_add_136_4_n60 ), .ZN(_add_0_root_add_136_4_n62 ) );
AND2_X2 _add_0_root_add_136_4_U61  ( .A1(N149), .A2(N117), .ZN(_add_0_root_add_136_4_n51 ) );
NOR2_X2 _add_0_root_add_136_4_U60  ( .A1(_add_0_root_add_136_4_n318 ), .A2(_add_0_root_add_136_4_n361 ), .ZN(_add_0_root_add_136_4_n340 ) );
NOR2_X2 _add_0_root_add_136_4_U59  ( .A1(_add_0_root_add_136_4_n5 ), .A2(_add_0_root_add_136_4_n160 ), .ZN(_add_0_root_add_136_4_n262 ) );
NOR2_X2 _add_0_root_add_136_4_U58  ( .A1(_add_0_root_add_136_4_n268 ), .A2(_add_0_root_add_136_4_n270 ), .ZN(_add_0_root_add_136_4_n287 ) );
NOR2_X1 _add_0_root_add_136_4_U57  ( .A1(_add_0_root_add_136_4_n130 ), .A2(_add_0_root_add_136_4_n350 ), .ZN(_add_0_root_add_136_4_n349 ) );
INV_X8 _add_0_root_add_136_4_U56  ( .A(_add_0_root_add_136_4_n165 ), .ZN(_add_0_root_add_136_4_n242 ) );
AND3_X4 _add_0_root_add_136_4_U55  ( .A1(_add_0_root_add_136_4_n164 ), .A2(_add_0_root_add_136_4_n49 ), .A3(_add_0_root_add_136_4_n6 ), .ZN(_add_0_root_add_136_4_n75 ) );
INV_X8 _add_0_root_add_136_4_U54  ( .A(_add_0_root_add_136_4_n184 ), .ZN(_add_0_root_add_136_4_n144 ) );
NOR2_X4 _add_0_root_add_136_4_U53  ( .A1(_add_0_root_add_136_4_n272 ), .A2(_add_0_root_add_136_4_n295 ), .ZN(_add_0_root_add_136_4_n292 ) );
INV_X8 _add_0_root_add_136_4_U52  ( .A(_add_0_root_add_136_4_n172 ), .ZN(_add_0_root_add_136_4_n303 ) );
NAND2_X4 _add_0_root_add_136_4_U51  ( .A1(_add_0_root_add_136_4_n18 ), .A2(_add_0_root_add_136_4_n239 ), .ZN(_add_0_root_add_136_4_n211 ) );
INV_X8 _add_0_root_add_136_4_U50  ( .A(_add_0_root_add_136_4_n142 ), .ZN(_add_0_root_add_136_4_n243 ) );
NOR2_X4 _add_0_root_add_136_4_U49  ( .A1(N153), .A2(N121), .ZN(_add_0_root_add_136_4_n212 ) );
NAND2_X4 _add_0_root_add_136_4_U48  ( .A1(N136), .A2(N104), .ZN(_add_0_root_add_136_4_n107 ) );
NOR2_X4 _add_0_root_add_136_4_U47  ( .A1(N102), .A2(N134), .ZN(_add_0_root_add_136_4_n431 ) );
NOR2_X2 _add_0_root_add_136_4_U46  ( .A1(_add_0_root_add_136_4_n84 ), .A2(_add_0_root_add_136_4_n112 ), .ZN(_add_0_root_add_136_4_n113 ) );
NOR2_X4 _add_0_root_add_136_4_U45  ( .A1(N101), .A2(N133), .ZN(_add_0_root_add_136_4_n435 ) );
NOR2_X4 _add_0_root_add_136_4_U44  ( .A1(N98), .A2(N130), .ZN(_add_0_root_add_136_4_n133 ) );
NAND2_X4 _add_0_root_add_136_4_U43  ( .A1(N128), .A2(N96), .ZN(_add_0_root_add_136_4_n258 ) );
NAND2_X2 _add_0_root_add_136_4_U42  ( .A1(_add_0_root_add_136_4_n71 ), .A2(_add_0_root_add_136_4_n377 ), .ZN(_add_0_root_add_136_4_n383 ) );
NAND2_X2 _add_0_root_add_136_4_U41  ( .A1(_add_0_root_add_136_4_n364 ), .A2(_add_0_root_add_136_4_n344 ), .ZN(_add_0_root_add_136_4_n362 ) );
NAND2_X2 _add_0_root_add_136_4_U40  ( .A1(_add_0_root_add_136_4_n302 ), .A2(_add_0_root_add_136_4_n296 ), .ZN(_add_0_root_add_136_4_n301 ) );
INV_X4 _add_0_root_add_136_4_U39  ( .A(_add_0_root_add_136_4_n301 ), .ZN(_add_0_root_add_136_4_n299 ) );
INV_X4 _add_0_root_add_136_4_U38  ( .A(_add_0_root_add_136_4_n313 ), .ZN(_add_0_root_add_136_4_n245 ) );
INV_X4 _add_0_root_add_136_4_U37  ( .A(_add_0_root_add_136_4_n372 ), .ZN(_add_0_root_add_136_4_n371 ) );
NAND2_X2 _add_0_root_add_136_4_U36  ( .A1(_add_0_root_add_136_4_n284 ), .A2(_add_0_root_add_136_4_n285 ), .ZN(_add_0_root_add_136_4_n283 ) );
NAND2_X2 _add_0_root_add_136_4_U35  ( .A1(_add_0_root_add_136_4_n375 ), .A2(_add_0_root_add_136_4_n356 ), .ZN(_add_0_root_add_136_4_n372 ) );
INV_X8 _add_0_root_add_136_4_U34  ( .A(_add_0_root_add_136_4_n273 ), .ZN(_add_0_root_add_136_4_n305 ) );
NOR2_X4 _add_0_root_add_136_4_U33  ( .A1(_add_0_root_add_136_4_n242 ), .A2(_add_0_root_add_136_4_n305 ), .ZN(_add_0_root_add_136_4_n302 ) );
AND2_X2 _add_0_root_add_136_4_U32  ( .A1(N135), .A2(N103), .ZN(_add_0_root_add_136_4_n85 ) );
NAND3_X2 _add_0_root_add_136_4_U31  ( .A1(_add_0_root_add_136_4_n96 ), .A2(_add_0_root_add_136_4_n107 ), .A3(_add_0_root_add_136_4_n108 ), .ZN(_add_0_root_add_136_4_n417 ) );
NOR2_X2 _add_0_root_add_136_4_U30  ( .A1(_add_0_root_add_136_4_n292 ), .A2(_add_0_root_add_136_4_n271 ), .ZN(_add_0_root_add_136_4_n263 ) );
NAND4_X1 _add_0_root_add_136_4_U29  ( .A1(_add_0_root_add_136_4_n140 ), .A2(_add_0_root_add_136_4_n141 ), .A3(_add_0_root_add_136_4_n50 ), .A4(_add_0_root_add_136_4_n243 ), .ZN(_add_0_root_add_136_4_n139 ) );
NOR2_X4 _add_0_root_add_136_4_U28  ( .A1(_add_0_root_add_136_4_n183 ), .A2(_add_0_root_add_136_4_n182 ), .ZN(_add_0_root_add_136_4_n426 ) );
NAND2_X4 _add_0_root_add_136_4_U27  ( .A1(_add_0_root_add_136_4_n426 ), .A2(_add_0_root_add_136_4_n427 ), .ZN(_add_0_root_add_136_4_n425 ) );
NOR2_X4 _add_0_root_add_136_4_U26  ( .A1(N135), .A2(N103), .ZN(_add_0_root_add_136_4_n34 ) );
INV_X4 _add_0_root_add_136_4_U25  ( .A(_add_0_root_add_136_4_n44 ), .ZN(_add_0_root_add_136_4_n45 ) );
NOR2_X4 _add_0_root_add_136_4_U24  ( .A1(N97), .A2(N129), .ZN(_add_0_root_add_136_4_n182 ) );
NAND2_X1 _add_0_root_add_136_4_U23  ( .A1(N129), .A2(N97), .ZN(_add_0_root_add_136_4_n428 ) );
NOR2_X4 _add_0_root_add_136_4_U22  ( .A1(_add_0_root_add_136_4_n408 ), .A2(_add_0_root_add_136_4_n409 ), .ZN(_add_0_root_add_136_4_n407 ) );
NOR2_X2 _add_0_root_add_136_4_U21  ( .A1(_add_0_root_add_136_4_n386 ), .A2(_add_0_root_add_136_4_n376 ), .ZN(_add_0_root_add_136_4_n385 ) );
OR2_X2 _add_0_root_add_136_4_U20  ( .A1(_add_0_root_add_136_4_n376 ), .A2(_add_0_root_add_136_4_n380 ), .ZN(_add_0_root_add_136_4_n81 ) );
BUF_X8 _add_0_root_add_136_4_U19  ( .A(_add_0_root_add_136_4_n250 ), .Z(_add_0_root_add_136_4_n8 ) );
NOR2_X1 _add_0_root_add_136_4_U18  ( .A1(N106), .A2(_add_0_root_add_136_4_n37 ), .ZN(_add_0_root_add_136_4_n414 ) );
NOR2_X4 _add_0_root_add_136_4_U17  ( .A1(_add_0_root_add_136_4_n207 ), .A2(_add_0_root_add_136_4_n208 ), .ZN(_add_0_root_add_136_4_n198 ) );
NOR2_X4 _add_0_root_add_136_4_U16  ( .A1(_add_0_root_add_136_4_n198 ), .A2(_add_0_root_add_136_4_n196 ), .ZN(_add_0_root_add_136_4_n197 ) );
INV_X2 _add_0_root_add_136_4_U15  ( .A(_add_0_root_add_136_4_n389 ), .ZN(_add_0_root_add_136_4_n17 ) );
INV_X4 _add_0_root_add_136_4_U14  ( .A(_add_0_root_add_136_4_n389 ), .ZN(_add_0_root_add_136_4_n7 ) );
NAND2_X4 _add_0_root_add_136_4_U13  ( .A1(_add_0_root_add_136_4_n245 ), .A2(_add_0_root_add_136_4_n164 ), .ZN(_add_0_root_add_136_4_n244 ) );
NAND3_X2 _add_0_root_add_136_4_U12  ( .A1(_add_0_root_add_136_4_n308 ), .A2(_add_0_root_add_136_4_n309 ), .A3(_add_0_root_add_136_4_n304 ), .ZN(_add_0_root_add_136_4_n6 ) );
NAND2_X2 _add_0_root_add_136_4_U11  ( .A1(_add_0_root_add_136_4_n231 ), .A2(_add_0_root_add_136_4_n244 ), .ZN(_add_0_root_add_136_4_n216 ) );
BUF_X8 _add_0_root_add_136_4_U10  ( .A(N152), .Z(_add_0_root_add_136_4_n52 ));
INV_X8 _add_0_root_add_136_4_U9  ( .A(_add_0_root_add_136_4_n5 ), .ZN(_add_0_root_add_136_4_n239 ) );
NOR2_X4 _add_0_root_add_136_4_U8  ( .A1(N152), .A2(N120), .ZN(_add_0_root_add_136_4_n5 ) );
INV_X1 _add_0_root_add_136_4_U7  ( .A(_add_0_root_add_136_4_n303 ), .ZN(_add_0_root_add_136_4_n4 ) );
NAND2_X4 _add_0_root_add_136_4_U6  ( .A1(_add_0_root_add_136_4_n381 ), .A2(_add_0_root_add_136_4_n382 ), .ZN(_add_0_root_add_136_4_n346 ) );
INV_X1 _add_0_root_add_136_4_U5  ( .A(_add_0_root_add_136_4_n358 ), .ZN(_add_0_root_add_136_4_n3 ) );
NOR2_X4 _add_0_root_add_136_4_U4  ( .A1(_add_0_root_add_136_4_n290 ), .A2(_add_0_root_add_136_4_n283 ), .ZN(_add_0_root_add_136_4_n286 ) );
INV_X4 _add_0_root_add_136_4_U3  ( .A(_add_0_root_add_136_4_n1 ), .ZN(_add_0_root_add_136_4_n2 ) );
INV_X1 _add_0_root_add_136_4_U2  ( .A(_add_0_root_add_136_4_n144 ), .ZN(_add_0_root_add_136_4_n1 ) );
endmodule
