
module sha1_exec ( clk, reset, start, data_in, load_in, cv, use_prev_cv, busy, 
        out_valid, cv_next );
  input [31:0] data_in;
  input [159:0] cv;
  output [159:0] cv_next;
  input clk, reset, start, load_in, use_prev_cv;
  output busy, out_valid;
  wire   N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,
         N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, n4654, n4655, n4656, n4658, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6117, n6118, n6139, n6140, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6569,
         n6570, n6571, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6856, n6859, n6862, n6865, n6868, n6871, n6874, n6877,
         n6880, n6883, n6884, n6885, n6886, n6889, n6892, n6895, n6898, n6901,
         n6904, n6907, n6910, n6913, n6916, n6917, n6918, n6919, n6922, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, \sha1_round/n825 ,
         \sha1_round/n824 , \sha1_round/n823 , \sha1_round/n822 ,
         \sha1_round/n821 , \sha1_round/n820 , \sha1_round/n819 ,
         \sha1_round/n818 , \sha1_round/n817 , \sha1_round/n816 ,
         \sha1_round/n815 , \sha1_round/n814 , \sha1_round/n813 ,
         \sha1_round/n812 , \sha1_round/n811 , \sha1_round/n810 ,
         \sha1_round/n809 , \sha1_round/n808 , \sha1_round/n807 ,
         \sha1_round/n806 , \sha1_round/n805 , \sha1_round/n804 ,
         \sha1_round/n803 , \sha1_round/n802 , \sha1_round/n801 ,
         \sha1_round/n800 , \sha1_round/n799 , \sha1_round/n798 ,
         \sha1_round/n797 , \sha1_round/n796 , \sha1_round/n795 ,
         \sha1_round/n794 , \sha1_round/n793 , \sha1_round/n792 ,
         \sha1_round/n791 , \sha1_round/n790 , \sha1_round/n789 ,
         \sha1_round/n788 , \sha1_round/n787 , \sha1_round/n786 ,
         \sha1_round/n785 , \sha1_round/n784 , \sha1_round/n783 ,
         \sha1_round/n782 , \sha1_round/n781 , \sha1_round/n780 ,
         \sha1_round/n779 , \sha1_round/n778 , \sha1_round/n777 ,
         \sha1_round/n776 , \sha1_round/n775 , \sha1_round/n774 ,
         \sha1_round/n773 , \sha1_round/n772 , \sha1_round/n771 ,
         \sha1_round/n770 , \sha1_round/n769 , \sha1_round/n768 ,
         \sha1_round/n767 , \sha1_round/n766 , \sha1_round/n765 ,
         \sha1_round/n764 , \sha1_round/n763 , \sha1_round/n762 ,
         \sha1_round/n761 , \sha1_round/n760 , \sha1_round/n759 ,
         \sha1_round/n758 , \sha1_round/n757 , \sha1_round/n756 ,
         \sha1_round/n755 , \sha1_round/n754 , \sha1_round/n753 ,
         \sha1_round/n752 , \sha1_round/n751 , \sha1_round/n750 ,
         \sha1_round/n749 , \sha1_round/n748 , \sha1_round/n747 ,
         \sha1_round/n746 , \sha1_round/n745 , \sha1_round/n744 ,
         \sha1_round/n743 , \sha1_round/n742 , \sha1_round/n741 ,
         \sha1_round/n740 , \sha1_round/n739 , \sha1_round/n738 ,
         \sha1_round/n737 , \sha1_round/n736 , \sha1_round/n735 ,
         \sha1_round/n734 , \sha1_round/n733 , \sha1_round/n732 ,
         \sha1_round/n731 , \sha1_round/n730 , \sha1_round/n729 ,
         \sha1_round/n728 , \sha1_round/n727 , \sha1_round/n726 ,
         \sha1_round/n725 , \sha1_round/n724 , \sha1_round/n723 ,
         \sha1_round/n722 , \sha1_round/n721 , \sha1_round/n720 ,
         \sha1_round/n719 , \sha1_round/n718 , \sha1_round/n717 ,
         \sha1_round/n716 , \sha1_round/n715 , \sha1_round/n714 ,
         \sha1_round/n713 , \sha1_round/n712 , \sha1_round/n711 ,
         \sha1_round/n710 , \sha1_round/n709 , \sha1_round/n708 ,
         \sha1_round/n707 , \sha1_round/n706 , \sha1_round/n705 ,
         \sha1_round/n704 , \sha1_round/n703 , \sha1_round/n702 ,
         \sha1_round/n701 , \sha1_round/n700 , \sha1_round/n699 ,
         \sha1_round/n698 , \sha1_round/n697 , \sha1_round/n696 ,
         \sha1_round/n695 , \sha1_round/n694 , \sha1_round/n693 ,
         \sha1_round/n692 , \sha1_round/n691 , \sha1_round/n690 ,
         \sha1_round/n689 , \sha1_round/n688 , \sha1_round/n687 ,
         \sha1_round/n686 , \sha1_round/n685 , \sha1_round/n684 ,
         \sha1_round/n683 , \sha1_round/n682 , \sha1_round/n681 ,
         \sha1_round/n680 , \sha1_round/n679 , \sha1_round/n678 ,
         \sha1_round/n677 , \sha1_round/n676 , \sha1_round/n675 ,
         \sha1_round/n674 , \sha1_round/n673 , \sha1_round/n672 ,
         \sha1_round/n671 , \sha1_round/n670 , \sha1_round/n669 ,
         \sha1_round/n668 , \sha1_round/n667 , \sha1_round/n666 ,
         \sha1_round/n665 , \sha1_round/n664 , \sha1_round/n663 ,
         \sha1_round/n662 , \sha1_round/n661 , \sha1_round/n660 ,
         \sha1_round/n659 , \sha1_round/n658 , \sha1_round/n657 ,
         \sha1_round/n656 , \sha1_round/n655 , \sha1_round/n654 ,
         \sha1_round/n653 , \sha1_round/n652 , \sha1_round/n651 ,
         \sha1_round/n650 , \sha1_round/n649 , \sha1_round/n648 ,
         \sha1_round/n647 , \sha1_round/n646 , \sha1_round/n645 ,
         \sha1_round/n644 , \sha1_round/n643 , \sha1_round/n642 ,
         \sha1_round/n641 , \sha1_round/n640 , \sha1_round/n639 ,
         \sha1_round/n638 , \sha1_round/n637 , \sha1_round/n636 ,
         \sha1_round/n635 , \sha1_round/n634 , \sha1_round/n633 ,
         \sha1_round/n632 , \sha1_round/n631 , \sha1_round/n630 ,
         \sha1_round/n629 , \sha1_round/n628 , \sha1_round/n627 ,
         \sha1_round/n626 , \sha1_round/n625 , \sha1_round/n624 ,
         \sha1_round/n623 , \sha1_round/n622 , \sha1_round/n621 ,
         \sha1_round/n620 , \sha1_round/n619 , \sha1_round/n618 ,
         \sha1_round/n617 , \sha1_round/n616 , \sha1_round/n615 ,
         \sha1_round/n614 , \sha1_round/n613 , \sha1_round/n612 ,
         \sha1_round/n611 , \sha1_round/n610 , \sha1_round/n609 ,
         \sha1_round/n608 , \sha1_round/n607 , \sha1_round/n606 ,
         \sha1_round/n605 , \sha1_round/n604 , \sha1_round/n603 ,
         \sha1_round/n602 , \sha1_round/n601 , \sha1_round/n600 ,
         \sha1_round/n599 , \sha1_round/n598 , \sha1_round/n597 ,
         \sha1_round/n596 , \sha1_round/n595 , \sha1_round/n594 ,
         \sha1_round/n593 , \sha1_round/n592 , \sha1_round/n591 ,
         \sha1_round/n590 , \sha1_round/n589 , \sha1_round/n588 ,
         \sha1_round/n587 , \sha1_round/n586 , \sha1_round/n585 ,
         \sha1_round/n584 , \sha1_round/n583 , \sha1_round/n582 ,
         \sha1_round/n581 , \sha1_round/n580 , \sha1_round/n579 ,
         \sha1_round/n578 , \sha1_round/n577 , \sha1_round/n576 ,
         \sha1_round/n575 , \sha1_round/n574 , \sha1_round/n573 ,
         \sha1_round/n572 , \sha1_round/n571 , \sha1_round/n570 ,
         \sha1_round/n569 , \sha1_round/n568 , \sha1_round/n567 ,
         \sha1_round/n566 , \sha1_round/n565 , \sha1_round/n564 ,
         \sha1_round/n563 , \sha1_round/n562 , \sha1_round/n561 ,
         \sha1_round/n560 , \sha1_round/n559 , \sha1_round/n558 ,
         \sha1_round/n557 , \sha1_round/n556 , \sha1_round/n555 ,
         \sha1_round/n554 , \sha1_round/n553 , \sha1_round/n552 ,
         \sha1_round/n551 , \sha1_round/n550 , \sha1_round/n549 ,
         \sha1_round/n548 , \sha1_round/n547 , \sha1_round/n546 ,
         \sha1_round/n545 , \sha1_round/n544 , \sha1_round/n543 ,
         \sha1_round/n542 , \sha1_round/n541 , \sha1_round/n540 ,
         \sha1_round/n539 , \sha1_round/n538 , \sha1_round/n537 ,
         \sha1_round/n536 , \sha1_round/n535 , \sha1_round/n534 ,
         \sha1_round/n533 , \sha1_round/n532 , \sha1_round/n531 ,
         \sha1_round/n530 , \sha1_round/n529 , \sha1_round/n528 ,
         \sha1_round/n527 , \sha1_round/n526 , \sha1_round/n525 ,
         \sha1_round/n524 , \sha1_round/n523 , \sha1_round/n522 ,
         \sha1_round/n521 , \sha1_round/n520 , \sha1_round/n519 ,
         \sha1_round/n518 , \sha1_round/n517 , \sha1_round/n516 ,
         \sha1_round/n515 , \sha1_round/n514 , \sha1_round/n513 ,
         \sha1_round/n512 , \sha1_round/n511 , \sha1_round/n510 ,
         \sha1_round/n509 , \sha1_round/n508 , \sha1_round/n380 ,
         \sha1_round/n379 , \sha1_round/n378 , \sha1_round/n377 ,
         \sha1_round/n376 , \sha1_round/n375 , \sha1_round/n374 ,
         \sha1_round/n373 , \sha1_round/n372 , \sha1_round/n371 ,
         \sha1_round/n370 , \sha1_round/n369 , \sha1_round/n368 ,
         \sha1_round/n367 , \sha1_round/n366 , \sha1_round/n365 ,
         \sha1_round/n364 , \sha1_round/n363 , \sha1_round/n362 ,
         \sha1_round/n361 , \sha1_round/n360 , \sha1_round/n359 ,
         \sha1_round/n358 , \sha1_round/n357 , \sha1_round/n356 ,
         \sha1_round/n355 , \sha1_round/n354 , \sha1_round/n353 ,
         \sha1_round/n352 , \sha1_round/n351 , \sha1_round/n350 ,
         \sha1_round/n349 , \sha1_round/n348 , \sha1_round/n3470 ,
         \sha1_round/n3460 , \sha1_round/n3450 , \sha1_round/n3440 ,
         \sha1_round/n3430 , \sha1_round/n3420 , \sha1_round/n3410 ,
         \sha1_round/n3400 , \sha1_round/n3390 , \sha1_round/n3380 ,
         \sha1_round/n3370 , \sha1_round/n3360 , \sha1_round/n3350 ,
         \sha1_round/n3340 , \sha1_round/n3330 , \sha1_round/n3320 ,
         \sha1_round/n3300 , \sha1_round/n3290 , \sha1_round/n3280 ,
         \sha1_round/n3270 , \sha1_round/n3260 , \sha1_round/n3250 ,
         \sha1_round/n3240 , \sha1_round/n3230 , \sha1_round/n3220 ,
         \sha1_round/n3210 , \sha1_round/n3200 , \sha1_round/n3190 ,
         \sha1_round/n3180 , \sha1_round/n3160 , \sha1_round/n3150 ,
         \sha1_round/n3140 , \sha1_round/n3130 , \sha1_round/n3120 ,
         \sha1_round/n3170 , \sha1_round/n168 , \sha1_round/n167 ,
         \sha1_round/n159 , \sha1_round/n158 , \sha1_round/n150 ,
         \sha1_round/n149 , \sha1_round/n141 , \sha1_round/n140 ,
         \sha1_round/n132 , \sha1_round/n131 , \sha1_round/n123 ,
         \sha1_round/n122 , \sha1_round/n114 , \sha1_round/n113 ,
         \sha1_round/n96 , \sha1_round/n95 , \sha1_round/n87 ,
         \sha1_round/n86 , \sha1_round/n2 , \sha1_round/N252 ,
         \sha1_round/N253 , \sha1_round/N254 , \sha1_round/N255 ,
         \sha1_round/N256 , \sha1_round/N257 , \sha1_round/N258 ,
         \sha1_round/N259 , \sha1_round/N260 , \sha1_round/N261 ,
         \sha1_round/N262 , \sha1_round/N263 , \sha1_round/N264 ,
         \sha1_round/N265 , \sha1_round/N266 , \sha1_round/N267 ,
         \sha1_round/N268 , \sha1_round/N269 , \sha1_round/N270 ,
         \sha1_round/N271 , \sha1_round/N272 , \sha1_round/N273 ,
         \sha1_round/N274 , \sha1_round/N275 , \sha1_round/N276 ,
         \sha1_round/N277 , \sha1_round/N278 , \sha1_round/N279 ,
         \sha1_round/N280 , \sha1_round/N281 , \sha1_round/N282 ,
         \sha1_round/N283 , \sha1_round/N284 , \sha1_round/N285 ,
         \sha1_round/N286 , \sha1_round/N287 , \sha1_round/N288 ,
         \sha1_round/N289 , \sha1_round/N290 , \sha1_round/N291 ,
         \sha1_round/N292 , \sha1_round/N293 , \sha1_round/N294 ,
         \sha1_round/N295 , \sha1_round/N296 , \sha1_round/N297 ,
         \sha1_round/N298 , \sha1_round/N299 , \sha1_round/N300 ,
         \sha1_round/N301 , \sha1_round/N302 , \sha1_round/N303 ,
         \sha1_round/N304 , \sha1_round/N305 , \sha1_round/N306 ,
         \sha1_round/N307 , \sha1_round/N308 , \sha1_round/N309 ,
         \sha1_round/N310 , \sha1_round/N311 , \sha1_round/N312 ,
         \sha1_round/N313 , \sha1_round/N314 , \sha1_round/N315 ,
         \sha1_round/N316 , \sha1_round/N317 , \sha1_round/N318 ,
         \sha1_round/N319 , \sha1_round/N320 , \sha1_round/N321 ,
         \sha1_round/N322 , \sha1_round/N323 , \sha1_round/N324 ,
         \sha1_round/N325 , \sha1_round/N326 , \sha1_round/N327 ,
         \sha1_round/N328 , \sha1_round/N329 , \sha1_round/N330 ,
         \sha1_round/N331 , \sha1_round/N332 , \sha1_round/N333 ,
         \sha1_round/N334 , \sha1_round/N335 , \sha1_round/N336 ,
         \sha1_round/N337 , \sha1_round/N338 , \sha1_round/N339 ,
         \sha1_round/N340 , \sha1_round/N341 , \sha1_round/N342 ,
         \sha1_round/N343 , \sha1_round/N344 , \sha1_round/N345 ,
         \sha1_round/N346 , \sha1_round/N347 , \sha1_round/k[3] ,
         \sha1_round/k[13] , \sha1_round/k[15] , \sha1_round/k_23 ,
         \sha1_round/k_26 , \sha1_round/k_27 , \sha1_round/k_30 ,
         \sha1_round/add_79_4/n345 , \sha1_round/add_79_4/n344 ,
         \sha1_round/add_79_4/n343 , \sha1_round/add_79_4/n342 ,
         \sha1_round/add_79_4/n341 , \sha1_round/add_79_4/n340 ,
         \sha1_round/add_79_4/n339 , \sha1_round/add_79_4/n338 ,
         \sha1_round/add_79_4/n337 , \sha1_round/add_79_4/n336 ,
         \sha1_round/add_79_4/n335 , \sha1_round/add_79_4/n334 ,
         \sha1_round/add_79_4/n333 , \sha1_round/add_79_4/n332 ,
         \sha1_round/add_79_4/n331 , \sha1_round/add_79_4/n330 ,
         \sha1_round/add_79_4/n329 , \sha1_round/add_79_4/n328 ,
         \sha1_round/add_79_4/n327 , \sha1_round/add_79_4/n326 ,
         \sha1_round/add_79_4/n325 , \sha1_round/add_79_4/n324 ,
         \sha1_round/add_79_4/n323 , \sha1_round/add_79_4/n322 ,
         \sha1_round/add_79_4/n321 , \sha1_round/add_79_4/n320 ,
         \sha1_round/add_79_4/n319 , \sha1_round/add_79_4/n318 ,
         \sha1_round/add_79_4/n317 , \sha1_round/add_79_4/n316 ,
         \sha1_round/add_79_4/n315 , \sha1_round/add_79_4/n314 ,
         \sha1_round/add_79_4/n313 , \sha1_round/add_79_4/n312 ,
         \sha1_round/add_79_4/n311 , \sha1_round/add_79_4/n310 ,
         \sha1_round/add_79_4/n309 , \sha1_round/add_79_4/n308 ,
         \sha1_round/add_79_4/n307 , \sha1_round/add_79_4/n306 ,
         \sha1_round/add_79_4/n305 , \sha1_round/add_79_4/n304 ,
         \sha1_round/add_79_4/n303 , \sha1_round/add_79_4/n302 ,
         \sha1_round/add_79_4/n301 , \sha1_round/add_79_4/n300 ,
         \sha1_round/add_79_4/n299 , \sha1_round/add_79_4/n298 ,
         \sha1_round/add_79_4/n297 , \sha1_round/add_79_4/n296 ,
         \sha1_round/add_79_4/n295 , \sha1_round/add_79_4/n294 ,
         \sha1_round/add_79_4/n293 , \sha1_round/add_79_4/n292 ,
         \sha1_round/add_79_4/n291 , \sha1_round/add_79_4/n290 ,
         \sha1_round/add_79_4/n289 , \sha1_round/add_79_4/n288 ,
         \sha1_round/add_79_4/n287 , \sha1_round/add_79_4/n286 ,
         \sha1_round/add_79_4/n285 , \sha1_round/add_79_4/n284 ,
         \sha1_round/add_79_4/n283 , \sha1_round/add_79_4/n282 ,
         \sha1_round/add_79_4/n281 , \sha1_round/add_79_4/n280 ,
         \sha1_round/add_79_4/n279 , \sha1_round/add_79_4/n278 ,
         \sha1_round/add_79_4/n277 , \sha1_round/add_79_4/n276 ,
         \sha1_round/add_79_4/n275 , \sha1_round/add_79_4/n274 ,
         \sha1_round/add_79_4/n273 , \sha1_round/add_79_4/n272 ,
         \sha1_round/add_79_4/n271 , \sha1_round/add_79_4/n270 ,
         \sha1_round/add_79_4/n269 , \sha1_round/add_79_4/n268 ,
         \sha1_round/add_79_4/n267 , \sha1_round/add_79_4/n266 ,
         \sha1_round/add_79_4/n265 , \sha1_round/add_79_4/n264 ,
         \sha1_round/add_79_4/n263 , \sha1_round/add_79_4/n262 ,
         \sha1_round/add_79_4/n261 , \sha1_round/add_79_4/n260 ,
         \sha1_round/add_79_4/n259 , \sha1_round/add_79_4/n258 ,
         \sha1_round/add_79_4/n257 , \sha1_round/add_79_4/n256 ,
         \sha1_round/add_79_4/n255 , \sha1_round/add_79_4/n254 ,
         \sha1_round/add_79_4/n253 , \sha1_round/add_79_4/n252 ,
         \sha1_round/add_79_4/n251 , \sha1_round/add_79_4/n250 ,
         \sha1_round/add_79_4/n249 , \sha1_round/add_79_4/n248 ,
         \sha1_round/add_79_4/n247 , \sha1_round/add_79_4/n246 ,
         \sha1_round/add_79_4/n245 , \sha1_round/add_79_4/n244 ,
         \sha1_round/add_79_4/n243 , \sha1_round/add_79_4/n242 ,
         \sha1_round/add_79_4/n241 , \sha1_round/add_79_4/n240 ,
         \sha1_round/add_79_4/n239 , \sha1_round/add_79_4/n238 ,
         \sha1_round/add_79_4/n237 , \sha1_round/add_79_4/n236 ,
         \sha1_round/add_79_4/n235 , \sha1_round/add_79_4/n234 ,
         \sha1_round/add_79_4/n233 , \sha1_round/add_79_4/n232 ,
         \sha1_round/add_79_4/n231 , \sha1_round/add_79_4/n230 ,
         \sha1_round/add_79_4/n229 , \sha1_round/add_79_4/n228 ,
         \sha1_round/add_79_4/n227 , \sha1_round/add_79_4/n226 ,
         \sha1_round/add_79_4/n225 , \sha1_round/add_79_4/n224 ,
         \sha1_round/add_79_4/n223 , \sha1_round/add_79_4/n222 ,
         \sha1_round/add_79_4/n221 , \sha1_round/add_79_4/n220 ,
         \sha1_round/add_79_4/n219 , \sha1_round/add_79_4/n218 ,
         \sha1_round/add_79_4/n217 , \sha1_round/add_79_4/n216 ,
         \sha1_round/add_79_4/n215 , \sha1_round/add_79_4/n214 ,
         \sha1_round/add_79_4/n213 , \sha1_round/add_79_4/n212 ,
         \sha1_round/add_79_4/n211 , \sha1_round/add_79_4/n210 ,
         \sha1_round/add_79_4/n209 , \sha1_round/add_79_4/n208 ,
         \sha1_round/add_79_4/n207 , \sha1_round/add_79_4/n206 ,
         \sha1_round/add_79_4/n205 , \sha1_round/add_79_4/n204 ,
         \sha1_round/add_79_4/n203 , \sha1_round/add_79_4/n202 ,
         \sha1_round/add_79_4/n201 , \sha1_round/add_79_4/n200 ,
         \sha1_round/add_79_4/n199 , \sha1_round/add_79_4/n198 ,
         \sha1_round/add_79_4/n197 , \sha1_round/add_79_4/n196 ,
         \sha1_round/add_79_4/n195 , \sha1_round/add_79_4/n194 ,
         \sha1_round/add_79_4/n193 , \sha1_round/add_79_4/n192 ,
         \sha1_round/add_79_4/n191 , \sha1_round/add_79_4/n190 ,
         \sha1_round/add_79_4/n189 , \sha1_round/add_79_4/n188 ,
         \sha1_round/add_79_4/n187 , \sha1_round/add_79_4/n186 ,
         \sha1_round/add_79_4/n185 , \sha1_round/add_79_4/n184 ,
         \sha1_round/add_79_4/n183 , \sha1_round/add_79_4/n182 ,
         \sha1_round/add_79_4/n181 , \sha1_round/add_79_4/n180 ,
         \sha1_round/add_79_4/n179 , \sha1_round/add_79_4/n178 ,
         \sha1_round/add_79_4/n177 , \sha1_round/add_79_4/n176 ,
         \sha1_round/add_79_4/n175 , \sha1_round/add_79_4/n174 ,
         \sha1_round/add_79_4/n173 , \sha1_round/add_79_4/n172 ,
         \sha1_round/add_79_4/n171 , \sha1_round/add_79_4/n170 ,
         \sha1_round/add_79_4/n169 , \sha1_round/add_79_4/n168 ,
         \sha1_round/add_79_4/n167 , \sha1_round/add_79_4/n166 ,
         \sha1_round/add_79_4/n165 , \sha1_round/add_79_4/n164 ,
         \sha1_round/add_79_4/n163 , \sha1_round/add_79_4/n162 ,
         \sha1_round/add_79_4/n161 , \sha1_round/add_79_4/n160 ,
         \sha1_round/add_79_4/n159 , \sha1_round/add_79_4/n158 ,
         \sha1_round/add_79_4/n157 , \sha1_round/add_79_4/n156 ,
         \sha1_round/add_79_4/n155 , \sha1_round/add_79_4/n154 ,
         \sha1_round/add_79_4/n153 , \sha1_round/add_79_4/n152 ,
         \sha1_round/add_79_4/n151 , \sha1_round/add_79_4/n150 ,
         \sha1_round/add_79_4/n149 , \sha1_round/add_79_4/n148 ,
         \sha1_round/add_79_4/n147 , \sha1_round/add_79_4/n146 ,
         \sha1_round/add_79_4/n145 , \sha1_round/add_79_4/n144 ,
         \sha1_round/add_79_4/n143 , \sha1_round/add_79_4/n142 ,
         \sha1_round/add_79_4/n141 , \sha1_round/add_79_4/n140 ,
         \sha1_round/add_79_4/n139 , \sha1_round/add_79_4/n138 ,
         \sha1_round/add_79_4/n137 , \sha1_round/add_79_4/n136 ,
         \sha1_round/add_79_4/n135 , \sha1_round/add_79_4/n134 ,
         \sha1_round/add_79_4/n133 , \sha1_round/add_79_4/n132 ,
         \sha1_round/add_79_4/n131 , \sha1_round/add_79_4/n130 ,
         \sha1_round/add_79_4/n129 , \sha1_round/add_79_4/n128 ,
         \sha1_round/add_79_4/n127 , \sha1_round/add_79_4/n126 ,
         \sha1_round/add_79_4/n125 , \sha1_round/add_79_4/n124 ,
         \sha1_round/add_79_4/n123 , \sha1_round/add_79_4/n122 ,
         \sha1_round/add_79_4/n121 , \sha1_round/add_79_4/n120 ,
         \sha1_round/add_79_4/n119 , \sha1_round/add_79_4/n118 ,
         \sha1_round/add_79_4/n117 , \sha1_round/add_79_4/n116 ,
         \sha1_round/add_79_4/n115 , \sha1_round/add_79_4/n114 ,
         \sha1_round/add_79_4/n113 , \sha1_round/add_79_4/n112 ,
         \sha1_round/add_79_4/n111 , \sha1_round/add_79_4/n110 ,
         \sha1_round/add_79_4/n109 , \sha1_round/add_79_4/n108 ,
         \sha1_round/add_79_4/n107 , \sha1_round/add_79_4/n106 ,
         \sha1_round/add_79_4/n105 , \sha1_round/add_79_4/n104 ,
         \sha1_round/add_79_4/n103 , \sha1_round/add_79_4/n102 ,
         \sha1_round/add_79_4/n101 , \sha1_round/add_79_4/n100 ,
         \sha1_round/add_79_4/n99 , \sha1_round/add_79_4/n98 ,
         \sha1_round/add_79_4/n97 , \sha1_round/add_79_4/n96 ,
         \sha1_round/add_79_4/n95 , \sha1_round/add_79_4/n94 ,
         \sha1_round/add_79_4/n93 , \sha1_round/add_79_4/n92 ,
         \sha1_round/add_79_4/n91 , \sha1_round/add_79_4/n90 ,
         \sha1_round/add_79_4/n89 , \sha1_round/add_79_4/n88 ,
         \sha1_round/add_79_4/n87 , \sha1_round/add_79_4/n86 ,
         \sha1_round/add_79_4/n85 , \sha1_round/add_79_4/n84 ,
         \sha1_round/add_79_4/n83 , \sha1_round/add_79_4/n82 ,
         \sha1_round/add_79_4/n81 , \sha1_round/add_79_4/n80 ,
         \sha1_round/add_79_4/n79 , \sha1_round/add_79_4/n78 ,
         \sha1_round/add_79_4/n77 , \sha1_round/add_79_4/n76 ,
         \sha1_round/add_79_4/n75 , \sha1_round/add_79_4/n74 ,
         \sha1_round/add_79_4/n73 , \sha1_round/add_79_4/n72 ,
         \sha1_round/add_79_4/n71 , \sha1_round/add_79_4/n70 ,
         \sha1_round/add_79_4/n69 , \sha1_round/add_79_4/n68 ,
         \sha1_round/add_79_4/n67 , \sha1_round/add_79_4/n66 ,
         \sha1_round/add_79_4/n65 , \sha1_round/add_79_4/n64 ,
         \sha1_round/add_79_4/n63 , \sha1_round/add_79_4/n62 ,
         \sha1_round/add_79_4/n61 , \sha1_round/add_79_4/n60 ,
         \sha1_round/add_79_4/n59 , \sha1_round/add_79_4/n58 ,
         \sha1_round/add_79_4/n57 , \sha1_round/add_79_4/n56 ,
         \sha1_round/add_79_4/n55 , \sha1_round/add_79_4/n54 ,
         \sha1_round/add_79_4/n53 , \sha1_round/add_79_4/n52 ,
         \sha1_round/add_79_4/n51 , \sha1_round/add_79_4/n50 ,
         \sha1_round/add_79_4/n49 , \sha1_round/add_79_4/n48 ,
         \sha1_round/add_79_4/n47 , \sha1_round/add_79_4/n46 ,
         \sha1_round/add_79_4/n45 , \sha1_round/add_79_4/n44 ,
         \sha1_round/add_79_4/n43 , \sha1_round/add_79_4/n42 ,
         \sha1_round/add_79_4/n41 , \sha1_round/add_79_4/n40 ,
         \sha1_round/add_79_4/n39 , \sha1_round/add_79_4/n38 ,
         \sha1_round/add_79_4/n37 , \sha1_round/add_79_4/n36 ,
         \sha1_round/add_79_4/n35 , \sha1_round/add_79_4/n34 ,
         \sha1_round/add_79_4/n33 , \sha1_round/add_79_4/n32 ,
         \sha1_round/add_79_4/n31 , \sha1_round/add_79_4/n30 ,
         \sha1_round/add_79_4/n29 , \sha1_round/add_79_4/n28 ,
         \sha1_round/add_79_4/n27 , \sha1_round/add_79_4/n26 ,
         \sha1_round/add_79_4/n25 , \sha1_round/add_79_4/n24 ,
         \sha1_round/add_79_4/n23 , \sha1_round/add_79_4/n22 ,
         \sha1_round/add_79_4/n21 , \sha1_round/add_79_4/n20 ,
         \sha1_round/add_79_4/n19 , \sha1_round/add_79_4/n18 ,
         \sha1_round/add_79_4/n17 , \sha1_round/add_79_4/n15 ,
         \sha1_round/add_79_4/n14 , \sha1_round/add_79_4/n13 ,
         \sha1_round/add_79_4/n12 , \sha1_round/add_79_4/n11 ,
         \sha1_round/add_79_4/n10 , \sha1_round/add_79_4/n9 ,
         \sha1_round/add_79_4/n8 , \sha1_round/add_79_4/n7 ,
         \sha1_round/add_79_4/n6 , \sha1_round/add_79_4/n5 ,
         \sha1_round/add_79_4/n4 , \sha1_round/add_79_4/n3 ,
         \sha1_round/add_79_4/n2 , \sha1_round/add_79_4/n1 ,
         \sha1_round/add_79_3/n387 , \sha1_round/add_79_3/n386 ,
         \sha1_round/add_79_3/n385 , \sha1_round/add_79_3/n384 ,
         \sha1_round/add_79_3/n383 , \sha1_round/add_79_3/n382 ,
         \sha1_round/add_79_3/n381 , \sha1_round/add_79_3/n380 ,
         \sha1_round/add_79_3/n379 , \sha1_round/add_79_3/n378 ,
         \sha1_round/add_79_3/n377 , \sha1_round/add_79_3/n376 ,
         \sha1_round/add_79_3/n375 , \sha1_round/add_79_3/n374 ,
         \sha1_round/add_79_3/n373 , \sha1_round/add_79_3/n372 ,
         \sha1_round/add_79_3/n371 , \sha1_round/add_79_3/n370 ,
         \sha1_round/add_79_3/n369 , \sha1_round/add_79_3/n368 ,
         \sha1_round/add_79_3/n367 , \sha1_round/add_79_3/n366 ,
         \sha1_round/add_79_3/n365 , \sha1_round/add_79_3/n364 ,
         \sha1_round/add_79_3/n363 , \sha1_round/add_79_3/n362 ,
         \sha1_round/add_79_3/n361 , \sha1_round/add_79_3/n360 ,
         \sha1_round/add_79_3/n359 , \sha1_round/add_79_3/n358 ,
         \sha1_round/add_79_3/n357 , \sha1_round/add_79_3/n356 ,
         \sha1_round/add_79_3/n355 , \sha1_round/add_79_3/n354 ,
         \sha1_round/add_79_3/n353 , \sha1_round/add_79_3/n352 ,
         \sha1_round/add_79_3/n351 , \sha1_round/add_79_3/n350 ,
         \sha1_round/add_79_3/n349 , \sha1_round/add_79_3/n348 ,
         \sha1_round/add_79_3/n347 , \sha1_round/add_79_3/n346 ,
         \sha1_round/add_79_3/n345 , \sha1_round/add_79_3/n344 ,
         \sha1_round/add_79_3/n343 , \sha1_round/add_79_3/n342 ,
         \sha1_round/add_79_3/n341 , \sha1_round/add_79_3/n340 ,
         \sha1_round/add_79_3/n339 , \sha1_round/add_79_3/n338 ,
         \sha1_round/add_79_3/n337 , \sha1_round/add_79_3/n336 ,
         \sha1_round/add_79_3/n335 , \sha1_round/add_79_3/n334 ,
         \sha1_round/add_79_3/n333 , \sha1_round/add_79_3/n332 ,
         \sha1_round/add_79_3/n331 , \sha1_round/add_79_3/n330 ,
         \sha1_round/add_79_3/n329 , \sha1_round/add_79_3/n328 ,
         \sha1_round/add_79_3/n327 , \sha1_round/add_79_3/n326 ,
         \sha1_round/add_79_3/n325 , \sha1_round/add_79_3/n324 ,
         \sha1_round/add_79_3/n323 , \sha1_round/add_79_3/n322 ,
         \sha1_round/add_79_3/n321 , \sha1_round/add_79_3/n320 ,
         \sha1_round/add_79_3/n319 , \sha1_round/add_79_3/n318 ,
         \sha1_round/add_79_3/n317 , \sha1_round/add_79_3/n316 ,
         \sha1_round/add_79_3/n315 , \sha1_round/add_79_3/n314 ,
         \sha1_round/add_79_3/n313 , \sha1_round/add_79_3/n312 ,
         \sha1_round/add_79_3/n311 , \sha1_round/add_79_3/n310 ,
         \sha1_round/add_79_3/n309 , \sha1_round/add_79_3/n308 ,
         \sha1_round/add_79_3/n307 , \sha1_round/add_79_3/n306 ,
         \sha1_round/add_79_3/n305 , \sha1_round/add_79_3/n304 ,
         \sha1_round/add_79_3/n303 , \sha1_round/add_79_3/n302 ,
         \sha1_round/add_79_3/n301 , \sha1_round/add_79_3/n300 ,
         \sha1_round/add_79_3/n299 , \sha1_round/add_79_3/n298 ,
         \sha1_round/add_79_3/n297 , \sha1_round/add_79_3/n296 ,
         \sha1_round/add_79_3/n295 , \sha1_round/add_79_3/n294 ,
         \sha1_round/add_79_3/n293 , \sha1_round/add_79_3/n292 ,
         \sha1_round/add_79_3/n291 , \sha1_round/add_79_3/n290 ,
         \sha1_round/add_79_3/n289 , \sha1_round/add_79_3/n288 ,
         \sha1_round/add_79_3/n287 , \sha1_round/add_79_3/n286 ,
         \sha1_round/add_79_3/n285 , \sha1_round/add_79_3/n284 ,
         \sha1_round/add_79_3/n283 , \sha1_round/add_79_3/n282 ,
         \sha1_round/add_79_3/n281 , \sha1_round/add_79_3/n280 ,
         \sha1_round/add_79_3/n279 , \sha1_round/add_79_3/n278 ,
         \sha1_round/add_79_3/n277 , \sha1_round/add_79_3/n276 ,
         \sha1_round/add_79_3/n275 , \sha1_round/add_79_3/n274 ,
         \sha1_round/add_79_3/n273 , \sha1_round/add_79_3/n272 ,
         \sha1_round/add_79_3/n271 , \sha1_round/add_79_3/n270 ,
         \sha1_round/add_79_3/n269 , \sha1_round/add_79_3/n268 ,
         \sha1_round/add_79_3/n267 , \sha1_round/add_79_3/n266 ,
         \sha1_round/add_79_3/n265 , \sha1_round/add_79_3/n264 ,
         \sha1_round/add_79_3/n263 , \sha1_round/add_79_3/n262 ,
         \sha1_round/add_79_3/n261 , \sha1_round/add_79_3/n260 ,
         \sha1_round/add_79_3/n259 , \sha1_round/add_79_3/n258 ,
         \sha1_round/add_79_3/n257 , \sha1_round/add_79_3/n256 ,
         \sha1_round/add_79_3/n255 , \sha1_round/add_79_3/n254 ,
         \sha1_round/add_79_3/n253 , \sha1_round/add_79_3/n252 ,
         \sha1_round/add_79_3/n251 , \sha1_round/add_79_3/n250 ,
         \sha1_round/add_79_3/n249 , \sha1_round/add_79_3/n248 ,
         \sha1_round/add_79_3/n247 , \sha1_round/add_79_3/n246 ,
         \sha1_round/add_79_3/n245 , \sha1_round/add_79_3/n244 ,
         \sha1_round/add_79_3/n243 , \sha1_round/add_79_3/n242 ,
         \sha1_round/add_79_3/n241 , \sha1_round/add_79_3/n240 ,
         \sha1_round/add_79_3/n239 , \sha1_round/add_79_3/n238 ,
         \sha1_round/add_79_3/n237 , \sha1_round/add_79_3/n236 ,
         \sha1_round/add_79_3/n235 , \sha1_round/add_79_3/n234 ,
         \sha1_round/add_79_3/n233 , \sha1_round/add_79_3/n232 ,
         \sha1_round/add_79_3/n231 , \sha1_round/add_79_3/n230 ,
         \sha1_round/add_79_3/n229 , \sha1_round/add_79_3/n228 ,
         \sha1_round/add_79_3/n227 , \sha1_round/add_79_3/n226 ,
         \sha1_round/add_79_3/n225 , \sha1_round/add_79_3/n224 ,
         \sha1_round/add_79_3/n223 , \sha1_round/add_79_3/n222 ,
         \sha1_round/add_79_3/n221 , \sha1_round/add_79_3/n220 ,
         \sha1_round/add_79_3/n219 , \sha1_round/add_79_3/n218 ,
         \sha1_round/add_79_3/n217 , \sha1_round/add_79_3/n216 ,
         \sha1_round/add_79_3/n215 , \sha1_round/add_79_3/n214 ,
         \sha1_round/add_79_3/n213 , \sha1_round/add_79_3/n212 ,
         \sha1_round/add_79_3/n211 , \sha1_round/add_79_3/n210 ,
         \sha1_round/add_79_3/n209 , \sha1_round/add_79_3/n208 ,
         \sha1_round/add_79_3/n207 , \sha1_round/add_79_3/n206 ,
         \sha1_round/add_79_3/n205 , \sha1_round/add_79_3/n204 ,
         \sha1_round/add_79_3/n203 , \sha1_round/add_79_3/n202 ,
         \sha1_round/add_79_3/n201 , \sha1_round/add_79_3/n200 ,
         \sha1_round/add_79_3/n199 , \sha1_round/add_79_3/n198 ,
         \sha1_round/add_79_3/n197 , \sha1_round/add_79_3/n196 ,
         \sha1_round/add_79_3/n195 , \sha1_round/add_79_3/n194 ,
         \sha1_round/add_79_3/n193 , \sha1_round/add_79_3/n192 ,
         \sha1_round/add_79_3/n191 , \sha1_round/add_79_3/n190 ,
         \sha1_round/add_79_3/n189 , \sha1_round/add_79_3/n188 ,
         \sha1_round/add_79_3/n187 , \sha1_round/add_79_3/n186 ,
         \sha1_round/add_79_3/n185 , \sha1_round/add_79_3/n184 ,
         \sha1_round/add_79_3/n183 , \sha1_round/add_79_3/n182 ,
         \sha1_round/add_79_3/n181 , \sha1_round/add_79_3/n180 ,
         \sha1_round/add_79_3/n179 , \sha1_round/add_79_3/n178 ,
         \sha1_round/add_79_3/n177 , \sha1_round/add_79_3/n176 ,
         \sha1_round/add_79_3/n175 , \sha1_round/add_79_3/n174 ,
         \sha1_round/add_79_3/n173 , \sha1_round/add_79_3/n172 ,
         \sha1_round/add_79_3/n171 , \sha1_round/add_79_3/n170 ,
         \sha1_round/add_79_3/n169 , \sha1_round/add_79_3/n168 ,
         \sha1_round/add_79_3/n167 , \sha1_round/add_79_3/n166 ,
         \sha1_round/add_79_3/n165 , \sha1_round/add_79_3/n164 ,
         \sha1_round/add_79_3/n163 , \sha1_round/add_79_3/n162 ,
         \sha1_round/add_79_3/n161 , \sha1_round/add_79_3/n160 ,
         \sha1_round/add_79_3/n159 , \sha1_round/add_79_3/n158 ,
         \sha1_round/add_79_3/n157 , \sha1_round/add_79_3/n156 ,
         \sha1_round/add_79_3/n155 , \sha1_round/add_79_3/n154 ,
         \sha1_round/add_79_3/n153 , \sha1_round/add_79_3/n152 ,
         \sha1_round/add_79_3/n151 , \sha1_round/add_79_3/n150 ,
         \sha1_round/add_79_3/n149 , \sha1_round/add_79_3/n148 ,
         \sha1_round/add_79_3/n147 , \sha1_round/add_79_3/n146 ,
         \sha1_round/add_79_3/n145 , \sha1_round/add_79_3/n144 ,
         \sha1_round/add_79_3/n143 , \sha1_round/add_79_3/n142 ,
         \sha1_round/add_79_3/n141 , \sha1_round/add_79_3/n140 ,
         \sha1_round/add_79_3/n139 , \sha1_round/add_79_3/n138 ,
         \sha1_round/add_79_3/n137 , \sha1_round/add_79_3/n136 ,
         \sha1_round/add_79_3/n135 , \sha1_round/add_79_3/n134 ,
         \sha1_round/add_79_3/n133 , \sha1_round/add_79_3/n132 ,
         \sha1_round/add_79_3/n131 , \sha1_round/add_79_3/n130 ,
         \sha1_round/add_79_3/n129 , \sha1_round/add_79_3/n128 ,
         \sha1_round/add_79_3/n127 , \sha1_round/add_79_3/n126 ,
         \sha1_round/add_79_3/n125 , \sha1_round/add_79_3/n124 ,
         \sha1_round/add_79_3/n123 , \sha1_round/add_79_3/n122 ,
         \sha1_round/add_79_3/n121 , \sha1_round/add_79_3/n120 ,
         \sha1_round/add_79_3/n119 , \sha1_round/add_79_3/n118 ,
         \sha1_round/add_79_3/n117 , \sha1_round/add_79_3/n116 ,
         \sha1_round/add_79_3/n115 , \sha1_round/add_79_3/n114 ,
         \sha1_round/add_79_3/n113 , \sha1_round/add_79_3/n112 ,
         \sha1_round/add_79_3/n111 , \sha1_round/add_79_3/n110 ,
         \sha1_round/add_79_3/n109 , \sha1_round/add_79_3/n108 ,
         \sha1_round/add_79_3/n107 , \sha1_round/add_79_3/n106 ,
         \sha1_round/add_79_3/n105 , \sha1_round/add_79_3/n104 ,
         \sha1_round/add_79_3/n103 , \sha1_round/add_79_3/n102 ,
         \sha1_round/add_79_3/n101 , \sha1_round/add_79_3/n100 ,
         \sha1_round/add_79_3/n99 , \sha1_round/add_79_3/n98 ,
         \sha1_round/add_79_3/n97 , \sha1_round/add_79_3/n96 ,
         \sha1_round/add_79_3/n95 , \sha1_round/add_79_3/n94 ,
         \sha1_round/add_79_3/n93 , \sha1_round/add_79_3/n92 ,
         \sha1_round/add_79_3/n91 , \sha1_round/add_79_3/n90 ,
         \sha1_round/add_79_3/n89 , \sha1_round/add_79_3/n88 ,
         \sha1_round/add_79_3/n87 , \sha1_round/add_79_3/n86 ,
         \sha1_round/add_79_3/n85 , \sha1_round/add_79_3/n84 ,
         \sha1_round/add_79_3/n83 , \sha1_round/add_79_3/n82 ,
         \sha1_round/add_79_3/n81 , \sha1_round/add_79_3/n80 ,
         \sha1_round/add_79_3/n79 , \sha1_round/add_79_3/n78 ,
         \sha1_round/add_79_3/n77 , \sha1_round/add_79_3/n76 ,
         \sha1_round/add_79_3/n75 , \sha1_round/add_79_3/n74 ,
         \sha1_round/add_79_3/n73 , \sha1_round/add_79_3/n72 ,
         \sha1_round/add_79_3/n71 , \sha1_round/add_79_3/n70 ,
         \sha1_round/add_79_3/n69 , \sha1_round/add_79_3/n68 ,
         \sha1_round/add_79_3/n67 , \sha1_round/add_79_3/n66 ,
         \sha1_round/add_79_3/n65 , \sha1_round/add_79_3/n64 ,
         \sha1_round/add_79_3/n63 , \sha1_round/add_79_3/n62 ,
         \sha1_round/add_79_3/n61 , \sha1_round/add_79_3/n60 ,
         \sha1_round/add_79_3/n58 , \sha1_round/add_79_3/n57 ,
         \sha1_round/add_79_3/n56 , \sha1_round/add_79_3/n55 ,
         \sha1_round/add_79_3/n54 , \sha1_round/add_79_3/n53 ,
         \sha1_round/add_79_3/n52 , \sha1_round/add_79_3/n51 ,
         \sha1_round/add_79_3/n50 , \sha1_round/add_79_3/n49 ,
         \sha1_round/add_79_3/n48 , \sha1_round/add_79_3/n47 ,
         \sha1_round/add_79_3/n46 , \sha1_round/add_79_3/n45 ,
         \sha1_round/add_79_3/n44 , \sha1_round/add_79_3/n43 ,
         \sha1_round/add_79_3/n42 , \sha1_round/add_79_3/n41 ,
         \sha1_round/add_79_3/n40 , \sha1_round/add_79_3/n39 ,
         \sha1_round/add_79_3/n38 , \sha1_round/add_79_3/n37 ,
         \sha1_round/add_79_3/n36 , \sha1_round/add_79_3/n35 ,
         \sha1_round/add_79_3/n34 , \sha1_round/add_79_3/n33 ,
         \sha1_round/add_79_3/n32 , \sha1_round/add_79_3/n31 ,
         \sha1_round/add_79_3/n30 , \sha1_round/add_79_3/n29 ,
         \sha1_round/add_79_3/n28 , \sha1_round/add_79_3/n27 ,
         \sha1_round/add_79_3/n26 , \sha1_round/add_79_3/n25 ,
         \sha1_round/add_79_3/n24 , \sha1_round/add_79_3/n23 ,
         \sha1_round/add_79_3/n22 , \sha1_round/add_79_3/n21 ,
         \sha1_round/add_79_3/n20 , \sha1_round/add_79_3/n19 ,
         \sha1_round/add_79_3/n18 , \sha1_round/add_79_3/n17 ,
         \sha1_round/add_79_3/n16 , \sha1_round/add_79_3/n15 ,
         \sha1_round/add_79_3/n14 , \sha1_round/add_79_3/n13 ,
         \sha1_round/add_79_3/n12 , \sha1_round/add_79_3/n11 ,
         \sha1_round/add_79_3/n10 , \sha1_round/add_79_3/n9 ,
         \sha1_round/add_79_3/n8 , \sha1_round/add_79_3/n7 ,
         \sha1_round/add_79_3/n6 , \sha1_round/add_79_3/n5 ,
         \sha1_round/add_79_3/n4 , \sha1_round/add_79_3/n3 ,
         \sha1_round/add_79_3/n1 , \sha1_round/add_79/n381 ,
         \sha1_round/add_79/n380 , \sha1_round/add_79/n379 ,
         \sha1_round/add_79/n378 , \sha1_round/add_79/n377 ,
         \sha1_round/add_79/n376 , \sha1_round/add_79/n375 ,
         \sha1_round/add_79/n374 , \sha1_round/add_79/n373 ,
         \sha1_round/add_79/n372 , \sha1_round/add_79/n371 ,
         \sha1_round/add_79/n370 , \sha1_round/add_79/n369 ,
         \sha1_round/add_79/n368 , \sha1_round/add_79/n367 ,
         \sha1_round/add_79/n366 , \sha1_round/add_79/n365 ,
         \sha1_round/add_79/n364 , \sha1_round/add_79/n363 ,
         \sha1_round/add_79/n362 , \sha1_round/add_79/n361 ,
         \sha1_round/add_79/n360 , \sha1_round/add_79/n359 ,
         \sha1_round/add_79/n358 , \sha1_round/add_79/n357 ,
         \sha1_round/add_79/n356 , \sha1_round/add_79/n355 ,
         \sha1_round/add_79/n354 , \sha1_round/add_79/n353 ,
         \sha1_round/add_79/n352 , \sha1_round/add_79/n351 ,
         \sha1_round/add_79/n350 , \sha1_round/add_79/n349 ,
         \sha1_round/add_79/n348 , \sha1_round/add_79/n347 ,
         \sha1_round/add_79/n346 , \sha1_round/add_79/n345 ,
         \sha1_round/add_79/n344 , \sha1_round/add_79/n343 ,
         \sha1_round/add_79/n342 , \sha1_round/add_79/n341 ,
         \sha1_round/add_79/n340 , \sha1_round/add_79/n339 ,
         \sha1_round/add_79/n338 , \sha1_round/add_79/n337 ,
         \sha1_round/add_79/n336 , \sha1_round/add_79/n335 ,
         \sha1_round/add_79/n334 , \sha1_round/add_79/n333 ,
         \sha1_round/add_79/n332 , \sha1_round/add_79/n331 ,
         \sha1_round/add_79/n330 , \sha1_round/add_79/n329 ,
         \sha1_round/add_79/n328 , \sha1_round/add_79/n327 ,
         \sha1_round/add_79/n326 , \sha1_round/add_79/n325 ,
         \sha1_round/add_79/n324 , \sha1_round/add_79/n323 ,
         \sha1_round/add_79/n322 , \sha1_round/add_79/n321 ,
         \sha1_round/add_79/n320 , \sha1_round/add_79/n319 ,
         \sha1_round/add_79/n318 , \sha1_round/add_79/n317 ,
         \sha1_round/add_79/n316 , \sha1_round/add_79/n315 ,
         \sha1_round/add_79/n314 , \sha1_round/add_79/n313 ,
         \sha1_round/add_79/n312 , \sha1_round/add_79/n311 ,
         \sha1_round/add_79/n310 , \sha1_round/add_79/n309 ,
         \sha1_round/add_79/n308 , \sha1_round/add_79/n307 ,
         \sha1_round/add_79/n306 , \sha1_round/add_79/n305 ,
         \sha1_round/add_79/n304 , \sha1_round/add_79/n303 ,
         \sha1_round/add_79/n302 , \sha1_round/add_79/n301 ,
         \sha1_round/add_79/n300 , \sha1_round/add_79/n299 ,
         \sha1_round/add_79/n298 , \sha1_round/add_79/n297 ,
         \sha1_round/add_79/n296 , \sha1_round/add_79/n295 ,
         \sha1_round/add_79/n294 , \sha1_round/add_79/n293 ,
         \sha1_round/add_79/n292 , \sha1_round/add_79/n291 ,
         \sha1_round/add_79/n290 , \sha1_round/add_79/n289 ,
         \sha1_round/add_79/n288 , \sha1_round/add_79/n287 ,
         \sha1_round/add_79/n286 , \sha1_round/add_79/n285 ,
         \sha1_round/add_79/n284 , \sha1_round/add_79/n283 ,
         \sha1_round/add_79/n282 , \sha1_round/add_79/n281 ,
         \sha1_round/add_79/n280 , \sha1_round/add_79/n279 ,
         \sha1_round/add_79/n278 , \sha1_round/add_79/n277 ,
         \sha1_round/add_79/n276 , \sha1_round/add_79/n275 ,
         \sha1_round/add_79/n274 , \sha1_round/add_79/n273 ,
         \sha1_round/add_79/n272 , \sha1_round/add_79/n271 ,
         \sha1_round/add_79/n270 , \sha1_round/add_79/n269 ,
         \sha1_round/add_79/n268 , \sha1_round/add_79/n267 ,
         \sha1_round/add_79/n266 , \sha1_round/add_79/n265 ,
         \sha1_round/add_79/n264 , \sha1_round/add_79/n263 ,
         \sha1_round/add_79/n262 , \sha1_round/add_79/n261 ,
         \sha1_round/add_79/n260 , \sha1_round/add_79/n259 ,
         \sha1_round/add_79/n258 , \sha1_round/add_79/n257 ,
         \sha1_round/add_79/n256 , \sha1_round/add_79/n255 ,
         \sha1_round/add_79/n254 , \sha1_round/add_79/n253 ,
         \sha1_round/add_79/n252 , \sha1_round/add_79/n251 ,
         \sha1_round/add_79/n250 , \sha1_round/add_79/n249 ,
         \sha1_round/add_79/n248 , \sha1_round/add_79/n247 ,
         \sha1_round/add_79/n246 , \sha1_round/add_79/n245 ,
         \sha1_round/add_79/n244 , \sha1_round/add_79/n243 ,
         \sha1_round/add_79/n242 , \sha1_round/add_79/n241 ,
         \sha1_round/add_79/n240 , \sha1_round/add_79/n239 ,
         \sha1_round/add_79/n238 , \sha1_round/add_79/n237 ,
         \sha1_round/add_79/n236 , \sha1_round/add_79/n235 ,
         \sha1_round/add_79/n234 , \sha1_round/add_79/n233 ,
         \sha1_round/add_79/n232 , \sha1_round/add_79/n231 ,
         \sha1_round/add_79/n230 , \sha1_round/add_79/n229 ,
         \sha1_round/add_79/n228 , \sha1_round/add_79/n227 ,
         \sha1_round/add_79/n226 , \sha1_round/add_79/n225 ,
         \sha1_round/add_79/n224 , \sha1_round/add_79/n223 ,
         \sha1_round/add_79/n222 , \sha1_round/add_79/n221 ,
         \sha1_round/add_79/n220 , \sha1_round/add_79/n219 ,
         \sha1_round/add_79/n218 , \sha1_round/add_79/n217 ,
         \sha1_round/add_79/n216 , \sha1_round/add_79/n215 ,
         \sha1_round/add_79/n214 , \sha1_round/add_79/n213 ,
         \sha1_round/add_79/n212 , \sha1_round/add_79/n211 ,
         \sha1_round/add_79/n210 , \sha1_round/add_79/n209 ,
         \sha1_round/add_79/n208 , \sha1_round/add_79/n207 ,
         \sha1_round/add_79/n206 , \sha1_round/add_79/n205 ,
         \sha1_round/add_79/n204 , \sha1_round/add_79/n203 ,
         \sha1_round/add_79/n202 , \sha1_round/add_79/n201 ,
         \sha1_round/add_79/n200 , \sha1_round/add_79/n199 ,
         \sha1_round/add_79/n198 , \sha1_round/add_79/n197 ,
         \sha1_round/add_79/n196 , \sha1_round/add_79/n195 ,
         \sha1_round/add_79/n194 , \sha1_round/add_79/n193 ,
         \sha1_round/add_79/n192 , \sha1_round/add_79/n191 ,
         \sha1_round/add_79/n190 , \sha1_round/add_79/n189 ,
         \sha1_round/add_79/n188 , \sha1_round/add_79/n187 ,
         \sha1_round/add_79/n186 , \sha1_round/add_79/n185 ,
         \sha1_round/add_79/n184 , \sha1_round/add_79/n183 ,
         \sha1_round/add_79/n182 , \sha1_round/add_79/n181 ,
         \sha1_round/add_79/n180 , \sha1_round/add_79/n179 ,
         \sha1_round/add_79/n178 , \sha1_round/add_79/n177 ,
         \sha1_round/add_79/n176 , \sha1_round/add_79/n175 ,
         \sha1_round/add_79/n174 , \sha1_round/add_79/n173 ,
         \sha1_round/add_79/n172 , \sha1_round/add_79/n171 ,
         \sha1_round/add_79/n170 , \sha1_round/add_79/n169 ,
         \sha1_round/add_79/n168 , \sha1_round/add_79/n167 ,
         \sha1_round/add_79/n166 , \sha1_round/add_79/n165 ,
         \sha1_round/add_79/n164 , \sha1_round/add_79/n163 ,
         \sha1_round/add_79/n162 , \sha1_round/add_79/n161 ,
         \sha1_round/add_79/n160 , \sha1_round/add_79/n159 ,
         \sha1_round/add_79/n158 , \sha1_round/add_79/n157 ,
         \sha1_round/add_79/n156 , \sha1_round/add_79/n155 ,
         \sha1_round/add_79/n154 , \sha1_round/add_79/n153 ,
         \sha1_round/add_79/n152 , \sha1_round/add_79/n151 ,
         \sha1_round/add_79/n150 , \sha1_round/add_79/n149 ,
         \sha1_round/add_79/n148 , \sha1_round/add_79/n147 ,
         \sha1_round/add_79/n146 , \sha1_round/add_79/n145 ,
         \sha1_round/add_79/n144 , \sha1_round/add_79/n143 ,
         \sha1_round/add_79/n142 , \sha1_round/add_79/n141 ,
         \sha1_round/add_79/n140 , \sha1_round/add_79/n139 ,
         \sha1_round/add_79/n138 , \sha1_round/add_79/n137 ,
         \sha1_round/add_79/n136 , \sha1_round/add_79/n135 ,
         \sha1_round/add_79/n134 , \sha1_round/add_79/n133 ,
         \sha1_round/add_79/n132 , \sha1_round/add_79/n131 ,
         \sha1_round/add_79/n130 , \sha1_round/add_79/n129 ,
         \sha1_round/add_79/n128 , \sha1_round/add_79/n127 ,
         \sha1_round/add_79/n126 , \sha1_round/add_79/n125 ,
         \sha1_round/add_79/n124 , \sha1_round/add_79/n123 ,
         \sha1_round/add_79/n122 , \sha1_round/add_79/n121 ,
         \sha1_round/add_79/n120 , \sha1_round/add_79/n119 ,
         \sha1_round/add_79/n118 , \sha1_round/add_79/n117 ,
         \sha1_round/add_79/n116 , \sha1_round/add_79/n115 ,
         \sha1_round/add_79/n114 , \sha1_round/add_79/n113 ,
         \sha1_round/add_79/n112 , \sha1_round/add_79/n111 ,
         \sha1_round/add_79/n110 , \sha1_round/add_79/n109 ,
         \sha1_round/add_79/n108 , \sha1_round/add_79/n107 ,
         \sha1_round/add_79/n106 , \sha1_round/add_79/n105 ,
         \sha1_round/add_79/n104 , \sha1_round/add_79/n103 ,
         \sha1_round/add_79/n102 , \sha1_round/add_79/n101 ,
         \sha1_round/add_79/n100 , \sha1_round/add_79/n99 ,
         \sha1_round/add_79/n98 , \sha1_round/add_79/n97 ,
         \sha1_round/add_79/n96 , \sha1_round/add_79/n95 ,
         \sha1_round/add_79/n94 , \sha1_round/add_79/n93 ,
         \sha1_round/add_79/n92 , \sha1_round/add_79/n91 ,
         \sha1_round/add_79/n90 , \sha1_round/add_79/n89 ,
         \sha1_round/add_79/n88 , \sha1_round/add_79/n87 ,
         \sha1_round/add_79/n86 , \sha1_round/add_79/n85 ,
         \sha1_round/add_79/n84 , \sha1_round/add_79/n83 ,
         \sha1_round/add_79/n82 , \sha1_round/add_79/n81 ,
         \sha1_round/add_79/n80 , \sha1_round/add_79/n79 ,
         \sha1_round/add_79/n78 , \sha1_round/add_79/n77 ,
         \sha1_round/add_79/n75 , \sha1_round/add_79/n74 ,
         \sha1_round/add_79/n73 , \sha1_round/add_79/n71 ,
         \sha1_round/add_79/n70 , \sha1_round/add_79/n69 ,
         \sha1_round/add_79/n68 , \sha1_round/add_79/n67 ,
         \sha1_round/add_79/n64 , \sha1_round/add_79/n63 ,
         \sha1_round/add_79/n62 , \sha1_round/add_79/n61 ,
         \sha1_round/add_79/n60 , \sha1_round/add_79/n59 ,
         \sha1_round/add_79/n58 , \sha1_round/add_79/n57 ,
         \sha1_round/add_79/n56 , \sha1_round/add_79/n55 ,
         \sha1_round/add_79/n54 , \sha1_round/add_79/n53 ,
         \sha1_round/add_79/n52 , \sha1_round/add_79/n51 ,
         \sha1_round/add_79/n50 , \sha1_round/add_79/n49 ,
         \sha1_round/add_79/n48 , \sha1_round/add_79/n47 ,
         \sha1_round/add_79/n46 , \sha1_round/add_79/n45 ,
         \sha1_round/add_79/n44 , \sha1_round/add_79/n43 ,
         \sha1_round/add_79/n42 , \sha1_round/add_79/n41 ,
         \sha1_round/add_79/n40 , \sha1_round/add_79/n39 ,
         \sha1_round/add_79/n38 , \sha1_round/add_79/n37 ,
         \sha1_round/add_79/n36 , \sha1_round/add_79/n35 ,
         \sha1_round/add_79/n34 , \sha1_round/add_79/n33 ,
         \sha1_round/add_79/n32 , \sha1_round/add_79/n31 ,
         \sha1_round/add_79/n30 , \sha1_round/add_79/n29 ,
         \sha1_round/add_79/n28 , \sha1_round/add_79/n27 ,
         \sha1_round/add_79/n26 , \sha1_round/add_79/n25 ,
         \sha1_round/add_79/n24 , \sha1_round/add_79/n23 ,
         \sha1_round/add_79/n22 , \sha1_round/add_79/n21 ,
         \sha1_round/add_79/n20 , \sha1_round/add_79/n19 ,
         \sha1_round/add_79/n18 , \sha1_round/add_79/n17 ,
         \sha1_round/add_79/n16 , \sha1_round/add_79/n15 ,
         \sha1_round/add_79/n14 , \sha1_round/add_79/n13 ,
         \sha1_round/add_79/n12 , \sha1_round/add_79/n11 ,
         \sha1_round/add_79/n8 , \sha1_round/add_79/n5 ,
         \sha1_round/add_79/n4 , \sha1_round/add_79/n2 ,
         \sha1_round/add_79/n1 , \sha1_round/add_79_2/n374 ,
         \sha1_round/add_79_2/n373 , \sha1_round/add_79_2/n372 ,
         \sha1_round/add_79_2/n371 , \sha1_round/add_79_2/n370 ,
         \sha1_round/add_79_2/n369 , \sha1_round/add_79_2/n368 ,
         \sha1_round/add_79_2/n367 , \sha1_round/add_79_2/n366 ,
         \sha1_round/add_79_2/n365 , \sha1_round/add_79_2/n364 ,
         \sha1_round/add_79_2/n363 , \sha1_round/add_79_2/n362 ,
         \sha1_round/add_79_2/n361 , \sha1_round/add_79_2/n360 ,
         \sha1_round/add_79_2/n359 , \sha1_round/add_79_2/n358 ,
         \sha1_round/add_79_2/n357 , \sha1_round/add_79_2/n356 ,
         \sha1_round/add_79_2/n355 , \sha1_round/add_79_2/n354 ,
         \sha1_round/add_79_2/n353 , \sha1_round/add_79_2/n352 ,
         \sha1_round/add_79_2/n351 , \sha1_round/add_79_2/n350 ,
         \sha1_round/add_79_2/n349 , \sha1_round/add_79_2/n348 ,
         \sha1_round/add_79_2/n347 , \sha1_round/add_79_2/n346 ,
         \sha1_round/add_79_2/n345 , \sha1_round/add_79_2/n344 ,
         \sha1_round/add_79_2/n343 , \sha1_round/add_79_2/n342 ,
         \sha1_round/add_79_2/n341 , \sha1_round/add_79_2/n340 ,
         \sha1_round/add_79_2/n339 , \sha1_round/add_79_2/n338 ,
         \sha1_round/add_79_2/n337 , \sha1_round/add_79_2/n336 ,
         \sha1_round/add_79_2/n335 , \sha1_round/add_79_2/n334 ,
         \sha1_round/add_79_2/n333 , \sha1_round/add_79_2/n332 ,
         \sha1_round/add_79_2/n331 , \sha1_round/add_79_2/n330 ,
         \sha1_round/add_79_2/n329 , \sha1_round/add_79_2/n328 ,
         \sha1_round/add_79_2/n327 , \sha1_round/add_79_2/n326 ,
         \sha1_round/add_79_2/n325 , \sha1_round/add_79_2/n324 ,
         \sha1_round/add_79_2/n323 , \sha1_round/add_79_2/n322 ,
         \sha1_round/add_79_2/n321 , \sha1_round/add_79_2/n320 ,
         \sha1_round/add_79_2/n319 , \sha1_round/add_79_2/n318 ,
         \sha1_round/add_79_2/n317 , \sha1_round/add_79_2/n316 ,
         \sha1_round/add_79_2/n315 , \sha1_round/add_79_2/n314 ,
         \sha1_round/add_79_2/n313 , \sha1_round/add_79_2/n312 ,
         \sha1_round/add_79_2/n311 , \sha1_round/add_79_2/n310 ,
         \sha1_round/add_79_2/n309 , \sha1_round/add_79_2/n308 ,
         \sha1_round/add_79_2/n307 , \sha1_round/add_79_2/n306 ,
         \sha1_round/add_79_2/n305 , \sha1_round/add_79_2/n304 ,
         \sha1_round/add_79_2/n303 , \sha1_round/add_79_2/n302 ,
         \sha1_round/add_79_2/n301 , \sha1_round/add_79_2/n300 ,
         \sha1_round/add_79_2/n299 , \sha1_round/add_79_2/n298 ,
         \sha1_round/add_79_2/n297 , \sha1_round/add_79_2/n296 ,
         \sha1_round/add_79_2/n295 , \sha1_round/add_79_2/n294 ,
         \sha1_round/add_79_2/n293 , \sha1_round/add_79_2/n292 ,
         \sha1_round/add_79_2/n291 , \sha1_round/add_79_2/n290 ,
         \sha1_round/add_79_2/n289 , \sha1_round/add_79_2/n288 ,
         \sha1_round/add_79_2/n287 , \sha1_round/add_79_2/n286 ,
         \sha1_round/add_79_2/n285 , \sha1_round/add_79_2/n284 ,
         \sha1_round/add_79_2/n283 , \sha1_round/add_79_2/n282 ,
         \sha1_round/add_79_2/n281 , \sha1_round/add_79_2/n280 ,
         \sha1_round/add_79_2/n279 , \sha1_round/add_79_2/n278 ,
         \sha1_round/add_79_2/n277 , \sha1_round/add_79_2/n276 ,
         \sha1_round/add_79_2/n275 , \sha1_round/add_79_2/n274 ,
         \sha1_round/add_79_2/n273 , \sha1_round/add_79_2/n272 ,
         \sha1_round/add_79_2/n271 , \sha1_round/add_79_2/n270 ,
         \sha1_round/add_79_2/n269 , \sha1_round/add_79_2/n268 ,
         \sha1_round/add_79_2/n267 , \sha1_round/add_79_2/n266 ,
         \sha1_round/add_79_2/n265 , \sha1_round/add_79_2/n264 ,
         \sha1_round/add_79_2/n263 , \sha1_round/add_79_2/n262 ,
         \sha1_round/add_79_2/n261 , \sha1_round/add_79_2/n260 ,
         \sha1_round/add_79_2/n259 , \sha1_round/add_79_2/n258 ,
         \sha1_round/add_79_2/n257 , \sha1_round/add_79_2/n256 ,
         \sha1_round/add_79_2/n255 , \sha1_round/add_79_2/n254 ,
         \sha1_round/add_79_2/n253 , \sha1_round/add_79_2/n252 ,
         \sha1_round/add_79_2/n251 , \sha1_round/add_79_2/n250 ,
         \sha1_round/add_79_2/n249 , \sha1_round/add_79_2/n248 ,
         \sha1_round/add_79_2/n247 , \sha1_round/add_79_2/n246 ,
         \sha1_round/add_79_2/n245 , \sha1_round/add_79_2/n244 ,
         \sha1_round/add_79_2/n243 , \sha1_round/add_79_2/n242 ,
         \sha1_round/add_79_2/n241 , \sha1_round/add_79_2/n240 ,
         \sha1_round/add_79_2/n239 , \sha1_round/add_79_2/n238 ,
         \sha1_round/add_79_2/n237 , \sha1_round/add_79_2/n236 ,
         \sha1_round/add_79_2/n235 , \sha1_round/add_79_2/n234 ,
         \sha1_round/add_79_2/n233 , \sha1_round/add_79_2/n232 ,
         \sha1_round/add_79_2/n231 , \sha1_round/add_79_2/n230 ,
         \sha1_round/add_79_2/n229 , \sha1_round/add_79_2/n228 ,
         \sha1_round/add_79_2/n227 , \sha1_round/add_79_2/n226 ,
         \sha1_round/add_79_2/n225 , \sha1_round/add_79_2/n224 ,
         \sha1_round/add_79_2/n223 , \sha1_round/add_79_2/n222 ,
         \sha1_round/add_79_2/n221 , \sha1_round/add_79_2/n220 ,
         \sha1_round/add_79_2/n219 , \sha1_round/add_79_2/n218 ,
         \sha1_round/add_79_2/n217 , \sha1_round/add_79_2/n216 ,
         \sha1_round/add_79_2/n215 , \sha1_round/add_79_2/n214 ,
         \sha1_round/add_79_2/n213 , \sha1_round/add_79_2/n212 ,
         \sha1_round/add_79_2/n211 , \sha1_round/add_79_2/n210 ,
         \sha1_round/add_79_2/n209 , \sha1_round/add_79_2/n208 ,
         \sha1_round/add_79_2/n207 , \sha1_round/add_79_2/n206 ,
         \sha1_round/add_79_2/n205 , \sha1_round/add_79_2/n204 ,
         \sha1_round/add_79_2/n203 , \sha1_round/add_79_2/n202 ,
         \sha1_round/add_79_2/n201 , \sha1_round/add_79_2/n200 ,
         \sha1_round/add_79_2/n199 , \sha1_round/add_79_2/n198 ,
         \sha1_round/add_79_2/n197 , \sha1_round/add_79_2/n196 ,
         \sha1_round/add_79_2/n195 , \sha1_round/add_79_2/n194 ,
         \sha1_round/add_79_2/n193 , \sha1_round/add_79_2/n192 ,
         \sha1_round/add_79_2/n191 , \sha1_round/add_79_2/n190 ,
         \sha1_round/add_79_2/n189 , \sha1_round/add_79_2/n188 ,
         \sha1_round/add_79_2/n187 , \sha1_round/add_79_2/n186 ,
         \sha1_round/add_79_2/n185 , \sha1_round/add_79_2/n184 ,
         \sha1_round/add_79_2/n183 , \sha1_round/add_79_2/n182 ,
         \sha1_round/add_79_2/n181 , \sha1_round/add_79_2/n180 ,
         \sha1_round/add_79_2/n179 , \sha1_round/add_79_2/n178 ,
         \sha1_round/add_79_2/n177 , \sha1_round/add_79_2/n176 ,
         \sha1_round/add_79_2/n175 , \sha1_round/add_79_2/n174 ,
         \sha1_round/add_79_2/n173 , \sha1_round/add_79_2/n172 ,
         \sha1_round/add_79_2/n171 , \sha1_round/add_79_2/n170 ,
         \sha1_round/add_79_2/n169 , \sha1_round/add_79_2/n168 ,
         \sha1_round/add_79_2/n167 , \sha1_round/add_79_2/n166 ,
         \sha1_round/add_79_2/n165 , \sha1_round/add_79_2/n164 ,
         \sha1_round/add_79_2/n163 , \sha1_round/add_79_2/n162 ,
         \sha1_round/add_79_2/n161 , \sha1_round/add_79_2/n160 ,
         \sha1_round/add_79_2/n159 , \sha1_round/add_79_2/n158 ,
         \sha1_round/add_79_2/n157 , \sha1_round/add_79_2/n156 ,
         \sha1_round/add_79_2/n155 , \sha1_round/add_79_2/n154 ,
         \sha1_round/add_79_2/n153 , \sha1_round/add_79_2/n152 ,
         \sha1_round/add_79_2/n151 , \sha1_round/add_79_2/n150 ,
         \sha1_round/add_79_2/n149 , \sha1_round/add_79_2/n148 ,
         \sha1_round/add_79_2/n147 , \sha1_round/add_79_2/n146 ,
         \sha1_round/add_79_2/n145 , \sha1_round/add_79_2/n144 ,
         \sha1_round/add_79_2/n143 , \sha1_round/add_79_2/n142 ,
         \sha1_round/add_79_2/n141 , \sha1_round/add_79_2/n140 ,
         \sha1_round/add_79_2/n139 , \sha1_round/add_79_2/n138 ,
         \sha1_round/add_79_2/n137 , \sha1_round/add_79_2/n136 ,
         \sha1_round/add_79_2/n135 , \sha1_round/add_79_2/n134 ,
         \sha1_round/add_79_2/n133 , \sha1_round/add_79_2/n132 ,
         \sha1_round/add_79_2/n131 , \sha1_round/add_79_2/n130 ,
         \sha1_round/add_79_2/n129 , \sha1_round/add_79_2/n128 ,
         \sha1_round/add_79_2/n127 , \sha1_round/add_79_2/n126 ,
         \sha1_round/add_79_2/n125 , \sha1_round/add_79_2/n124 ,
         \sha1_round/add_79_2/n123 , \sha1_round/add_79_2/n122 ,
         \sha1_round/add_79_2/n121 , \sha1_round/add_79_2/n120 ,
         \sha1_round/add_79_2/n119 , \sha1_round/add_79_2/n118 ,
         \sha1_round/add_79_2/n117 , \sha1_round/add_79_2/n116 ,
         \sha1_round/add_79_2/n115 , \sha1_round/add_79_2/n114 ,
         \sha1_round/add_79_2/n113 , \sha1_round/add_79_2/n112 ,
         \sha1_round/add_79_2/n111 , \sha1_round/add_79_2/n110 ,
         \sha1_round/add_79_2/n109 , \sha1_round/add_79_2/n108 ,
         \sha1_round/add_79_2/n107 , \sha1_round/add_79_2/n106 ,
         \sha1_round/add_79_2/n105 , \sha1_round/add_79_2/n104 ,
         \sha1_round/add_79_2/n103 , \sha1_round/add_79_2/n102 ,
         \sha1_round/add_79_2/n101 , \sha1_round/add_79_2/n100 ,
         \sha1_round/add_79_2/n99 , \sha1_round/add_79_2/n98 ,
         \sha1_round/add_79_2/n97 , \sha1_round/add_79_2/n96 ,
         \sha1_round/add_79_2/n95 , \sha1_round/add_79_2/n94 ,
         \sha1_round/add_79_2/n93 , \sha1_round/add_79_2/n92 ,
         \sha1_round/add_79_2/n91 , \sha1_round/add_79_2/n90 ,
         \sha1_round/add_79_2/n89 , \sha1_round/add_79_2/n88 ,
         \sha1_round/add_79_2/n87 , \sha1_round/add_79_2/n86 ,
         \sha1_round/add_79_2/n85 , \sha1_round/add_79_2/n84 ,
         \sha1_round/add_79_2/n83 , \sha1_round/add_79_2/n82 ,
         \sha1_round/add_79_2/n81 , \sha1_round/add_79_2/n80 ,
         \sha1_round/add_79_2/n79 , \sha1_round/add_79_2/n78 ,
         \sha1_round/add_79_2/n77 , \sha1_round/add_79_2/n76 ,
         \sha1_round/add_79_2/n75 , \sha1_round/add_79_2/n74 ,
         \sha1_round/add_79_2/n73 , \sha1_round/add_79_2/n72 ,
         \sha1_round/add_79_2/n71 , \sha1_round/add_79_2/n70 ,
         \sha1_round/add_79_2/n69 , \sha1_round/add_79_2/n68 ,
         \sha1_round/add_79_2/n67 , \sha1_round/add_79_2/n66 ,
         \sha1_round/add_79_2/n65 , \sha1_round/add_79_2/n64 ,
         \sha1_round/add_79_2/n63 , \sha1_round/add_79_2/n62 ,
         \sha1_round/add_79_2/n61 , \sha1_round/add_79_2/n60 ,
         \sha1_round/add_79_2/n59 , \sha1_round/add_79_2/n58 ,
         \sha1_round/add_79_2/n57 , \sha1_round/add_79_2/n56 ,
         \sha1_round/add_79_2/n55 , \sha1_round/add_79_2/n54 ,
         \sha1_round/add_79_2/n53 , \sha1_round/add_79_2/n52 ,
         \sha1_round/add_79_2/n51 , \sha1_round/add_79_2/n50 ,
         \sha1_round/add_79_2/n49 , \sha1_round/add_79_2/n48 ,
         \sha1_round/add_79_2/n47 , \sha1_round/add_79_2/n46 ,
         \sha1_round/add_79_2/n45 , \sha1_round/add_79_2/n44 ,
         \sha1_round/add_79_2/n43 , \sha1_round/add_79_2/n42 ,
         \sha1_round/add_79_2/n41 , \sha1_round/add_79_2/n40 ,
         \sha1_round/add_79_2/n39 , \sha1_round/add_79_2/n38 ,
         \sha1_round/add_79_2/n37 , \sha1_round/add_79_2/n36 ,
         \sha1_round/add_79_2/n35 , \sha1_round/add_79_2/n34 ,
         \sha1_round/add_79_2/n33 , \sha1_round/add_79_2/n32 ,
         \sha1_round/add_79_2/n31 , \sha1_round/add_79_2/n29 ,
         \sha1_round/add_79_2/n28 , \sha1_round/add_79_2/n27 ,
         \sha1_round/add_79_2/n25 , \sha1_round/add_79_2/n24 ,
         \sha1_round/add_79_2/n23 , \sha1_round/add_79_2/n22 ,
         \sha1_round/add_79_2/n21 , \sha1_round/add_79_2/n20 ,
         \sha1_round/add_79_2/n19 , \sha1_round/add_79_2/n18 ,
         \sha1_round/add_79_2/n17 , \sha1_round/add_79_2/n16 ,
         \sha1_round/add_79_2/n15 , \sha1_round/add_79_2/n14 ,
         \sha1_round/add_79_2/n13 , \sha1_round/add_79_2/n12 ,
         \sha1_round/add_79_2/n11 , \sha1_round/add_79_2/n10 ,
         \sha1_round/add_79_2/n9 , \sha1_round/add_79_2/n8 ,
         \sha1_round/add_79_2/n7 , \sha1_round/add_79_2/n6 ,
         \sha1_round/add_79_2/n5 , \sha1_round/add_79_2/n4 ,
         \sha1_round/add_79_2/n3 , \sha1_round/add_79_2/n2 ,
         \sha1_round/add_79_2/n1 , \rnd_cnt_reg/n12 , \rnd_cnt_reg/n10 ,
         \rnd_cnt_reg/n70 , \rnd_cnt_reg/n60 , \rnd_cnt_reg/n40 ,
         \rnd_cnt_reg/n2 , \rnd_cnt_reg/N9 , \rnd_cnt_reg/N8 ,
         \rnd_cnt_reg/N7 , \rnd_cnt_reg/N6 , \rnd_cnt_reg/N5 ,
         \rnd_cnt_reg/N4 , \rnd_cnt_reg/N3 , \state_reg/n2 , \state_reg/N4 ,
         \state_reg/N3 , \w_reg/n1070 , \w_reg/n1060 , \w_reg/n1050 ,
         \w_reg/n1040 , \w_reg/n1030 , \w_reg/n1020 , \w_reg/n1010 ,
         \w_reg/n1000 , \w_reg/n990 , \w_reg/n980 , \w_reg/n970 , \w_reg/n960 ,
         \w_reg/n950 , \w_reg/n940 , \w_reg/n930 , \w_reg/n920 , \w_reg/n910 ,
         \w_reg/n900 , \w_reg/n890 , \w_reg/n880 , \w_reg/n870 , \w_reg/n860 ,
         \w_reg/n850 , \w_reg/n840 , \w_reg/n830 , \w_reg/n820 , \w_reg/n810 ,
         \w_reg/n800 , \w_reg/n790 , \w_reg/n780 , \w_reg/n770 , \w_reg/n760 ,
         \w_reg/n750 , \w_reg/n740 , \w_reg/n730 , \w_reg/n720 , \w_reg/n710 ,
         \w_reg/n700 , \w_reg/n690 , \w_reg/n680 , \w_reg/n670 , \w_reg/n660 ,
         \w_reg/n650 , \w_reg/n640 , \w_reg/n630 , \w_reg/n620 , \w_reg/n610 ,
         \w_reg/n600 , \w_reg/N514 , \w_reg/N513 , \w_reg/N512 , \w_reg/N511 ,
         \w_reg/N510 , \w_reg/N509 , \w_reg/N508 , \w_reg/N507 , \w_reg/N506 ,
         \w_reg/N505 , \w_reg/N504 , \w_reg/N503 , \w_reg/N502 , \w_reg/N501 ,
         \w_reg/N500 , \w_reg/N499 , \w_reg/N498 , \w_reg/N497 , \w_reg/N496 ,
         \w_reg/N495 , \w_reg/N494 , \w_reg/N493 , \w_reg/N492 , \w_reg/N491 ,
         \w_reg/N490 , \w_reg/N489 , \w_reg/N488 , \w_reg/N487 , \w_reg/N486 ,
         \w_reg/N485 , \w_reg/N484 , \w_reg/N483 , \w_reg/N482 , \w_reg/N481 ,
         \w_reg/N480 , \w_reg/N479 , \w_reg/N478 , \w_reg/N477 , \w_reg/N476 ,
         \w_reg/N475 , \w_reg/N474 , \w_reg/N473 , \w_reg/N472 , \w_reg/N471 ,
         \w_reg/N470 , \w_reg/N469 , \w_reg/N468 , \w_reg/N467 , \w_reg/N466 ,
         \w_reg/N465 , \w_reg/N464 , \w_reg/N463 , \w_reg/N462 , \w_reg/N461 ,
         \w_reg/N460 , \w_reg/N459 , \w_reg/N458 , \w_reg/N457 , \w_reg/N456 ,
         \w_reg/N455 , \w_reg/N454 , \w_reg/N453 , \w_reg/N452 , \w_reg/N451 ,
         \w_reg/N450 , \w_reg/N449 , \w_reg/N448 , \w_reg/N447 , \w_reg/N446 ,
         \w_reg/N445 , \w_reg/N444 , \w_reg/N443 , \w_reg/N442 , \w_reg/N441 ,
         \w_reg/N440 , \w_reg/N439 , \w_reg/N438 , \w_reg/N437 , \w_reg/N436 ,
         \w_reg/N435 , \w_reg/N434 , \w_reg/N433 , \w_reg/N432 , \w_reg/N431 ,
         \w_reg/N430 , \w_reg/N429 , \w_reg/N428 , \w_reg/N427 , \w_reg/N426 ,
         \w_reg/N425 , \w_reg/N424 , \w_reg/N423 , \w_reg/N422 , \w_reg/N421 ,
         \w_reg/N420 , \w_reg/N419 , \w_reg/N418 , \w_reg/N417 , \w_reg/N416 ,
         \w_reg/N415 , \w_reg/N414 , \w_reg/N413 , \w_reg/N412 , \w_reg/N411 ,
         \w_reg/N410 , \w_reg/N409 , \w_reg/N408 , \w_reg/N407 , \w_reg/N406 ,
         \w_reg/N405 , \w_reg/N404 , \w_reg/N403 , \w_reg/N402 , \w_reg/N401 ,
         \w_reg/N400 , \w_reg/N399 , \w_reg/N398 , \w_reg/N397 , \w_reg/N396 ,
         \w_reg/N395 , \w_reg/N394 , \w_reg/N393 , \w_reg/N392 , \w_reg/N391 ,
         \w_reg/N390 , \w_reg/N389 , \w_reg/N388 , \w_reg/N387 , \w_reg/N386 ,
         \w_reg/N385 , \w_reg/N384 , \w_reg/N383 , \w_reg/N382 , \w_reg/N381 ,
         \w_reg/N380 , \w_reg/N379 , \w_reg/N378 , \w_reg/N377 , \w_reg/N376 ,
         \w_reg/N375 , \w_reg/N374 , \w_reg/N373 , \w_reg/N372 , \w_reg/N371 ,
         \w_reg/N370 , \w_reg/N369 , \w_reg/N368 , \w_reg/N367 , \w_reg/N366 ,
         \w_reg/N365 , \w_reg/N364 , \w_reg/N363 , \w_reg/N362 , \w_reg/N361 ,
         \w_reg/N360 , \w_reg/N359 , \w_reg/N358 , \w_reg/N357 , \w_reg/N356 ,
         \w_reg/N355 , \w_reg/N354 , \w_reg/N353 , \w_reg/N352 , \w_reg/N351 ,
         \w_reg/N350 , \w_reg/N349 , \w_reg/N348 , \w_reg/N347 , \w_reg/N346 ,
         \w_reg/N345 , \w_reg/N344 , \w_reg/N343 , \w_reg/N342 , \w_reg/N341 ,
         \w_reg/N340 , \w_reg/N339 , \w_reg/N338 , \w_reg/N337 , \w_reg/N336 ,
         \w_reg/N335 , \w_reg/N334 , \w_reg/N333 , \w_reg/N332 , \w_reg/N331 ,
         \w_reg/N330 , \w_reg/N329 , \w_reg/N328 , \w_reg/N327 , \w_reg/N326 ,
         \w_reg/N325 , \w_reg/N324 , \w_reg/N323 , \w_reg/N322 , \w_reg/N321 ,
         \w_reg/N320 , \w_reg/N319 , \w_reg/N318 , \w_reg/N317 , \w_reg/N316 ,
         \w_reg/N315 , \w_reg/N314 , \w_reg/N313 , \w_reg/N312 , \w_reg/N311 ,
         \w_reg/N310 , \w_reg/N309 , \w_reg/N308 , \w_reg/N307 , \w_reg/N306 ,
         \w_reg/N305 , \w_reg/N304 , \w_reg/N303 , \w_reg/N302 , \w_reg/N301 ,
         \w_reg/N300 , \w_reg/N299 , \w_reg/N298 , \w_reg/N297 , \w_reg/N296 ,
         \w_reg/N295 , \w_reg/N294 , \w_reg/N293 , \w_reg/N292 , \w_reg/N291 ,
         \w_reg/N290 , \w_reg/N289 , \w_reg/N288 , \w_reg/N287 , \w_reg/N286 ,
         \w_reg/N285 , \w_reg/N284 , \w_reg/N283 , \w_reg/N282 , \w_reg/N281 ,
         \w_reg/N280 , \w_reg/N279 , \w_reg/N278 , \w_reg/N277 , \w_reg/N276 ,
         \w_reg/N275 , \w_reg/N274 , \w_reg/N273 , \w_reg/N272 , \w_reg/N271 ,
         \w_reg/N270 , \w_reg/N269 , \w_reg/N268 , \w_reg/N267 , \w_reg/N266 ,
         \w_reg/N265 , \w_reg/N264 , \w_reg/N263 , \w_reg/N262 , \w_reg/N261 ,
         \w_reg/N260 , \w_reg/N259 , \w_reg/N258 , \w_reg/N257 , \w_reg/N256 ,
         \w_reg/N255 , \w_reg/N254 , \w_reg/N253 , \w_reg/N252 , \w_reg/N251 ,
         \w_reg/N250 , \w_reg/N249 , \w_reg/N248 , \w_reg/N247 , \w_reg/N246 ,
         \w_reg/N245 , \w_reg/N244 , \w_reg/N243 , \w_reg/N242 , \w_reg/N241 ,
         \w_reg/N240 , \w_reg/N239 , \w_reg/N238 , \w_reg/N237 , \w_reg/N236 ,
         \w_reg/N235 , \w_reg/N234 , \w_reg/N233 , \w_reg/N232 , \w_reg/N231 ,
         \w_reg/N230 , \w_reg/N229 , \w_reg/N228 , \w_reg/N227 , \w_reg/N226 ,
         \w_reg/N225 , \w_reg/N224 , \w_reg/N223 , \w_reg/N222 , \w_reg/N221 ,
         \w_reg/N220 , \w_reg/N219 , \w_reg/N218 , \w_reg/N217 , \w_reg/N216 ,
         \w_reg/N215 , \w_reg/N214 , \w_reg/N213 , \w_reg/N212 , \w_reg/N211 ,
         \w_reg/N210 , \w_reg/N209 , \w_reg/N208 , \w_reg/N207 , \w_reg/N206 ,
         \w_reg/N205 , \w_reg/N204 , \w_reg/N203 , \w_reg/N202 , \w_reg/N201 ,
         \w_reg/N200 , \w_reg/N199 , \w_reg/N198 , \w_reg/N197 , \w_reg/N196 ,
         \w_reg/N195 , \w_reg/N194 , \w_reg/N193 , \w_reg/N192 , \w_reg/N191 ,
         \w_reg/N190 , \w_reg/N189 , \w_reg/N188 , \w_reg/N187 , \w_reg/N186 ,
         \w_reg/N185 , \w_reg/N184 , \w_reg/N183 , \w_reg/N182 , \w_reg/N181 ,
         \w_reg/N180 , \w_reg/N179 , \w_reg/N178 , \w_reg/N177 , \w_reg/N176 ,
         \w_reg/N175 , \w_reg/N174 , \w_reg/N173 , \w_reg/N172 , \w_reg/N171 ,
         \w_reg/N170 , \w_reg/N169 , \w_reg/N168 , \w_reg/N167 , \w_reg/N166 ,
         \w_reg/N165 , \w_reg/N164 , \w_reg/N163 , \w_reg/N162 , \w_reg/N161 ,
         \w_reg/N160 , \w_reg/N159 , \w_reg/N158 , \w_reg/N157 , \w_reg/N156 ,
         \w_reg/N155 , \w_reg/N154 , \w_reg/N153 , \w_reg/N152 , \w_reg/N151 ,
         \w_reg/N150 , \w_reg/N149 , \w_reg/N148 , \w_reg/N147 , \w_reg/N146 ,
         \w_reg/N145 , \w_reg/N144 , \w_reg/N143 , \w_reg/N142 , \w_reg/N141 ,
         \w_reg/N140 , \w_reg/N139 , \w_reg/N138 , \w_reg/N137 , \w_reg/N136 ,
         \w_reg/N135 , \w_reg/N134 , \w_reg/N133 , \w_reg/N132 , \w_reg/N131 ,
         \w_reg/N130 , \w_reg/N129 , \w_reg/N128 , \w_reg/N127 , \w_reg/N126 ,
         \w_reg/N125 , \w_reg/N124 , \w_reg/N123 , \w_reg/N122 , \w_reg/N121 ,
         \w_reg/N120 , \w_reg/N119 , \w_reg/N118 , \w_reg/N117 , \w_reg/N116 ,
         \w_reg/N115 , \w_reg/N114 , \w_reg/N113 , \w_reg/N112 , \w_reg/N111 ,
         \w_reg/N110 , \w_reg/N109 , \w_reg/N108 , \w_reg/N107 , \w_reg/N106 ,
         \w_reg/N105 , \w_reg/N104 , \w_reg/N103 , \w_reg/N102 , \w_reg/N101 ,
         \w_reg/N100 , \w_reg/N99 , \w_reg/N98 , \w_reg/N97 , \w_reg/N96 ,
         \w_reg/N95 , \w_reg/N94 , \w_reg/N93 , \w_reg/N92 , \w_reg/N91 ,
         \w_reg/N90 , \w_reg/N89 , \w_reg/N88 , \w_reg/N87 , \w_reg/N86 ,
         \w_reg/N85 , \w_reg/N84 , \w_reg/N83 , \w_reg/N82 , \w_reg/N81 ,
         \w_reg/N80 , \w_reg/N79 , \w_reg/N78 , \w_reg/N77 , \w_reg/N76 ,
         \w_reg/N75 , \w_reg/N74 , \w_reg/N73 , \w_reg/N72 , \w_reg/N71 ,
         \w_reg/N70 , \w_reg/N69 , \w_reg/N68 , \w_reg/N67 , \w_reg/N66 ,
         \w_reg/N65 , \w_reg/N64 , \w_reg/N63 , \w_reg/N62 , \w_reg/N61 ,
         \w_reg/N60 , \w_reg/N59 , \w_reg/N58 , \w_reg/N57 , \w_reg/N56 ,
         \w_reg/N55 , \w_reg/N54 , \w_reg/N53 , \w_reg/N52 , \w_reg/N51 ,
         \w_reg/N50 , \w_reg/N49 , \w_reg/N48 , \w_reg/N47 , \w_reg/N46 ,
         \w_reg/N45 , \w_reg/N44 , \w_reg/N43 , \w_reg/N42 , \w_reg/N41 ,
         \w_reg/N40 , \w_reg/N39 , \w_reg/N38 , \w_reg/N37 , \w_reg/N36 ,
         \w_reg/N35 , \w_reg/N34 , \w_reg/N33 , \w_reg/N32 , \w_reg/N31 ,
         \w_reg/N30 , \w_reg/N29 , \w_reg/N28 , \w_reg/N27 , \w_reg/N26 ,
         \w_reg/N25 , \w_reg/N24 , \w_reg/N23 , \w_reg/N22 , \w_reg/N21 ,
         \w_reg/N20 , \w_reg/N19 , \w_reg/N18 , \w_reg/N17 , \w_reg/N16 ,
         \w_reg/N15 , \w_reg/N14 , \w_reg/N13 , \w_reg/N12 , \w_reg/N11 ,
         \w_reg/N10 , \w_reg/N9 , \w_reg/N8 , \w_reg/N7 , \w_reg/N6 ,
         \w_reg/N5 , \w_reg/N4 , \w_reg/N3 , \cv_reg/n330 , \cv_reg/n320 ,
         \cv_reg/n310 , \cv_reg/n300 , \cv_reg/n290 , \cv_reg/n280 ,
         \cv_reg/n270 , \cv_reg/n260 , \cv_reg/n250 , \cv_reg/n240 ,
         \cv_reg/n230 , \cv_reg/n220 , \cv_reg/n210 , \cv_reg/n200 ,
         \cv_reg/n190 , \cv_reg/n180 , \cv_reg/n170 , \cv_reg/N162 ,
         \cv_reg/N161 , \cv_reg/N160 , \cv_reg/N159 , \cv_reg/N158 ,
         \cv_reg/N157 , \cv_reg/N156 , \cv_reg/N155 , \cv_reg/N154 ,
         \cv_reg/N153 , \cv_reg/N152 , \cv_reg/N151 , \cv_reg/N150 ,
         \cv_reg/N149 , \cv_reg/N148 , \cv_reg/N147 , \cv_reg/N146 ,
         \cv_reg/N145 , \cv_reg/N144 , \cv_reg/N143 , \cv_reg/N142 ,
         \cv_reg/N141 , \cv_reg/N140 , \cv_reg/N139 , \cv_reg/N138 ,
         \cv_reg/N137 , \cv_reg/N136 , \cv_reg/N135 , \cv_reg/N134 ,
         \cv_reg/N133 , \cv_reg/N132 , \cv_reg/N131 , \cv_reg/N130 ,
         \cv_reg/N129 , \cv_reg/N128 , \cv_reg/N127 , \cv_reg/N126 ,
         \cv_reg/N125 , \cv_reg/N124 , \cv_reg/N123 , \cv_reg/N122 ,
         \cv_reg/N121 , \cv_reg/N120 , \cv_reg/N119 , \cv_reg/N118 ,
         \cv_reg/N117 , \cv_reg/N116 , \cv_reg/N115 , \cv_reg/N114 ,
         \cv_reg/N113 , \cv_reg/N112 , \cv_reg/N111 , \cv_reg/N110 ,
         \cv_reg/N109 , \cv_reg/N108 , \cv_reg/N107 , \cv_reg/N106 ,
         \cv_reg/N105 , \cv_reg/N104 , \cv_reg/N103 , \cv_reg/N102 ,
         \cv_reg/N101 , \cv_reg/N100 , \cv_reg/N99 , \cv_reg/N98 ,
         \cv_reg/N97 , \cv_reg/N96 , \cv_reg/N95 , \cv_reg/N94 , \cv_reg/N93 ,
         \cv_reg/N92 , \cv_reg/N91 , \cv_reg/N90 , \cv_reg/N89 , \cv_reg/N88 ,
         \cv_reg/N87 , \cv_reg/N86 , \cv_reg/N85 , \cv_reg/N84 , \cv_reg/N83 ,
         \cv_reg/N82 , \cv_reg/N81 , \cv_reg/N80 , \cv_reg/N79 , \cv_reg/N78 ,
         \cv_reg/N77 , \cv_reg/N76 , \cv_reg/N75 , \cv_reg/N74 , \cv_reg/N73 ,
         \cv_reg/N72 , \cv_reg/N71 , \cv_reg/N70 , \cv_reg/N69 , \cv_reg/N68 ,
         \cv_reg/N67 , \cv_reg/N66 , \cv_reg/N65 , \cv_reg/N64 , \cv_reg/N63 ,
         \cv_reg/N62 , \cv_reg/N61 , \cv_reg/N60 , \cv_reg/N59 , \cv_reg/N58 ,
         \cv_reg/N57 , \cv_reg/N56 , \cv_reg/N55 , \cv_reg/N54 , \cv_reg/N53 ,
         \cv_reg/N52 , \cv_reg/N51 , \cv_reg/N50 , \cv_reg/N49 , \cv_reg/N48 ,
         \cv_reg/N47 , \cv_reg/N46 , \cv_reg/N45 , \cv_reg/N44 , \cv_reg/N43 ,
         \cv_reg/N42 , \cv_reg/N41 , \cv_reg/N40 , \cv_reg/N39 , \cv_reg/N38 ,
         \cv_reg/N37 , \cv_reg/N36 , \cv_reg/N35 , \cv_reg/N34 , \cv_reg/N33 ,
         \cv_reg/N32 , \cv_reg/N31 , \cv_reg/N30 , \cv_reg/N29 , \cv_reg/N28 ,
         \cv_reg/N27 , \cv_reg/N26 , \cv_reg/N25 , \cv_reg/N24 , \cv_reg/N23 ,
         \cv_reg/N22 , \cv_reg/N21 , \cv_reg/N20 , \cv_reg/N19 , \cv_reg/N18 ,
         \cv_reg/N17 , \cv_reg/N16 , \cv_reg/N15 , \cv_reg/N14 , \cv_reg/N13 ,
         \cv_reg/N12 , \cv_reg/N11 , \cv_reg/N10 , \cv_reg/N9 , \cv_reg/N8 ,
         \cv_reg/N7 , \cv_reg/N6 , \cv_reg/N5 , \cv_reg/N4 , \cv_reg/N3 ,
         \rnd_reg/n320 , \rnd_reg/n310 , \rnd_reg/n300 , \rnd_reg/n290 ,
         \rnd_reg/n280 , \rnd_reg/n270 , \rnd_reg/n260 , \rnd_reg/n250 ,
         \rnd_reg/n240 , \rnd_reg/n230 , \rnd_reg/n220 , \rnd_reg/n210 ,
         \rnd_reg/n200 , \rnd_reg/n190 , \rnd_reg/n180 , \rnd_reg/n170 ,
         \rnd_reg/N162 , \rnd_reg/N161 , \rnd_reg/N160 , \rnd_reg/N159 ,
         \rnd_reg/N158 , \rnd_reg/N157 , \rnd_reg/N156 , \rnd_reg/N155 ,
         \rnd_reg/N154 , \rnd_reg/N153 , \rnd_reg/N152 , \rnd_reg/N151 ,
         \rnd_reg/N150 , \rnd_reg/N149 , \rnd_reg/N148 , \rnd_reg/N147 ,
         \rnd_reg/N146 , \rnd_reg/N145 , \rnd_reg/N144 , \rnd_reg/N143 ,
         \rnd_reg/N142 , \rnd_reg/N141 , \rnd_reg/N140 , \rnd_reg/N139 ,
         \rnd_reg/N138 , \rnd_reg/N137 , \rnd_reg/N136 , \rnd_reg/N135 ,
         \rnd_reg/N134 , \rnd_reg/N133 , \rnd_reg/N132 , \rnd_reg/N131 ,
         \rnd_reg/N130 , \rnd_reg/N129 , \rnd_reg/N128 , \rnd_reg/N127 ,
         \rnd_reg/N126 , \rnd_reg/N125 , \rnd_reg/N124 , \rnd_reg/N123 ,
         \rnd_reg/N122 , \rnd_reg/N121 , \rnd_reg/N120 , \rnd_reg/N119 ,
         \rnd_reg/N118 , \rnd_reg/N117 , \rnd_reg/N116 , \rnd_reg/N115 ,
         \rnd_reg/N114 , \rnd_reg/N113 , \rnd_reg/N112 , \rnd_reg/N111 ,
         \rnd_reg/N110 , \rnd_reg/N109 , \rnd_reg/N108 , \rnd_reg/N107 ,
         \rnd_reg/N106 , \rnd_reg/N105 , \rnd_reg/N104 , \rnd_reg/N103 ,
         \rnd_reg/N102 , \rnd_reg/N101 , \rnd_reg/N100 , \rnd_reg/N99 ,
         \rnd_reg/N98 , \rnd_reg/N97 , \rnd_reg/N96 , \rnd_reg/N95 ,
         \rnd_reg/N94 , \rnd_reg/N93 , \rnd_reg/N92 , \rnd_reg/N91 ,
         \rnd_reg/N90 , \rnd_reg/N89 , \rnd_reg/N88 , \rnd_reg/N87 ,
         \rnd_reg/N86 , \rnd_reg/N85 , \rnd_reg/N84 , \rnd_reg/N83 ,
         \rnd_reg/N82 , \rnd_reg/N81 , \rnd_reg/N80 , \rnd_reg/N79 ,
         \rnd_reg/N78 , \rnd_reg/N77 , \rnd_reg/N76 , \rnd_reg/N75 ,
         \rnd_reg/N74 , \rnd_reg/N73 , \rnd_reg/N72 , \rnd_reg/N71 ,
         \rnd_reg/N70 , \rnd_reg/N69 , \rnd_reg/N68 , \rnd_reg/N67 ,
         \rnd_reg/N66 , \rnd_reg/N65 , \rnd_reg/N64 , \rnd_reg/N63 ,
         \rnd_reg/N62 , \rnd_reg/N61 , \rnd_reg/N60 , \rnd_reg/N59 ,
         \rnd_reg/N58 , \rnd_reg/N57 , \rnd_reg/N56 , \rnd_reg/N55 ,
         \rnd_reg/N54 , \rnd_reg/N53 , \rnd_reg/N52 , \rnd_reg/N51 ,
         \rnd_reg/N50 , \rnd_reg/N49 , \rnd_reg/N48 , \rnd_reg/N47 ,
         \rnd_reg/N46 , \rnd_reg/N45 , \rnd_reg/N44 , \rnd_reg/N43 ,
         \rnd_reg/N42 , \rnd_reg/N41 , \rnd_reg/N40 , \rnd_reg/N39 ,
         \rnd_reg/N38 , \rnd_reg/N37 , \rnd_reg/N36 , \rnd_reg/N35 ,
         \rnd_reg/N34 , \rnd_reg/N33 , \rnd_reg/N32 , \rnd_reg/N31 ,
         \rnd_reg/N30 , \rnd_reg/N29 , \rnd_reg/N28 , \rnd_reg/N27 ,
         \rnd_reg/N26 , \rnd_reg/N25 , \rnd_reg/N24 , \rnd_reg/N23 ,
         \rnd_reg/N22 , \rnd_reg/N21 , \rnd_reg/N20 , \rnd_reg/N19 ,
         \rnd_reg/N18 , \rnd_reg/N17 , \rnd_reg/N16 , \rnd_reg/N15 ,
         \rnd_reg/N14 , \rnd_reg/N13 , \rnd_reg/N12 , \rnd_reg/N11 ,
         \rnd_reg/N10 , \rnd_reg/N9 , \rnd_reg/N8 , \rnd_reg/N7 , \rnd_reg/N6 ,
         \rnd_reg/N5 , \rnd_reg/N4 , \rnd_reg/N3 , \cv_next_reg/n320 ,
         \cv_next_reg/n310 , \cv_next_reg/n300 , \cv_next_reg/n290 ,
         \cv_next_reg/n280 , \cv_next_reg/n270 , \cv_next_reg/n260 ,
         \cv_next_reg/n250 , \cv_next_reg/n240 , \cv_next_reg/n230 ,
         \cv_next_reg/n220 , \cv_next_reg/n210 , \cv_next_reg/n200 ,
         \cv_next_reg/n190 , \cv_next_reg/n180 , \cv_next_reg/n170 ,
         \cv_next_reg/N162 , \cv_next_reg/N161 , \cv_next_reg/N160 ,
         \cv_next_reg/N159 , \cv_next_reg/N158 , \cv_next_reg/N157 ,
         \cv_next_reg/N156 , \cv_next_reg/N155 , \cv_next_reg/N154 ,
         \cv_next_reg/N153 , \cv_next_reg/N152 , \cv_next_reg/N151 ,
         \cv_next_reg/N150 , \cv_next_reg/N149 , \cv_next_reg/N148 ,
         \cv_next_reg/N147 , \cv_next_reg/N146 , \cv_next_reg/N145 ,
         \cv_next_reg/N144 , \cv_next_reg/N143 , \cv_next_reg/N142 ,
         \cv_next_reg/N141 , \cv_next_reg/N140 , \cv_next_reg/N139 ,
         \cv_next_reg/N138 , \cv_next_reg/N137 , \cv_next_reg/N136 ,
         \cv_next_reg/N135 , \cv_next_reg/N134 , \cv_next_reg/N133 ,
         \cv_next_reg/N132 , \cv_next_reg/N131 , \cv_next_reg/N130 ,
         \cv_next_reg/N129 , \cv_next_reg/N128 , \cv_next_reg/N127 ,
         \cv_next_reg/N126 , \cv_next_reg/N125 , \cv_next_reg/N124 ,
         \cv_next_reg/N123 , \cv_next_reg/N122 , \cv_next_reg/N121 ,
         \cv_next_reg/N120 , \cv_next_reg/N119 , \cv_next_reg/N118 ,
         \cv_next_reg/N117 , \cv_next_reg/N116 , \cv_next_reg/N115 ,
         \cv_next_reg/N114 , \cv_next_reg/N113 , \cv_next_reg/N112 ,
         \cv_next_reg/N111 , \cv_next_reg/N110 , \cv_next_reg/N109 ,
         \cv_next_reg/N108 , \cv_next_reg/N107 , \cv_next_reg/N106 ,
         \cv_next_reg/N105 , \cv_next_reg/N104 , \cv_next_reg/N103 ,
         \cv_next_reg/N102 , \cv_next_reg/N101 , \cv_next_reg/N100 ,
         \cv_next_reg/N99 , \cv_next_reg/N98 , \cv_next_reg/N97 ,
         \cv_next_reg/N96 , \cv_next_reg/N95 , \cv_next_reg/N94 ,
         \cv_next_reg/N93 , \cv_next_reg/N92 , \cv_next_reg/N91 ,
         \cv_next_reg/N90 , \cv_next_reg/N89 , \cv_next_reg/N88 ,
         \cv_next_reg/N87 , \cv_next_reg/N86 , \cv_next_reg/N85 ,
         \cv_next_reg/N84 , \cv_next_reg/N83 , \cv_next_reg/N82 ,
         \cv_next_reg/N81 , \cv_next_reg/N80 , \cv_next_reg/N79 ,
         \cv_next_reg/N78 , \cv_next_reg/N77 , \cv_next_reg/N76 ,
         \cv_next_reg/N75 , \cv_next_reg/N74 , \cv_next_reg/N73 ,
         \cv_next_reg/N72 , \cv_next_reg/N71 , \cv_next_reg/N70 ,
         \cv_next_reg/N69 , \cv_next_reg/N68 , \cv_next_reg/N67 ,
         \cv_next_reg/N66 , \cv_next_reg/N65 , \cv_next_reg/N64 ,
         \cv_next_reg/N63 , \cv_next_reg/N62 , \cv_next_reg/N61 ,
         \cv_next_reg/N60 , \cv_next_reg/N59 , \cv_next_reg/N58 ,
         \cv_next_reg/N57 , \cv_next_reg/N56 , \cv_next_reg/N55 ,
         \cv_next_reg/N54 , \cv_next_reg/N53 , \cv_next_reg/N52 ,
         \cv_next_reg/N51 , \cv_next_reg/N50 , \cv_next_reg/N49 ,
         \cv_next_reg/N48 , \cv_next_reg/N47 , \cv_next_reg/N46 ,
         \cv_next_reg/N45 , \cv_next_reg/N44 , \cv_next_reg/N43 ,
         \cv_next_reg/N42 , \cv_next_reg/N41 , \cv_next_reg/N40 ,
         \cv_next_reg/N39 , \cv_next_reg/N38 , \cv_next_reg/N37 ,
         \cv_next_reg/N36 , \cv_next_reg/N35 , \cv_next_reg/N34 ,
         \cv_next_reg/N33 , \cv_next_reg/N32 , \cv_next_reg/N31 ,
         \cv_next_reg/N30 , \cv_next_reg/N29 , \cv_next_reg/N28 ,
         \cv_next_reg/N27 , \cv_next_reg/N26 , \cv_next_reg/N25 ,
         \cv_next_reg/N24 , \cv_next_reg/N23 , \cv_next_reg/N22 ,
         \cv_next_reg/N21 , \cv_next_reg/N20 , \cv_next_reg/N19 ,
         \cv_next_reg/N18 , \cv_next_reg/N17 , \cv_next_reg/N16 ,
         \cv_next_reg/N15 , \cv_next_reg/N14 , \cv_next_reg/N13 ,
         \cv_next_reg/N12 , \cv_next_reg/N11 , \cv_next_reg/N10 ,
         \cv_next_reg/N9 , \cv_next_reg/N8 , \cv_next_reg/N7 ,
         \cv_next_reg/N6 , \cv_next_reg/N5 , \cv_next_reg/N4 ,
         \cv_next_reg/N3 , \add_98_2/n379 , \add_98_2/n378 , \add_98_2/n377 ,
         \add_98_2/n376 , \add_98_2/n375 , \add_98_2/n374 , \add_98_2/n373 ,
         \add_98_2/n372 , \add_98_2/n371 , \add_98_2/n370 , \add_98_2/n369 ,
         \add_98_2/n368 , \add_98_2/n367 , \add_98_2/n366 , \add_98_2/n365 ,
         \add_98_2/n364 , \add_98_2/n363 , \add_98_2/n362 , \add_98_2/n361 ,
         \add_98_2/n360 , \add_98_2/n359 , \add_98_2/n358 , \add_98_2/n357 ,
         \add_98_2/n356 , \add_98_2/n355 , \add_98_2/n354 , \add_98_2/n353 ,
         \add_98_2/n352 , \add_98_2/n351 , \add_98_2/n350 , \add_98_2/n349 ,
         \add_98_2/n348 , \add_98_2/n347 , \add_98_2/n346 , \add_98_2/n345 ,
         \add_98_2/n344 , \add_98_2/n343 , \add_98_2/n342 , \add_98_2/n341 ,
         \add_98_2/n340 , \add_98_2/n339 , \add_98_2/n338 , \add_98_2/n337 ,
         \add_98_2/n336 , \add_98_2/n335 , \add_98_2/n334 , \add_98_2/n333 ,
         \add_98_2/n332 , \add_98_2/n331 , \add_98_2/n330 , \add_98_2/n329 ,
         \add_98_2/n328 , \add_98_2/n327 , \add_98_2/n326 , \add_98_2/n325 ,
         \add_98_2/n324 , \add_98_2/n323 , \add_98_2/n322 , \add_98_2/n321 ,
         \add_98_2/n320 , \add_98_2/n319 , \add_98_2/n318 , \add_98_2/n317 ,
         \add_98_2/n316 , \add_98_2/n315 , \add_98_2/n314 , \add_98_2/n313 ,
         \add_98_2/n312 , \add_98_2/n311 , \add_98_2/n310 , \add_98_2/n309 ,
         \add_98_2/n308 , \add_98_2/n307 , \add_98_2/n306 , \add_98_2/n305 ,
         \add_98_2/n304 , \add_98_2/n303 , \add_98_2/n302 , \add_98_2/n301 ,
         \add_98_2/n300 , \add_98_2/n299 , \add_98_2/n298 , \add_98_2/n297 ,
         \add_98_2/n296 , \add_98_2/n295 , \add_98_2/n294 , \add_98_2/n293 ,
         \add_98_2/n292 , \add_98_2/n291 , \add_98_2/n290 , \add_98_2/n289 ,
         \add_98_2/n288 , \add_98_2/n287 , \add_98_2/n286 , \add_98_2/n285 ,
         \add_98_2/n284 , \add_98_2/n283 , \add_98_2/n282 , \add_98_2/n281 ,
         \add_98_2/n280 , \add_98_2/n279 , \add_98_2/n278 , \add_98_2/n277 ,
         \add_98_2/n276 , \add_98_2/n275 , \add_98_2/n274 , \add_98_2/n273 ,
         \add_98_2/n272 , \add_98_2/n271 , \add_98_2/n270 , \add_98_2/n269 ,
         \add_98_2/n268 , \add_98_2/n267 , \add_98_2/n266 , \add_98_2/n265 ,
         \add_98_2/n264 , \add_98_2/n263 , \add_98_2/n262 , \add_98_2/n261 ,
         \add_98_2/n260 , \add_98_2/n259 , \add_98_2/n258 , \add_98_2/n257 ,
         \add_98_2/n256 , \add_98_2/n255 , \add_98_2/n254 , \add_98_2/n253 ,
         \add_98_2/n252 , \add_98_2/n251 , \add_98_2/n250 , \add_98_2/n249 ,
         \add_98_2/n248 , \add_98_2/n247 , \add_98_2/n246 , \add_98_2/n245 ,
         \add_98_2/n244 , \add_98_2/n243 , \add_98_2/n242 , \add_98_2/n241 ,
         \add_98_2/n240 , \add_98_2/n239 , \add_98_2/n238 , \add_98_2/n237 ,
         \add_98_2/n236 , \add_98_2/n235 , \add_98_2/n234 , \add_98_2/n233 ,
         \add_98_2/n232 , \add_98_2/n231 , \add_98_2/n230 , \add_98_2/n229 ,
         \add_98_2/n228 , \add_98_2/n227 , \add_98_2/n226 , \add_98_2/n225 ,
         \add_98_2/n224 , \add_98_2/n223 , \add_98_2/n222 , \add_98_2/n221 ,
         \add_98_2/n220 , \add_98_2/n219 , \add_98_2/n218 , \add_98_2/n217 ,
         \add_98_2/n216 , \add_98_2/n215 , \add_98_2/n214 , \add_98_2/n213 ,
         \add_98_2/n212 , \add_98_2/n211 , \add_98_2/n210 , \add_98_2/n209 ,
         \add_98_2/n208 , \add_98_2/n207 , \add_98_2/n206 , \add_98_2/n205 ,
         \add_98_2/n204 , \add_98_2/n203 , \add_98_2/n202 , \add_98_2/n201 ,
         \add_98_2/n200 , \add_98_2/n199 , \add_98_2/n198 , \add_98_2/n197 ,
         \add_98_2/n196 , \add_98_2/n195 , \add_98_2/n194 , \add_98_2/n193 ,
         \add_98_2/n192 , \add_98_2/n191 , \add_98_2/n190 , \add_98_2/n189 ,
         \add_98_2/n188 , \add_98_2/n187 , \add_98_2/n186 , \add_98_2/n185 ,
         \add_98_2/n184 , \add_98_2/n183 , \add_98_2/n182 , \add_98_2/n181 ,
         \add_98_2/n180 , \add_98_2/n179 , \add_98_2/n178 , \add_98_2/n177 ,
         \add_98_2/n176 , \add_98_2/n175 , \add_98_2/n174 , \add_98_2/n173 ,
         \add_98_2/n172 , \add_98_2/n171 , \add_98_2/n170 , \add_98_2/n169 ,
         \add_98_2/n168 , \add_98_2/n167 , \add_98_2/n166 , \add_98_2/n165 ,
         \add_98_2/n164 , \add_98_2/n163 , \add_98_2/n162 , \add_98_2/n161 ,
         \add_98_2/n160 , \add_98_2/n159 , \add_98_2/n158 , \add_98_2/n157 ,
         \add_98_2/n156 , \add_98_2/n155 , \add_98_2/n154 , \add_98_2/n153 ,
         \add_98_2/n152 , \add_98_2/n151 , \add_98_2/n150 , \add_98_2/n149 ,
         \add_98_2/n148 , \add_98_2/n147 , \add_98_2/n146 , \add_98_2/n145 ,
         \add_98_2/n144 , \add_98_2/n143 , \add_98_2/n142 , \add_98_2/n141 ,
         \add_98_2/n140 , \add_98_2/n139 , \add_98_2/n138 , \add_98_2/n137 ,
         \add_98_2/n136 , \add_98_2/n135 , \add_98_2/n134 , \add_98_2/n133 ,
         \add_98_2/n132 , \add_98_2/n131 , \add_98_2/n130 , \add_98_2/n129 ,
         \add_98_2/n128 , \add_98_2/n127 , \add_98_2/n126 , \add_98_2/n125 ,
         \add_98_2/n124 , \add_98_2/n123 , \add_98_2/n122 , \add_98_2/n121 ,
         \add_98_2/n120 , \add_98_2/n119 , \add_98_2/n118 , \add_98_2/n117 ,
         \add_98_2/n116 , \add_98_2/n115 , \add_98_2/n114 , \add_98_2/n113 ,
         \add_98_2/n112 , \add_98_2/n111 , \add_98_2/n110 , \add_98_2/n109 ,
         \add_98_2/n108 , \add_98_2/n107 , \add_98_2/n106 , \add_98_2/n105 ,
         \add_98_2/n104 , \add_98_2/n103 , \add_98_2/n102 , \add_98_2/n101 ,
         \add_98_2/n100 , \add_98_2/n99 , \add_98_2/n98 , \add_98_2/n97 ,
         \add_98_2/n96 , \add_98_2/n95 , \add_98_2/n94 , \add_98_2/n93 ,
         \add_98_2/n92 , \add_98_2/n91 , \add_98_2/n90 , \add_98_2/n89 ,
         \add_98_2/n88 , \add_98_2/n87 , \add_98_2/n86 , \add_98_2/n85 ,
         \add_98_2/n84 , \add_98_2/n83 , \add_98_2/n82 , \add_98_2/n81 ,
         \add_98_2/n80 , \add_98_2/n79 , \add_98_2/n78 , \add_98_2/n77 ,
         \add_98_2/n76 , \add_98_2/n75 , \add_98_2/n74 , \add_98_2/n73 ,
         \add_98_2/n72 , \add_98_2/n71 , \add_98_2/n70 , \add_98_2/n69 ,
         \add_98_2/n68 , \add_98_2/n67 , \add_98_2/n66 , \add_98_2/n65 ,
         \add_98_2/n64 , \add_98_2/n63 , \add_98_2/n62 , \add_98_2/n61 ,
         \add_98_2/n60 , \add_98_2/n59 , \add_98_2/n58 , \add_98_2/n57 ,
         \add_98_2/n56 , \add_98_2/n55 , \add_98_2/n54 , \add_98_2/n53 ,
         \add_98_2/n52 , \add_98_2/n51 , \add_98_2/n50 , \add_98_2/n49 ,
         \add_98_2/n48 , \add_98_2/n47 , \add_98_2/n46 , \add_98_2/n45 ,
         \add_98_2/n44 , \add_98_2/n43 , \add_98_2/n42 , \add_98_2/n41 ,
         \add_98_2/n40 , \add_98_2/n39 , \add_98_2/n38 , \add_98_2/n37 ,
         \add_98_2/n36 , \add_98_2/n35 , \add_98_2/n34 , \add_98_2/n33 ,
         \add_98_2/n32 , \add_98_2/n31 , \add_98_2/n30 , \add_98_2/n29 ,
         \add_98_2/n28 , \add_98_2/n26 , \add_98_2/n25 , \add_98_2/n24 ,
         \add_98_2/n23 , \add_98_2/n22 , \add_98_2/n21 , \add_98_2/n20 ,
         \add_98_2/n19 , \add_98_2/n18 , \add_98_2/n17 , \add_98_2/n16 ,
         \add_98_2/n15 , \add_98_2/n14 , \add_98_2/n13 , \add_98_2/n12 ,
         \add_98_2/n11 , \add_98_2/n10 , \add_98_2/n9 , \add_98_2/n8 ,
         \add_98_2/n7 , \add_98_2/n6 , \add_98_2/n5 , \add_98_2/n4 ,
         \add_98_2/n3 , \add_98_2/n2 , \add_98_2/n1 , \add_98_3/n381 ,
         \add_98_3/n380 , \add_98_3/n379 , \add_98_3/n378 , \add_98_3/n377 ,
         \add_98_3/n376 , \add_98_3/n375 , \add_98_3/n374 , \add_98_3/n373 ,
         \add_98_3/n372 , \add_98_3/n371 , \add_98_3/n370 , \add_98_3/n369 ,
         \add_98_3/n368 , \add_98_3/n367 , \add_98_3/n366 , \add_98_3/n365 ,
         \add_98_3/n364 , \add_98_3/n363 , \add_98_3/n362 , \add_98_3/n361 ,
         \add_98_3/n360 , \add_98_3/n359 , \add_98_3/n358 , \add_98_3/n357 ,
         \add_98_3/n356 , \add_98_3/n355 , \add_98_3/n354 , \add_98_3/n353 ,
         \add_98_3/n352 , \add_98_3/n351 , \add_98_3/n350 , \add_98_3/n349 ,
         \add_98_3/n348 , \add_98_3/n347 , \add_98_3/n346 , \add_98_3/n345 ,
         \add_98_3/n344 , \add_98_3/n343 , \add_98_3/n342 , \add_98_3/n341 ,
         \add_98_3/n340 , \add_98_3/n339 , \add_98_3/n338 , \add_98_3/n337 ,
         \add_98_3/n336 , \add_98_3/n335 , \add_98_3/n334 , \add_98_3/n333 ,
         \add_98_3/n332 , \add_98_3/n331 , \add_98_3/n330 , \add_98_3/n329 ,
         \add_98_3/n328 , \add_98_3/n327 , \add_98_3/n326 , \add_98_3/n325 ,
         \add_98_3/n324 , \add_98_3/n323 , \add_98_3/n322 , \add_98_3/n321 ,
         \add_98_3/n320 , \add_98_3/n319 , \add_98_3/n318 , \add_98_3/n317 ,
         \add_98_3/n316 , \add_98_3/n315 , \add_98_3/n314 , \add_98_3/n313 ,
         \add_98_3/n312 , \add_98_3/n311 , \add_98_3/n310 , \add_98_3/n309 ,
         \add_98_3/n308 , \add_98_3/n307 , \add_98_3/n306 , \add_98_3/n305 ,
         \add_98_3/n304 , \add_98_3/n303 , \add_98_3/n302 , \add_98_3/n301 ,
         \add_98_3/n300 , \add_98_3/n299 , \add_98_3/n298 , \add_98_3/n297 ,
         \add_98_3/n296 , \add_98_3/n295 , \add_98_3/n294 , \add_98_3/n293 ,
         \add_98_3/n292 , \add_98_3/n291 , \add_98_3/n290 , \add_98_3/n289 ,
         \add_98_3/n288 , \add_98_3/n287 , \add_98_3/n286 , \add_98_3/n285 ,
         \add_98_3/n284 , \add_98_3/n283 , \add_98_3/n282 , \add_98_3/n281 ,
         \add_98_3/n280 , \add_98_3/n279 , \add_98_3/n278 , \add_98_3/n277 ,
         \add_98_3/n276 , \add_98_3/n275 , \add_98_3/n274 , \add_98_3/n273 ,
         \add_98_3/n272 , \add_98_3/n271 , \add_98_3/n270 , \add_98_3/n269 ,
         \add_98_3/n268 , \add_98_3/n267 , \add_98_3/n266 , \add_98_3/n265 ,
         \add_98_3/n264 , \add_98_3/n263 , \add_98_3/n262 , \add_98_3/n261 ,
         \add_98_3/n260 , \add_98_3/n259 , \add_98_3/n258 , \add_98_3/n257 ,
         \add_98_3/n256 , \add_98_3/n255 , \add_98_3/n254 , \add_98_3/n253 ,
         \add_98_3/n252 , \add_98_3/n251 , \add_98_3/n250 , \add_98_3/n249 ,
         \add_98_3/n248 , \add_98_3/n247 , \add_98_3/n246 , \add_98_3/n245 ,
         \add_98_3/n244 , \add_98_3/n243 , \add_98_3/n242 , \add_98_3/n241 ,
         \add_98_3/n240 , \add_98_3/n239 , \add_98_3/n238 , \add_98_3/n237 ,
         \add_98_3/n236 , \add_98_3/n235 , \add_98_3/n234 , \add_98_3/n233 ,
         \add_98_3/n232 , \add_98_3/n231 , \add_98_3/n230 , \add_98_3/n229 ,
         \add_98_3/n228 , \add_98_3/n227 , \add_98_3/n226 , \add_98_3/n225 ,
         \add_98_3/n224 , \add_98_3/n223 , \add_98_3/n222 , \add_98_3/n221 ,
         \add_98_3/n220 , \add_98_3/n219 , \add_98_3/n218 , \add_98_3/n217 ,
         \add_98_3/n216 , \add_98_3/n215 , \add_98_3/n214 , \add_98_3/n213 ,
         \add_98_3/n212 , \add_98_3/n211 , \add_98_3/n210 , \add_98_3/n209 ,
         \add_98_3/n208 , \add_98_3/n207 , \add_98_3/n206 , \add_98_3/n205 ,
         \add_98_3/n204 , \add_98_3/n203 , \add_98_3/n202 , \add_98_3/n201 ,
         \add_98_3/n200 , \add_98_3/n199 , \add_98_3/n198 , \add_98_3/n197 ,
         \add_98_3/n196 , \add_98_3/n195 , \add_98_3/n194 , \add_98_3/n193 ,
         \add_98_3/n192 , \add_98_3/n191 , \add_98_3/n190 , \add_98_3/n189 ,
         \add_98_3/n188 , \add_98_3/n187 , \add_98_3/n186 , \add_98_3/n185 ,
         \add_98_3/n184 , \add_98_3/n183 , \add_98_3/n182 , \add_98_3/n181 ,
         \add_98_3/n180 , \add_98_3/n179 , \add_98_3/n178 , \add_98_3/n177 ,
         \add_98_3/n176 , \add_98_3/n175 , \add_98_3/n174 , \add_98_3/n173 ,
         \add_98_3/n172 , \add_98_3/n171 , \add_98_3/n170 , \add_98_3/n169 ,
         \add_98_3/n168 , \add_98_3/n167 , \add_98_3/n166 , \add_98_3/n165 ,
         \add_98_3/n164 , \add_98_3/n163 , \add_98_3/n162 , \add_98_3/n161 ,
         \add_98_3/n160 , \add_98_3/n159 , \add_98_3/n158 , \add_98_3/n157 ,
         \add_98_3/n156 , \add_98_3/n155 , \add_98_3/n154 , \add_98_3/n153 ,
         \add_98_3/n152 , \add_98_3/n151 , \add_98_3/n150 , \add_98_3/n149 ,
         \add_98_3/n148 , \add_98_3/n147 , \add_98_3/n146 , \add_98_3/n145 ,
         \add_98_3/n144 , \add_98_3/n143 , \add_98_3/n142 , \add_98_3/n141 ,
         \add_98_3/n140 , \add_98_3/n139 , \add_98_3/n138 , \add_98_3/n137 ,
         \add_98_3/n136 , \add_98_3/n135 , \add_98_3/n134 , \add_98_3/n133 ,
         \add_98_3/n132 , \add_98_3/n131 , \add_98_3/n130 , \add_98_3/n129 ,
         \add_98_3/n128 , \add_98_3/n127 , \add_98_3/n126 , \add_98_3/n125 ,
         \add_98_3/n124 , \add_98_3/n123 , \add_98_3/n122 , \add_98_3/n121 ,
         \add_98_3/n120 , \add_98_3/n119 , \add_98_3/n118 , \add_98_3/n117 ,
         \add_98_3/n116 , \add_98_3/n115 , \add_98_3/n114 , \add_98_3/n113 ,
         \add_98_3/n112 , \add_98_3/n111 , \add_98_3/n110 , \add_98_3/n109 ,
         \add_98_3/n108 , \add_98_3/n107 , \add_98_3/n106 , \add_98_3/n105 ,
         \add_98_3/n104 , \add_98_3/n103 , \add_98_3/n102 , \add_98_3/n101 ,
         \add_98_3/n100 , \add_98_3/n99 , \add_98_3/n98 , \add_98_3/n97 ,
         \add_98_3/n96 , \add_98_3/n95 , \add_98_3/n94 , \add_98_3/n93 ,
         \add_98_3/n92 , \add_98_3/n91 , \add_98_3/n90 , \add_98_3/n89 ,
         \add_98_3/n88 , \add_98_3/n87 , \add_98_3/n86 , \add_98_3/n85 ,
         \add_98_3/n84 , \add_98_3/n83 , \add_98_3/n82 , \add_98_3/n81 ,
         \add_98_3/n80 , \add_98_3/n79 , \add_98_3/n78 , \add_98_3/n77 ,
         \add_98_3/n76 , \add_98_3/n75 , \add_98_3/n74 , \add_98_3/n73 ,
         \add_98_3/n72 , \add_98_3/n71 , \add_98_3/n70 , \add_98_3/n69 ,
         \add_98_3/n68 , \add_98_3/n67 , \add_98_3/n66 , \add_98_3/n65 ,
         \add_98_3/n64 , \add_98_3/n63 , \add_98_3/n62 , \add_98_3/n61 ,
         \add_98_3/n60 , \add_98_3/n59 , \add_98_3/n58 , \add_98_3/n57 ,
         \add_98_3/n56 , \add_98_3/n55 , \add_98_3/n54 , \add_98_3/n53 ,
         \add_98_3/n52 , \add_98_3/n51 , \add_98_3/n50 , \add_98_3/n49 ,
         \add_98_3/n48 , \add_98_3/n47 , \add_98_3/n46 , \add_98_3/n45 ,
         \add_98_3/n44 , \add_98_3/n43 , \add_98_3/n42 , \add_98_3/n41 ,
         \add_98_3/n40 , \add_98_3/n39 , \add_98_3/n38 , \add_98_3/n37 ,
         \add_98_3/n36 , \add_98_3/n35 , \add_98_3/n34 , \add_98_3/n33 ,
         \add_98_3/n32 , \add_98_3/n31 , \add_98_3/n30 , \add_98_3/n29 ,
         \add_98_3/n28 , \add_98_3/n26 , \add_98_3/n25 , \add_98_3/n24 ,
         \add_98_3/n23 , \add_98_3/n22 , \add_98_3/n21 , \add_98_3/n20 ,
         \add_98_3/n19 , \add_98_3/n18 , \add_98_3/n17 , \add_98_3/n16 ,
         \add_98_3/n15 , \add_98_3/n14 , \add_98_3/n13 , \add_98_3/n12 ,
         \add_98_3/n11 , \add_98_3/n10 , \add_98_3/n9 , \add_98_3/n8 ,
         \add_98_3/n7 , \add_98_3/n6 , \add_98_3/n5 , \add_98_3/n4 ,
         \add_98_3/n3 , \add_98_3/n2 , \add_98_3/n1 , \add_98_5/n392 ,
         \add_98_5/n391 , \add_98_5/n390 , \add_98_5/n389 , \add_98_5/n388 ,
         \add_98_5/n387 , \add_98_5/n386 , \add_98_5/n385 , \add_98_5/n384 ,
         \add_98_5/n383 , \add_98_5/n382 , \add_98_5/n381 , \add_98_5/n380 ,
         \add_98_5/n379 , \add_98_5/n378 , \add_98_5/n377 , \add_98_5/n376 ,
         \add_98_5/n375 , \add_98_5/n374 , \add_98_5/n373 , \add_98_5/n372 ,
         \add_98_5/n371 , \add_98_5/n370 , \add_98_5/n369 , \add_98_5/n368 ,
         \add_98_5/n367 , \add_98_5/n366 , \add_98_5/n365 , \add_98_5/n364 ,
         \add_98_5/n363 , \add_98_5/n362 , \add_98_5/n361 , \add_98_5/n360 ,
         \add_98_5/n359 , \add_98_5/n358 , \add_98_5/n357 , \add_98_5/n356 ,
         \add_98_5/n355 , \add_98_5/n354 , \add_98_5/n353 , \add_98_5/n352 ,
         \add_98_5/n351 , \add_98_5/n350 , \add_98_5/n349 , \add_98_5/n348 ,
         \add_98_5/n347 , \add_98_5/n346 , \add_98_5/n345 , \add_98_5/n344 ,
         \add_98_5/n343 , \add_98_5/n342 , \add_98_5/n341 , \add_98_5/n340 ,
         \add_98_5/n339 , \add_98_5/n338 , \add_98_5/n337 , \add_98_5/n336 ,
         \add_98_5/n335 , \add_98_5/n334 , \add_98_5/n333 , \add_98_5/n332 ,
         \add_98_5/n331 , \add_98_5/n330 , \add_98_5/n329 , \add_98_5/n328 ,
         \add_98_5/n327 , \add_98_5/n326 , \add_98_5/n325 , \add_98_5/n324 ,
         \add_98_5/n323 , \add_98_5/n322 , \add_98_5/n321 , \add_98_5/n320 ,
         \add_98_5/n319 , \add_98_5/n318 , \add_98_5/n317 , \add_98_5/n316 ,
         \add_98_5/n315 , \add_98_5/n314 , \add_98_5/n313 , \add_98_5/n312 ,
         \add_98_5/n311 , \add_98_5/n310 , \add_98_5/n309 , \add_98_5/n308 ,
         \add_98_5/n307 , \add_98_5/n306 , \add_98_5/n305 , \add_98_5/n304 ,
         \add_98_5/n303 , \add_98_5/n302 , \add_98_5/n301 , \add_98_5/n300 ,
         \add_98_5/n299 , \add_98_5/n298 , \add_98_5/n297 , \add_98_5/n296 ,
         \add_98_5/n295 , \add_98_5/n294 , \add_98_5/n293 , \add_98_5/n292 ,
         \add_98_5/n291 , \add_98_5/n290 , \add_98_5/n289 , \add_98_5/n288 ,
         \add_98_5/n287 , \add_98_5/n286 , \add_98_5/n285 , \add_98_5/n284 ,
         \add_98_5/n283 , \add_98_5/n282 , \add_98_5/n281 , \add_98_5/n280 ,
         \add_98_5/n279 , \add_98_5/n278 , \add_98_5/n277 , \add_98_5/n276 ,
         \add_98_5/n275 , \add_98_5/n274 , \add_98_5/n273 , \add_98_5/n272 ,
         \add_98_5/n271 , \add_98_5/n270 , \add_98_5/n269 , \add_98_5/n268 ,
         \add_98_5/n267 , \add_98_5/n266 , \add_98_5/n265 , \add_98_5/n264 ,
         \add_98_5/n263 , \add_98_5/n262 , \add_98_5/n261 , \add_98_5/n260 ,
         \add_98_5/n259 , \add_98_5/n258 , \add_98_5/n257 , \add_98_5/n256 ,
         \add_98_5/n255 , \add_98_5/n254 , \add_98_5/n253 , \add_98_5/n252 ,
         \add_98_5/n251 , \add_98_5/n250 , \add_98_5/n249 , \add_98_5/n248 ,
         \add_98_5/n247 , \add_98_5/n246 , \add_98_5/n245 , \add_98_5/n244 ,
         \add_98_5/n243 , \add_98_5/n242 , \add_98_5/n241 , \add_98_5/n240 ,
         \add_98_5/n239 , \add_98_5/n238 , \add_98_5/n237 , \add_98_5/n236 ,
         \add_98_5/n235 , \add_98_5/n234 , \add_98_5/n233 , \add_98_5/n232 ,
         \add_98_5/n231 , \add_98_5/n230 , \add_98_5/n229 , \add_98_5/n228 ,
         \add_98_5/n227 , \add_98_5/n226 , \add_98_5/n225 , \add_98_5/n224 ,
         \add_98_5/n223 , \add_98_5/n222 , \add_98_5/n221 , \add_98_5/n220 ,
         \add_98_5/n219 , \add_98_5/n218 , \add_98_5/n217 , \add_98_5/n216 ,
         \add_98_5/n215 , \add_98_5/n214 , \add_98_5/n213 , \add_98_5/n212 ,
         \add_98_5/n211 , \add_98_5/n210 , \add_98_5/n209 , \add_98_5/n208 ,
         \add_98_5/n207 , \add_98_5/n206 , \add_98_5/n205 , \add_98_5/n204 ,
         \add_98_5/n203 , \add_98_5/n202 , \add_98_5/n201 , \add_98_5/n200 ,
         \add_98_5/n199 , \add_98_5/n198 , \add_98_5/n197 , \add_98_5/n196 ,
         \add_98_5/n195 , \add_98_5/n194 , \add_98_5/n193 , \add_98_5/n192 ,
         \add_98_5/n191 , \add_98_5/n190 , \add_98_5/n189 , \add_98_5/n188 ,
         \add_98_5/n187 , \add_98_5/n186 , \add_98_5/n185 , \add_98_5/n184 ,
         \add_98_5/n183 , \add_98_5/n182 , \add_98_5/n181 , \add_98_5/n180 ,
         \add_98_5/n179 , \add_98_5/n178 , \add_98_5/n177 , \add_98_5/n176 ,
         \add_98_5/n175 , \add_98_5/n174 , \add_98_5/n173 , \add_98_5/n172 ,
         \add_98_5/n171 , \add_98_5/n170 , \add_98_5/n169 , \add_98_5/n168 ,
         \add_98_5/n167 , \add_98_5/n166 , \add_98_5/n165 , \add_98_5/n164 ,
         \add_98_5/n163 , \add_98_5/n162 , \add_98_5/n161 , \add_98_5/n160 ,
         \add_98_5/n159 , \add_98_5/n158 , \add_98_5/n157 , \add_98_5/n156 ,
         \add_98_5/n155 , \add_98_5/n154 , \add_98_5/n153 , \add_98_5/n152 ,
         \add_98_5/n151 , \add_98_5/n150 , \add_98_5/n149 , \add_98_5/n148 ,
         \add_98_5/n147 , \add_98_5/n146 , \add_98_5/n145 , \add_98_5/n144 ,
         \add_98_5/n143 , \add_98_5/n142 , \add_98_5/n141 , \add_98_5/n140 ,
         \add_98_5/n139 , \add_98_5/n138 , \add_98_5/n137 , \add_98_5/n136 ,
         \add_98_5/n135 , \add_98_5/n134 , \add_98_5/n133 , \add_98_5/n132 ,
         \add_98_5/n131 , \add_98_5/n130 , \add_98_5/n129 , \add_98_5/n128 ,
         \add_98_5/n127 , \add_98_5/n126 , \add_98_5/n125 , \add_98_5/n124 ,
         \add_98_5/n123 , \add_98_5/n122 , \add_98_5/n121 , \add_98_5/n120 ,
         \add_98_5/n119 , \add_98_5/n118 , \add_98_5/n117 , \add_98_5/n116 ,
         \add_98_5/n115 , \add_98_5/n114 , \add_98_5/n113 , \add_98_5/n112 ,
         \add_98_5/n111 , \add_98_5/n110 , \add_98_5/n109 , \add_98_5/n108 ,
         \add_98_5/n107 , \add_98_5/n106 , \add_98_5/n105 , \add_98_5/n104 ,
         \add_98_5/n103 , \add_98_5/n102 , \add_98_5/n101 , \add_98_5/n100 ,
         \add_98_5/n99 , \add_98_5/n98 , \add_98_5/n97 , \add_98_5/n96 ,
         \add_98_5/n95 , \add_98_5/n94 , \add_98_5/n93 , \add_98_5/n92 ,
         \add_98_5/n91 , \add_98_5/n90 , \add_98_5/n89 , \add_98_5/n88 ,
         \add_98_5/n87 , \add_98_5/n86 , \add_98_5/n85 , \add_98_5/n84 ,
         \add_98_5/n83 , \add_98_5/n82 , \add_98_5/n81 , \add_98_5/n80 ,
         \add_98_5/n79 , \add_98_5/n78 , \add_98_5/n77 , \add_98_5/n76 ,
         \add_98_5/n75 , \add_98_5/n74 , \add_98_5/n73 , \add_98_5/n72 ,
         \add_98_5/n71 , \add_98_5/n70 , \add_98_5/n69 , \add_98_5/n68 ,
         \add_98_5/n67 , \add_98_5/n66 , \add_98_5/n65 , \add_98_5/n64 ,
         \add_98_5/n63 , \add_98_5/n62 , \add_98_5/n61 , \add_98_5/n60 ,
         \add_98_5/n59 , \add_98_5/n58 , \add_98_5/n57 , \add_98_5/n56 ,
         \add_98_5/n55 , \add_98_5/n54 , \add_98_5/n53 , \add_98_5/n52 ,
         \add_98_5/n51 , \add_98_5/n50 , \add_98_5/n49 , \add_98_5/n48 ,
         \add_98_5/n47 , \add_98_5/n46 , \add_98_5/n45 , \add_98_5/n44 ,
         \add_98_5/n43 , \add_98_5/n42 , \add_98_5/n41 , \add_98_5/n40 ,
         \add_98_5/n39 , \add_98_5/n38 , \add_98_5/n37 , \add_98_5/n36 ,
         \add_98_5/n35 , \add_98_5/n34 , \add_98_5/n33 , \add_98_5/n32 ,
         \add_98_5/n31 , \add_98_5/n29 , \add_98_5/n28 , \add_98_5/n27 ,
         \add_98_5/n26 , \add_98_5/n25 , \add_98_5/n24 , \add_98_5/n23 ,
         \add_98_5/n22 , \add_98_5/n21 , \add_98_5/n20 , \add_98_5/n19 ,
         \add_98_5/n18 , \add_98_5/n17 , \add_98_5/n16 , \add_98_5/n15 ,
         \add_98_5/n14 , \add_98_5/n13 , \add_98_5/n12 , \add_98_5/n11 ,
         \add_98_5/n10 , \add_98_5/n9 , \add_98_5/n8 , \add_98_5/n7 ,
         \add_98_5/n6 , \add_98_5/n5 , \add_98_5/n4 , \add_98_5/n3 ,
         \add_98_5/n2 , \add_98_5/n1 , \add_98/n394 , \add_98/n393 ,
         \add_98/n392 , \add_98/n391 , \add_98/n390 , \add_98/n389 ,
         \add_98/n388 , \add_98/n387 , \add_98/n386 , \add_98/n385 ,
         \add_98/n384 , \add_98/n383 , \add_98/n382 , \add_98/n381 ,
         \add_98/n380 , \add_98/n379 , \add_98/n378 , \add_98/n377 ,
         \add_98/n376 , \add_98/n375 , \add_98/n374 , \add_98/n373 ,
         \add_98/n372 , \add_98/n371 , \add_98/n370 , \add_98/n369 ,
         \add_98/n368 , \add_98/n367 , \add_98/n366 , \add_98/n365 ,
         \add_98/n364 , \add_98/n363 , \add_98/n362 , \add_98/n361 ,
         \add_98/n360 , \add_98/n359 , \add_98/n358 , \add_98/n357 ,
         \add_98/n356 , \add_98/n355 , \add_98/n354 , \add_98/n353 ,
         \add_98/n352 , \add_98/n351 , \add_98/n350 , \add_98/n349 ,
         \add_98/n348 , \add_98/n347 , \add_98/n346 , \add_98/n345 ,
         \add_98/n344 , \add_98/n343 , \add_98/n342 , \add_98/n341 ,
         \add_98/n340 , \add_98/n339 , \add_98/n338 , \add_98/n337 ,
         \add_98/n336 , \add_98/n335 , \add_98/n334 , \add_98/n333 ,
         \add_98/n332 , \add_98/n331 , \add_98/n330 , \add_98/n329 ,
         \add_98/n328 , \add_98/n327 , \add_98/n326 , \add_98/n325 ,
         \add_98/n324 , \add_98/n323 , \add_98/n322 , \add_98/n321 ,
         \add_98/n320 , \add_98/n319 , \add_98/n318 , \add_98/n317 ,
         \add_98/n316 , \add_98/n315 , \add_98/n314 , \add_98/n313 ,
         \add_98/n312 , \add_98/n311 , \add_98/n310 , \add_98/n309 ,
         \add_98/n308 , \add_98/n307 , \add_98/n306 , \add_98/n305 ,
         \add_98/n304 , \add_98/n303 , \add_98/n302 , \add_98/n301 ,
         \add_98/n300 , \add_98/n299 , \add_98/n298 , \add_98/n297 ,
         \add_98/n296 , \add_98/n295 , \add_98/n294 , \add_98/n293 ,
         \add_98/n292 , \add_98/n291 , \add_98/n290 , \add_98/n289 ,
         \add_98/n288 , \add_98/n287 , \add_98/n286 , \add_98/n285 ,
         \add_98/n284 , \add_98/n283 , \add_98/n282 , \add_98/n281 ,
         \add_98/n280 , \add_98/n279 , \add_98/n278 , \add_98/n277 ,
         \add_98/n276 , \add_98/n275 , \add_98/n274 , \add_98/n273 ,
         \add_98/n272 , \add_98/n271 , \add_98/n270 , \add_98/n269 ,
         \add_98/n268 , \add_98/n267 , \add_98/n266 , \add_98/n265 ,
         \add_98/n264 , \add_98/n263 , \add_98/n262 , \add_98/n261 ,
         \add_98/n260 , \add_98/n259 , \add_98/n258 , \add_98/n257 ,
         \add_98/n256 , \add_98/n255 , \add_98/n254 , \add_98/n253 ,
         \add_98/n252 , \add_98/n251 , \add_98/n250 , \add_98/n249 ,
         \add_98/n248 , \add_98/n247 , \add_98/n246 , \add_98/n245 ,
         \add_98/n244 , \add_98/n243 , \add_98/n242 , \add_98/n241 ,
         \add_98/n240 , \add_98/n239 , \add_98/n238 , \add_98/n237 ,
         \add_98/n236 , \add_98/n235 , \add_98/n234 , \add_98/n233 ,
         \add_98/n232 , \add_98/n231 , \add_98/n230 , \add_98/n229 ,
         \add_98/n228 , \add_98/n227 , \add_98/n226 , \add_98/n225 ,
         \add_98/n224 , \add_98/n223 , \add_98/n222 , \add_98/n221 ,
         \add_98/n220 , \add_98/n219 , \add_98/n218 , \add_98/n217 ,
         \add_98/n216 , \add_98/n215 , \add_98/n214 , \add_98/n213 ,
         \add_98/n212 , \add_98/n211 , \add_98/n210 , \add_98/n209 ,
         \add_98/n208 , \add_98/n207 , \add_98/n206 , \add_98/n205 ,
         \add_98/n204 , \add_98/n203 , \add_98/n202 , \add_98/n201 ,
         \add_98/n200 , \add_98/n199 , \add_98/n198 , \add_98/n197 ,
         \add_98/n196 , \add_98/n195 , \add_98/n194 , \add_98/n193 ,
         \add_98/n192 , \add_98/n191 , \add_98/n190 , \add_98/n189 ,
         \add_98/n188 , \add_98/n187 , \add_98/n186 , \add_98/n185 ,
         \add_98/n184 , \add_98/n183 , \add_98/n182 , \add_98/n181 ,
         \add_98/n180 , \add_98/n179 , \add_98/n178 , \add_98/n177 ,
         \add_98/n176 , \add_98/n175 , \add_98/n174 , \add_98/n173 ,
         \add_98/n172 , \add_98/n171 , \add_98/n170 , \add_98/n169 ,
         \add_98/n168 , \add_98/n167 , \add_98/n166 , \add_98/n165 ,
         \add_98/n164 , \add_98/n163 , \add_98/n162 , \add_98/n161 ,
         \add_98/n160 , \add_98/n159 , \add_98/n158 , \add_98/n157 ,
         \add_98/n156 , \add_98/n155 , \add_98/n154 , \add_98/n153 ,
         \add_98/n152 , \add_98/n151 , \add_98/n150 , \add_98/n149 ,
         \add_98/n148 , \add_98/n147 , \add_98/n146 , \add_98/n145 ,
         \add_98/n144 , \add_98/n143 , \add_98/n142 , \add_98/n141 ,
         \add_98/n140 , \add_98/n139 , \add_98/n138 , \add_98/n137 ,
         \add_98/n136 , \add_98/n135 , \add_98/n134 , \add_98/n133 ,
         \add_98/n132 , \add_98/n131 , \add_98/n130 , \add_98/n129 ,
         \add_98/n128 , \add_98/n127 , \add_98/n126 , \add_98/n125 ,
         \add_98/n124 , \add_98/n123 , \add_98/n122 , \add_98/n121 ,
         \add_98/n120 , \add_98/n119 , \add_98/n118 , \add_98/n117 ,
         \add_98/n116 , \add_98/n115 , \add_98/n114 , \add_98/n113 ,
         \add_98/n112 , \add_98/n111 , \add_98/n110 , \add_98/n109 ,
         \add_98/n108 , \add_98/n107 , \add_98/n106 , \add_98/n105 ,
         \add_98/n104 , \add_98/n103 , \add_98/n102 , \add_98/n101 ,
         \add_98/n100 , \add_98/n99 , \add_98/n98 , \add_98/n97 , \add_98/n96 ,
         \add_98/n95 , \add_98/n94 , \add_98/n93 , \add_98/n92 , \add_98/n91 ,
         \add_98/n90 , \add_98/n89 , \add_98/n88 , \add_98/n87 , \add_98/n86 ,
         \add_98/n85 , \add_98/n84 , \add_98/n83 , \add_98/n82 , \add_98/n81 ,
         \add_98/n80 , \add_98/n79 , \add_98/n78 , \add_98/n77 , \add_98/n76 ,
         \add_98/n75 , \add_98/n74 , \add_98/n73 , \add_98/n72 , \add_98/n71 ,
         \add_98/n70 , \add_98/n69 , \add_98/n68 , \add_98/n67 , \add_98/n66 ,
         \add_98/n65 , \add_98/n64 , \add_98/n63 , \add_98/n62 , \add_98/n61 ,
         \add_98/n60 , \add_98/n59 , \add_98/n58 , \add_98/n57 , \add_98/n56 ,
         \add_98/n55 , \add_98/n54 , \add_98/n53 , \add_98/n52 , \add_98/n51 ,
         \add_98/n50 , \add_98/n49 , \add_98/n48 , \add_98/n47 , \add_98/n46 ,
         \add_98/n45 , \add_98/n44 , \add_98/n43 , \add_98/n42 , \add_98/n41 ,
         \add_98/n40 , \add_98/n39 , \add_98/n38 , \add_98/n37 , \add_98/n36 ,
         \add_98/n35 , \add_98/n34 , \add_98/n32 , \add_98/n31 , \add_98/n30 ,
         \add_98/n29 , \add_98/n28 , \add_98/n27 , \add_98/n26 , \add_98/n25 ,
         \add_98/n24 , \add_98/n23 , \add_98/n22 , \add_98/n21 , \add_98/n20 ,
         \add_98/n19 , \add_98/n18 , \add_98/n17 , \add_98/n16 , \add_98/n15 ,
         \add_98/n14 , \add_98/n13 , \add_98/n12 , \add_98/n11 , \add_98/n10 ,
         \add_98/n9 , \add_98/n8 , \add_98/n7 , \add_98/n6 , \add_98/n5 ,
         \add_98/n4 , \add_98/n3 , \add_98/n2 , \add_98/n1 , \add_98_4/n389 ,
         \add_98_4/n388 , \add_98_4/n387 , \add_98_4/n386 , \add_98_4/n385 ,
         \add_98_4/n384 , \add_98_4/n383 , \add_98_4/n382 , \add_98_4/n381 ,
         \add_98_4/n380 , \add_98_4/n379 , \add_98_4/n378 , \add_98_4/n377 ,
         \add_98_4/n376 , \add_98_4/n375 , \add_98_4/n374 , \add_98_4/n373 ,
         \add_98_4/n372 , \add_98_4/n371 , \add_98_4/n370 , \add_98_4/n369 ,
         \add_98_4/n368 , \add_98_4/n367 , \add_98_4/n366 , \add_98_4/n365 ,
         \add_98_4/n364 , \add_98_4/n363 , \add_98_4/n362 , \add_98_4/n361 ,
         \add_98_4/n360 , \add_98_4/n359 , \add_98_4/n358 , \add_98_4/n357 ,
         \add_98_4/n356 , \add_98_4/n355 , \add_98_4/n354 , \add_98_4/n353 ,
         \add_98_4/n352 , \add_98_4/n351 , \add_98_4/n350 , \add_98_4/n349 ,
         \add_98_4/n348 , \add_98_4/n347 , \add_98_4/n346 , \add_98_4/n345 ,
         \add_98_4/n344 , \add_98_4/n343 , \add_98_4/n342 , \add_98_4/n341 ,
         \add_98_4/n340 , \add_98_4/n339 , \add_98_4/n338 , \add_98_4/n337 ,
         \add_98_4/n336 , \add_98_4/n335 , \add_98_4/n334 , \add_98_4/n333 ,
         \add_98_4/n332 , \add_98_4/n331 , \add_98_4/n330 , \add_98_4/n329 ,
         \add_98_4/n328 , \add_98_4/n327 , \add_98_4/n326 , \add_98_4/n325 ,
         \add_98_4/n324 , \add_98_4/n323 , \add_98_4/n322 , \add_98_4/n321 ,
         \add_98_4/n320 , \add_98_4/n319 , \add_98_4/n318 , \add_98_4/n317 ,
         \add_98_4/n316 , \add_98_4/n315 , \add_98_4/n314 , \add_98_4/n313 ,
         \add_98_4/n312 , \add_98_4/n311 , \add_98_4/n310 , \add_98_4/n309 ,
         \add_98_4/n308 , \add_98_4/n307 , \add_98_4/n306 , \add_98_4/n305 ,
         \add_98_4/n304 , \add_98_4/n303 , \add_98_4/n302 , \add_98_4/n301 ,
         \add_98_4/n300 , \add_98_4/n299 , \add_98_4/n298 , \add_98_4/n297 ,
         \add_98_4/n296 , \add_98_4/n295 , \add_98_4/n294 , \add_98_4/n293 ,
         \add_98_4/n292 , \add_98_4/n291 , \add_98_4/n290 , \add_98_4/n289 ,
         \add_98_4/n288 , \add_98_4/n287 , \add_98_4/n286 , \add_98_4/n285 ,
         \add_98_4/n284 , \add_98_4/n283 , \add_98_4/n282 , \add_98_4/n281 ,
         \add_98_4/n280 , \add_98_4/n279 , \add_98_4/n278 , \add_98_4/n277 ,
         \add_98_4/n276 , \add_98_4/n275 , \add_98_4/n274 , \add_98_4/n273 ,
         \add_98_4/n272 , \add_98_4/n271 , \add_98_4/n270 , \add_98_4/n269 ,
         \add_98_4/n268 , \add_98_4/n267 , \add_98_4/n266 , \add_98_4/n265 ,
         \add_98_4/n264 , \add_98_4/n263 , \add_98_4/n262 , \add_98_4/n261 ,
         \add_98_4/n260 , \add_98_4/n259 , \add_98_4/n258 , \add_98_4/n257 ,
         \add_98_4/n256 , \add_98_4/n255 , \add_98_4/n254 , \add_98_4/n253 ,
         \add_98_4/n252 , \add_98_4/n251 , \add_98_4/n250 , \add_98_4/n249 ,
         \add_98_4/n248 , \add_98_4/n247 , \add_98_4/n246 , \add_98_4/n245 ,
         \add_98_4/n244 , \add_98_4/n243 , \add_98_4/n242 , \add_98_4/n241 ,
         \add_98_4/n240 , \add_98_4/n239 , \add_98_4/n238 , \add_98_4/n237 ,
         \add_98_4/n236 , \add_98_4/n235 , \add_98_4/n234 , \add_98_4/n233 ,
         \add_98_4/n232 , \add_98_4/n231 , \add_98_4/n230 , \add_98_4/n229 ,
         \add_98_4/n228 , \add_98_4/n227 , \add_98_4/n226 , \add_98_4/n225 ,
         \add_98_4/n224 , \add_98_4/n223 , \add_98_4/n222 , \add_98_4/n221 ,
         \add_98_4/n220 , \add_98_4/n219 , \add_98_4/n218 , \add_98_4/n217 ,
         \add_98_4/n216 , \add_98_4/n215 , \add_98_4/n214 , \add_98_4/n213 ,
         \add_98_4/n212 , \add_98_4/n211 , \add_98_4/n210 , \add_98_4/n209 ,
         \add_98_4/n208 , \add_98_4/n207 , \add_98_4/n206 , \add_98_4/n205 ,
         \add_98_4/n204 , \add_98_4/n203 , \add_98_4/n202 , \add_98_4/n201 ,
         \add_98_4/n200 , \add_98_4/n199 , \add_98_4/n198 , \add_98_4/n197 ,
         \add_98_4/n196 , \add_98_4/n195 , \add_98_4/n194 , \add_98_4/n193 ,
         \add_98_4/n192 , \add_98_4/n191 , \add_98_4/n190 , \add_98_4/n189 ,
         \add_98_4/n188 , \add_98_4/n187 , \add_98_4/n186 , \add_98_4/n185 ,
         \add_98_4/n184 , \add_98_4/n183 , \add_98_4/n182 , \add_98_4/n181 ,
         \add_98_4/n180 , \add_98_4/n179 , \add_98_4/n178 , \add_98_4/n177 ,
         \add_98_4/n176 , \add_98_4/n175 , \add_98_4/n174 , \add_98_4/n173 ,
         \add_98_4/n172 , \add_98_4/n171 , \add_98_4/n170 , \add_98_4/n169 ,
         \add_98_4/n168 , \add_98_4/n167 , \add_98_4/n166 , \add_98_4/n165 ,
         \add_98_4/n164 , \add_98_4/n163 , \add_98_4/n162 , \add_98_4/n161 ,
         \add_98_4/n160 , \add_98_4/n159 , \add_98_4/n158 , \add_98_4/n157 ,
         \add_98_4/n156 , \add_98_4/n155 , \add_98_4/n154 , \add_98_4/n153 ,
         \add_98_4/n152 , \add_98_4/n151 , \add_98_4/n150 , \add_98_4/n149 ,
         \add_98_4/n148 , \add_98_4/n147 , \add_98_4/n146 , \add_98_4/n145 ,
         \add_98_4/n144 , \add_98_4/n143 , \add_98_4/n142 , \add_98_4/n141 ,
         \add_98_4/n140 , \add_98_4/n139 , \add_98_4/n138 , \add_98_4/n137 ,
         \add_98_4/n136 , \add_98_4/n135 , \add_98_4/n134 , \add_98_4/n133 ,
         \add_98_4/n132 , \add_98_4/n131 , \add_98_4/n130 , \add_98_4/n129 ,
         \add_98_4/n128 , \add_98_4/n127 , \add_98_4/n126 , \add_98_4/n125 ,
         \add_98_4/n124 , \add_98_4/n123 , \add_98_4/n122 , \add_98_4/n121 ,
         \add_98_4/n120 , \add_98_4/n119 , \add_98_4/n118 , \add_98_4/n117 ,
         \add_98_4/n116 , \add_98_4/n115 , \add_98_4/n114 , \add_98_4/n113 ,
         \add_98_4/n112 , \add_98_4/n111 , \add_98_4/n110 , \add_98_4/n109 ,
         \add_98_4/n108 , \add_98_4/n107 , \add_98_4/n106 , \add_98_4/n105 ,
         \add_98_4/n104 , \add_98_4/n103 , \add_98_4/n102 , \add_98_4/n101 ,
         \add_98_4/n100 , \add_98_4/n99 , \add_98_4/n98 , \add_98_4/n97 ,
         \add_98_4/n96 , \add_98_4/n95 , \add_98_4/n94 , \add_98_4/n93 ,
         \add_98_4/n92 , \add_98_4/n91 , \add_98_4/n90 , \add_98_4/n89 ,
         \add_98_4/n88 , \add_98_4/n87 , \add_98_4/n86 , \add_98_4/n85 ,
         \add_98_4/n84 , \add_98_4/n83 , \add_98_4/n82 , \add_98_4/n81 ,
         \add_98_4/n80 , \add_98_4/n79 , \add_98_4/n78 , \add_98_4/n77 ,
         \add_98_4/n76 , \add_98_4/n75 , \add_98_4/n74 , \add_98_4/n73 ,
         \add_98_4/n72 , \add_98_4/n71 , \add_98_4/n70 , \add_98_4/n69 ,
         \add_98_4/n68 , \add_98_4/n67 , \add_98_4/n66 , \add_98_4/n65 ,
         \add_98_4/n64 , \add_98_4/n63 , \add_98_4/n62 , \add_98_4/n61 ,
         \add_98_4/n60 , \add_98_4/n59 , \add_98_4/n58 , \add_98_4/n57 ,
         \add_98_4/n56 , \add_98_4/n55 , \add_98_4/n54 , \add_98_4/n53 ,
         \add_98_4/n52 , \add_98_4/n51 , \add_98_4/n50 , \add_98_4/n49 ,
         \add_98_4/n48 , \add_98_4/n47 , \add_98_4/n46 , \add_98_4/n45 ,
         \add_98_4/n44 , \add_98_4/n43 , \add_98_4/n42 , \add_98_4/n41 ,
         \add_98_4/n40 , \add_98_4/n39 , \add_98_4/n38 , \add_98_4/n37 ,
         \add_98_4/n36 , \add_98_4/n35 , \add_98_4/n34 , \add_98_4/n33 ,
         \add_98_4/n32 , \add_98_4/n31 , \add_98_4/n30 , \add_98_4/n29 ,
         \add_98_4/n27 , \add_98_4/n26 , \add_98_4/n25 , \add_98_4/n24 ,
         \add_98_4/n23 , \add_98_4/n22 , \add_98_4/n21 , \add_98_4/n20 ,
         \add_98_4/n19 , \add_98_4/n18 , \add_98_4/n17 , \add_98_4/n16 ,
         \add_98_4/n15 , \add_98_4/n14 , \add_98_4/n13 , \add_98_4/n12 ,
         \add_98_4/n11 , \add_98_4/n10 , \add_98_4/n9 , \add_98_4/n8 ,
         \add_98_4/n7 , \add_98_4/n6 , \add_98_4/n5 , \add_98_4/n4 ,
         \add_98_4/n3 , \add_98_4/n2 , \add_98_4/n1 ;
  wire   [6:0] rnd_cnt_q;
  wire   [511:0] w_d;
  wire   [479:0] w_q;
  wire   [1:0] state;
  wire   [31:0] w;
  wire   [159:0] rnd_q;
  wire   [159:0] sha1_round_wire;
  wire   [159:0] rnd_d;
  wire   [159:0] cv_d;
  wire   [159:0] cv_q;
  wire   [159:0] cv_next_d;
  wire   [6:0] rnd_cnt_d;
  wire   [1:0] next_state;
  wire   [31:0] \sha1_round/f ;

  NAND2_X2 U3406 ( .A1(w[9]), .A2(n7159), .ZN(n4656) );
  NAND2_X2 U3407 ( .A1(w_q[9]), .A2(n7279), .ZN(n4655) );
  NAND2_X2 U3409 ( .A1(n4660), .A2(n4661), .ZN(w_d[99]) );
  NAND2_X2 U3410 ( .A1(w_q[67]), .A2(n7216), .ZN(n4661) );
  NAND2_X2 U3411 ( .A1(w_q[99]), .A2(n7279), .ZN(n4660) );
  NAND2_X2 U3412 ( .A1(n4663), .A2(n4664), .ZN(w_d[98]) );
  NAND2_X2 U3413 ( .A1(w_q[66]), .A2(n7216), .ZN(n4664) );
  NAND2_X2 U3414 ( .A1(w_q[98]), .A2(n7279), .ZN(n4663) );
  NAND2_X2 U3415 ( .A1(n4665), .A2(n4666), .ZN(w_d[97]) );
  NAND2_X2 U3416 ( .A1(w_q[65]), .A2(n7216), .ZN(n4666) );
  NAND2_X2 U3417 ( .A1(w_q[97]), .A2(n7279), .ZN(n4665) );
  NAND2_X2 U3418 ( .A1(n4667), .A2(n4668), .ZN(w_d[96]) );
  NAND2_X2 U3419 ( .A1(w_q[64]), .A2(n7216), .ZN(n4668) );
  NAND2_X2 U3420 ( .A1(w_q[96]), .A2(n7279), .ZN(n4667) );
  NAND2_X2 U3422 ( .A1(w[8]), .A2(n7159), .ZN(n4671) );
  NAND2_X2 U3423 ( .A1(w_q[8]), .A2(n7279), .ZN(n4670) );
  NAND2_X2 U3426 ( .A1(w[7]), .A2(n7159), .ZN(n4674) );
  NAND2_X2 U3427 ( .A1(w_q[7]), .A2(n7278), .ZN(n4673) );
  NAND2_X2 U3430 ( .A1(w[6]), .A2(n7159), .ZN(n4677) );
  NAND2_X2 U3431 ( .A1(w_q[6]), .A2(n7278), .ZN(n4676) );
  NAND2_X2 U3433 ( .A1(n4678), .A2(n4679), .ZN(w_d[63]) );
  NAND2_X2 U3434 ( .A1(w_q[31]), .A2(n7216), .ZN(n4679) );
  NAND2_X2 U3435 ( .A1(w_q[63]), .A2(n7278), .ZN(n4678) );
  NAND2_X2 U3436 ( .A1(n4680), .A2(n4681), .ZN(w_d[62]) );
  NAND2_X2 U3437 ( .A1(w_q[30]), .A2(n7216), .ZN(n4681) );
  NAND2_X2 U3438 ( .A1(w_q[62]), .A2(n7278), .ZN(n4680) );
  NAND2_X2 U3439 ( .A1(n4682), .A2(n4683), .ZN(w_d[61]) );
  NAND2_X2 U3440 ( .A1(w_q[29]), .A2(n7216), .ZN(n4683) );
  NAND2_X2 U3441 ( .A1(w_q[61]), .A2(n7278), .ZN(n4682) );
  NAND2_X2 U3442 ( .A1(n4684), .A2(n4685), .ZN(w_d[60]) );
  NAND2_X2 U3443 ( .A1(w_q[28]), .A2(n7215), .ZN(n4685) );
  NAND2_X2 U3444 ( .A1(w_q[60]), .A2(n7278), .ZN(n4684) );
  NAND2_X2 U3446 ( .A1(w[5]), .A2(n7159), .ZN(n4688) );
  NAND2_X2 U3447 ( .A1(w_q[5]), .A2(n7278), .ZN(n4687) );
  NAND2_X2 U3449 ( .A1(n4689), .A2(n4690), .ZN(w_d[59]) );
  NAND2_X2 U3450 ( .A1(w_q[27]), .A2(n7215), .ZN(n4690) );
  NAND2_X2 U3451 ( .A1(w_q[59]), .A2(n7278), .ZN(n4689) );
  NAND2_X2 U3452 ( .A1(n4691), .A2(n4692), .ZN(w_d[58]) );
  NAND2_X2 U3453 ( .A1(w_q[26]), .A2(n7215), .ZN(n4692) );
  NAND2_X2 U3454 ( .A1(w_q[58]), .A2(n7278), .ZN(n4691) );
  NAND2_X2 U3455 ( .A1(n4693), .A2(n4694), .ZN(w_d[57]) );
  NAND2_X2 U3456 ( .A1(w_q[25]), .A2(n7215), .ZN(n4694) );
  NAND2_X2 U3457 ( .A1(w_q[57]), .A2(n7278), .ZN(n4693) );
  NAND2_X2 U3458 ( .A1(n4695), .A2(n4696), .ZN(w_d[56]) );
  NAND2_X2 U3459 ( .A1(w_q[24]), .A2(n7215), .ZN(n4696) );
  NAND2_X2 U3460 ( .A1(w_q[56]), .A2(n7278), .ZN(n4695) );
  NAND2_X2 U3461 ( .A1(n4697), .A2(n4698), .ZN(w_d[55]) );
  NAND2_X2 U3462 ( .A1(w_q[23]), .A2(n7215), .ZN(n4698) );
  NAND2_X2 U3463 ( .A1(w_q[55]), .A2(n7277), .ZN(n4697) );
  NAND2_X2 U3464 ( .A1(n4699), .A2(n4700), .ZN(w_d[54]) );
  NAND2_X2 U3465 ( .A1(w_q[22]), .A2(n7215), .ZN(n4700) );
  NAND2_X2 U3466 ( .A1(w_q[54]), .A2(n7277), .ZN(n4699) );
  NAND2_X2 U3467 ( .A1(n4701), .A2(n4702), .ZN(w_d[53]) );
  NAND2_X2 U3468 ( .A1(w_q[21]), .A2(n7215), .ZN(n4702) );
  NAND2_X2 U3469 ( .A1(w_q[53]), .A2(n7277), .ZN(n4701) );
  NAND2_X2 U3470 ( .A1(n4703), .A2(n4704), .ZN(w_d[52]) );
  NAND2_X2 U3471 ( .A1(w_q[20]), .A2(n7215), .ZN(n4704) );
  NAND2_X2 U3472 ( .A1(w_q[52]), .A2(n7277), .ZN(n4703) );
  NAND2_X2 U3473 ( .A1(n4705), .A2(n4706), .ZN(w_d[51]) );
  NAND2_X2 U3474 ( .A1(w_q[19]), .A2(n7215), .ZN(n4706) );
  NAND2_X2 U3475 ( .A1(w_q[51]), .A2(n7277), .ZN(n4705) );
  NAND2_X2 U3476 ( .A1(n4707), .A2(n4708), .ZN(w_d[511]) );
  NAND2_X2 U3477 ( .A1(n7179), .A2(n4709), .ZN(n4708) );
  XOR2_X2 U3478 ( .A(n4710), .B(n4711), .Z(n4709) );
  XOR2_X2 U3479 ( .A(w_d[254]), .B(n4712), .Z(n4711) );
  XOR2_X2 U3480 ( .A(w_d[94]), .B(w_d[446]), .Z(n4710) );
  NAND2_X2 U3481 ( .A1(n4713), .A2(n4714), .ZN(w_d[94]) );
  NAND2_X2 U3482 ( .A1(w_q[62]), .A2(n7215), .ZN(n4714) );
  NAND2_X2 U3483 ( .A1(w_q[94]), .A2(n7277), .ZN(n4713) );
  NAND2_X2 U3484 ( .A1(n4715), .A2(n7181), .ZN(n4707) );
  NAND2_X2 U3485 ( .A1(n4717), .A2(n4718), .ZN(w_d[510]) );
  NAND2_X2 U3486 ( .A1(n7179), .A2(n4719), .ZN(n4718) );
  XOR2_X2 U3487 ( .A(n4720), .B(n4721), .Z(n4719) );
  XOR2_X2 U3488 ( .A(w_d[253]), .B(n4722), .Z(n4721) );
  XOR2_X2 U3489 ( .A(w_d[93]), .B(w_d[445]), .Z(n4720) );
  NAND2_X2 U3490 ( .A1(n4723), .A2(n4724), .ZN(w_d[93]) );
  NAND2_X2 U3491 ( .A1(w_q[61]), .A2(n7220), .ZN(n4724) );
  NAND2_X2 U3492 ( .A1(w_q[93]), .A2(n7277), .ZN(n4723) );
  NAND2_X2 U3493 ( .A1(n4712), .A2(n7181), .ZN(n4717) );
  NAND2_X2 U3494 ( .A1(n4725), .A2(n4726), .ZN(n4712) );
  NAND2_X2 U3495 ( .A1(w_q[478]), .A2(n7225), .ZN(n4726) );
  NAND2_X2 U3496 ( .A1(w[30]), .A2(n7277), .ZN(n4725) );
  NAND2_X2 U3497 ( .A1(n4727), .A2(n4728), .ZN(w_d[50]) );
  NAND2_X2 U3498 ( .A1(w_q[18]), .A2(n7196), .ZN(n4728) );
  NAND2_X2 U3499 ( .A1(w_q[50]), .A2(n7277), .ZN(n4727) );
  NAND2_X2 U3500 ( .A1(n4729), .A2(n4730), .ZN(w_d[509]) );
  NAND2_X2 U3501 ( .A1(n7179), .A2(n4731), .ZN(n4730) );
  XOR2_X2 U3502 ( .A(n4732), .B(n4733), .Z(n4731) );
  XOR2_X2 U3503 ( .A(w_d[252]), .B(n4734), .Z(n4733) );
  XOR2_X2 U3504 ( .A(w_d[92]), .B(w_d[444]), .Z(n4732) );
  NAND2_X2 U3505 ( .A1(n4735), .A2(n4736), .ZN(w_d[92]) );
  NAND2_X2 U3506 ( .A1(w_q[60]), .A2(n7219), .ZN(n4736) );
  NAND2_X2 U3507 ( .A1(w_q[92]), .A2(n7277), .ZN(n4735) );
  NAND2_X2 U3508 ( .A1(n4722), .A2(n7181), .ZN(n4729) );
  NAND2_X2 U3509 ( .A1(n4737), .A2(n4738), .ZN(n4722) );
  NAND2_X2 U3510 ( .A1(w_q[477]), .A2(n7224), .ZN(n4738) );
  NAND2_X2 U3511 ( .A1(w[29]), .A2(n7277), .ZN(n4737) );
  NAND2_X2 U3512 ( .A1(n4739), .A2(n4740), .ZN(w_d[508]) );
  NAND2_X2 U3513 ( .A1(n7179), .A2(n4741), .ZN(n4740) );
  XOR2_X2 U3514 ( .A(n4742), .B(n4743), .Z(n4741) );
  XOR2_X2 U3515 ( .A(w_d[251]), .B(n4744), .Z(n4743) );
  XOR2_X2 U3516 ( .A(w_d[91]), .B(w_d[443]), .Z(n4742) );
  NAND2_X2 U3517 ( .A1(n4745), .A2(n4746), .ZN(w_d[91]) );
  NAND2_X2 U3518 ( .A1(w_q[59]), .A2(n7226), .ZN(n4746) );
  NAND2_X2 U3519 ( .A1(w_q[91]), .A2(n7236), .ZN(n4745) );
  NAND2_X2 U3520 ( .A1(n4734), .A2(n7181), .ZN(n4739) );
  NAND2_X2 U3521 ( .A1(n4747), .A2(n4748), .ZN(n4734) );
  NAND2_X2 U3522 ( .A1(w_q[476]), .A2(n7223), .ZN(n4748) );
  NAND2_X2 U3523 ( .A1(w[28]), .A2(n7231), .ZN(n4747) );
  NAND2_X2 U3524 ( .A1(n4749), .A2(n4750), .ZN(w_d[507]) );
  NAND2_X2 U3525 ( .A1(n7179), .A2(n4751), .ZN(n4750) );
  XOR2_X2 U3526 ( .A(n4752), .B(n4753), .Z(n4751) );
  XOR2_X2 U3527 ( .A(w_d[250]), .B(n4754), .Z(n4753) );
  XOR2_X2 U3528 ( .A(w_d[90]), .B(w_d[442]), .Z(n4752) );
  NAND2_X2 U3529 ( .A1(n4755), .A2(n4756), .ZN(w_d[90]) );
  NAND2_X2 U3530 ( .A1(w_q[58]), .A2(n7220), .ZN(n4756) );
  NAND2_X2 U3531 ( .A1(w_q[90]), .A2(n7232), .ZN(n4755) );
  NAND2_X2 U3532 ( .A1(n4744), .A2(n7181), .ZN(n4749) );
  NAND2_X2 U3533 ( .A1(n4757), .A2(n4758), .ZN(n4744) );
  NAND2_X2 U3534 ( .A1(w_q[475]), .A2(n7222), .ZN(n4758) );
  NAND2_X2 U3535 ( .A1(w[27]), .A2(n7233), .ZN(n4757) );
  NAND2_X2 U3536 ( .A1(n4759), .A2(n4760), .ZN(w_d[506]) );
  NAND2_X2 U3537 ( .A1(n7179), .A2(n4761), .ZN(n4760) );
  XOR2_X2 U3538 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR2_X2 U3539 ( .A(w_d[249]), .B(n4764), .Z(n4763) );
  XOR2_X2 U3540 ( .A(w_d[89]), .B(w_d[441]), .Z(n4762) );
  NAND2_X2 U3541 ( .A1(n4765), .A2(n4766), .ZN(w_d[89]) );
  NAND2_X2 U3542 ( .A1(w_q[57]), .A2(n7219), .ZN(n4766) );
  NAND2_X2 U3543 ( .A1(w_q[89]), .A2(n7236), .ZN(n4765) );
  NAND2_X2 U3544 ( .A1(n4754), .A2(n7181), .ZN(n4759) );
  NAND2_X2 U3545 ( .A1(n4767), .A2(n4768), .ZN(n4754) );
  NAND2_X2 U3546 ( .A1(w_q[474]), .A2(n7221), .ZN(n4768) );
  NAND2_X2 U3547 ( .A1(w[26]), .A2(n7234), .ZN(n4767) );
  NAND2_X2 U3548 ( .A1(n4769), .A2(n4770), .ZN(w_d[505]) );
  NAND2_X2 U3549 ( .A1(n7179), .A2(n4771), .ZN(n4770) );
  XOR2_X2 U3550 ( .A(n4772), .B(n4773), .Z(n4771) );
  XOR2_X2 U3551 ( .A(w_d[248]), .B(n4774), .Z(n4773) );
  XOR2_X2 U3552 ( .A(w_d[88]), .B(w_d[440]), .Z(n4772) );
  NAND2_X2 U3553 ( .A1(n4775), .A2(n4776), .ZN(w_d[88]) );
  NAND2_X2 U3554 ( .A1(w_q[56]), .A2(n7219), .ZN(n4776) );
  NAND2_X2 U3555 ( .A1(w_q[88]), .A2(n7235), .ZN(n4775) );
  NAND2_X2 U3556 ( .A1(n4764), .A2(n7181), .ZN(n4769) );
  NAND2_X2 U3557 ( .A1(n4777), .A2(n4778), .ZN(n4764) );
  NAND2_X2 U3558 ( .A1(w_q[473]), .A2(n7225), .ZN(n4778) );
  NAND2_X2 U3559 ( .A1(w[25]), .A2(n7238), .ZN(n4777) );
  NAND2_X2 U3560 ( .A1(n4779), .A2(n4780), .ZN(w_d[504]) );
  NAND2_X2 U3561 ( .A1(n7179), .A2(n4781), .ZN(n4780) );
  XOR2_X2 U3562 ( .A(n4782), .B(n4783), .Z(n4781) );
  XOR2_X2 U3563 ( .A(w_d[247]), .B(n4784), .Z(n4783) );
  XOR2_X2 U3564 ( .A(w_d[87]), .B(w_d[439]), .Z(n4782) );
  NAND2_X2 U3565 ( .A1(n4785), .A2(n4786), .ZN(w_d[87]) );
  NAND2_X2 U3566 ( .A1(w_q[55]), .A2(n7226), .ZN(n4786) );
  NAND2_X2 U3567 ( .A1(w_q[87]), .A2(n7238), .ZN(n4785) );
  NAND2_X2 U3568 ( .A1(n4774), .A2(n7181), .ZN(n4779) );
  NAND2_X2 U3569 ( .A1(n4787), .A2(n4788), .ZN(n4774) );
  NAND2_X2 U3570 ( .A1(w_q[472]), .A2(n7224), .ZN(n4788) );
  NAND2_X2 U3571 ( .A1(w[24]), .A2(n7230), .ZN(n4787) );
  NAND2_X2 U3572 ( .A1(n4789), .A2(n4790), .ZN(w_d[503]) );
  NAND2_X2 U3573 ( .A1(n7179), .A2(n4791), .ZN(n4790) );
  XOR2_X2 U3574 ( .A(n4792), .B(n4793), .Z(n4791) );
  XOR2_X2 U3575 ( .A(w_d[246]), .B(n4794), .Z(n4793) );
  XOR2_X2 U3576 ( .A(w_d[86]), .B(w_d[438]), .Z(n4792) );
  NAND2_X2 U3577 ( .A1(n4795), .A2(n4796), .ZN(w_d[86]) );
  NAND2_X2 U3578 ( .A1(w_q[54]), .A2(n7219), .ZN(n4796) );
  NAND2_X2 U3579 ( .A1(w_q[86]), .A2(n7236), .ZN(n4795) );
  NAND2_X2 U3580 ( .A1(n4784), .A2(n7181), .ZN(n4789) );
  NAND2_X2 U3581 ( .A1(n4797), .A2(n4798), .ZN(n4784) );
  NAND2_X2 U3582 ( .A1(w_q[471]), .A2(n7223), .ZN(n4798) );
  NAND2_X2 U3583 ( .A1(w[23]), .A2(n7276), .ZN(n4797) );
  NAND2_X2 U3584 ( .A1(n4799), .A2(n4800), .ZN(w_d[502]) );
  NAND2_X2 U3585 ( .A1(n7179), .A2(n4801), .ZN(n4800) );
  XOR2_X2 U3586 ( .A(n4802), .B(n4803), .Z(n4801) );
  XOR2_X2 U3587 ( .A(w_d[245]), .B(n4804), .Z(n4803) );
  XOR2_X2 U3588 ( .A(w_d[85]), .B(w_d[437]), .Z(n4802) );
  NAND2_X2 U3589 ( .A1(n4805), .A2(n4806), .ZN(w_d[85]) );
  NAND2_X2 U3590 ( .A1(w_q[53]), .A2(n7220), .ZN(n4806) );
  NAND2_X2 U3591 ( .A1(w_q[85]), .A2(n7276), .ZN(n4805) );
  NAND2_X2 U3592 ( .A1(n4794), .A2(n7181), .ZN(n4799) );
  NAND2_X2 U3593 ( .A1(n4807), .A2(n4808), .ZN(n4794) );
  NAND2_X2 U3594 ( .A1(w_q[470]), .A2(n7222), .ZN(n4808) );
  NAND2_X2 U3595 ( .A1(w[22]), .A2(n7276), .ZN(n4807) );
  NAND2_X2 U3596 ( .A1(n4809), .A2(n4810), .ZN(w_d[501]) );
  NAND2_X2 U3597 ( .A1(n7178), .A2(n4811), .ZN(n4810) );
  XOR2_X2 U3598 ( .A(n4812), .B(n4813), .Z(n4811) );
  XOR2_X2 U3599 ( .A(w_d[244]), .B(n4814), .Z(n4813) );
  XOR2_X2 U3600 ( .A(w_d[84]), .B(w_d[436]), .Z(n4812) );
  NAND2_X2 U3601 ( .A1(n4815), .A2(n4816), .ZN(w_d[84]) );
  NAND2_X2 U3602 ( .A1(w_q[52]), .A2(n7226), .ZN(n4816) );
  NAND2_X2 U3603 ( .A1(w_q[84]), .A2(n7276), .ZN(n4815) );
  NAND2_X2 U3604 ( .A1(n4804), .A2(n7181), .ZN(n4809) );
  NAND2_X2 U3605 ( .A1(n4817), .A2(n4818), .ZN(n4804) );
  NAND2_X2 U3606 ( .A1(w_q[469]), .A2(n7221), .ZN(n4818) );
  NAND2_X2 U3607 ( .A1(w[21]), .A2(n7276), .ZN(n4817) );
  NAND2_X2 U3608 ( .A1(n4819), .A2(n4820), .ZN(w_d[500]) );
  NAND2_X2 U3609 ( .A1(n7178), .A2(n4821), .ZN(n4820) );
  XOR2_X2 U3610 ( .A(n4822), .B(n4823), .Z(n4821) );
  XOR2_X2 U3611 ( .A(w_d[243]), .B(n4824), .Z(n4823) );
  XOR2_X2 U3612 ( .A(w_d[83]), .B(w_d[435]), .Z(n4822) );
  NAND2_X2 U3613 ( .A1(n4825), .A2(n4826), .ZN(w_d[83]) );
  NAND2_X2 U3614 ( .A1(w_q[51]), .A2(n7220), .ZN(n4826) );
  NAND2_X2 U3615 ( .A1(w_q[83]), .A2(n7276), .ZN(n4825) );
  NAND2_X2 U3616 ( .A1(n4814), .A2(n7180), .ZN(n4819) );
  NAND2_X2 U3617 ( .A1(n4827), .A2(n4828), .ZN(n4814) );
  NAND2_X2 U3618 ( .A1(w_q[468]), .A2(n7225), .ZN(n4828) );
  NAND2_X2 U3619 ( .A1(w[20]), .A2(n7276), .ZN(n4827) );
  NAND2_X2 U3621 ( .A1(w[4]), .A2(n7159), .ZN(n4831) );
  NAND2_X2 U3622 ( .A1(w_q[4]), .A2(n7276), .ZN(n4830) );
  NAND2_X2 U3624 ( .A1(n4832), .A2(n4833), .ZN(w_d[49]) );
  NAND2_X2 U3625 ( .A1(w_q[17]), .A2(n7197), .ZN(n4833) );
  NAND2_X2 U3626 ( .A1(w_q[49]), .A2(n7276), .ZN(n4832) );
  NAND2_X2 U3627 ( .A1(n4834), .A2(n4835), .ZN(w_d[499]) );
  NAND2_X2 U3628 ( .A1(n7178), .A2(n4836), .ZN(n4835) );
  XOR2_X2 U3629 ( .A(n4837), .B(n4838), .Z(n4836) );
  XOR2_X2 U3630 ( .A(w_d[242]), .B(n4839), .Z(n4838) );
  XOR2_X2 U3631 ( .A(w_d[82]), .B(w_d[434]), .Z(n4837) );
  NAND2_X2 U3632 ( .A1(n4840), .A2(n4841), .ZN(w_d[82]) );
  NAND2_X2 U3633 ( .A1(w_q[50]), .A2(n7226), .ZN(n4841) );
  NAND2_X2 U3634 ( .A1(w_q[82]), .A2(n7276), .ZN(n4840) );
  NAND2_X2 U3635 ( .A1(n4824), .A2(n7180), .ZN(n4834) );
  NAND2_X2 U3636 ( .A1(n4842), .A2(n4843), .ZN(n4824) );
  NAND2_X2 U3637 ( .A1(w_q[467]), .A2(n7224), .ZN(n4843) );
  NAND2_X2 U3638 ( .A1(w[19]), .A2(n7276), .ZN(n4842) );
  NAND2_X2 U3639 ( .A1(n4844), .A2(n4845), .ZN(w_d[498]) );
  NAND2_X2 U3640 ( .A1(n7178), .A2(n4846), .ZN(n4845) );
  XOR2_X2 U3641 ( .A(n4847), .B(n4848), .Z(n4846) );
  XOR2_X2 U3642 ( .A(w_d[241]), .B(n4849), .Z(n4848) );
  XOR2_X2 U3643 ( .A(w_d[81]), .B(w_d[433]), .Z(n4847) );
  NAND2_X2 U3644 ( .A1(n4850), .A2(n4851), .ZN(w_d[81]) );
  NAND2_X2 U3645 ( .A1(w_q[49]), .A2(n7220), .ZN(n4851) );
  NAND2_X2 U3646 ( .A1(w_q[81]), .A2(n7235), .ZN(n4850) );
  NAND2_X2 U3647 ( .A1(n4839), .A2(n7180), .ZN(n4844) );
  NAND2_X2 U3648 ( .A1(n4852), .A2(n4853), .ZN(n4839) );
  NAND2_X2 U3649 ( .A1(w_q[466]), .A2(n7221), .ZN(n4853) );
  NAND2_X2 U3650 ( .A1(w[18]), .A2(n7230), .ZN(n4852) );
  NAND2_X2 U3651 ( .A1(n4854), .A2(n4855), .ZN(w_d[497]) );
  NAND2_X2 U3652 ( .A1(n7178), .A2(n4856), .ZN(n4855) );
  XOR2_X2 U3653 ( .A(n4857), .B(n4858), .Z(n4856) );
  XOR2_X2 U3654 ( .A(w_d[240]), .B(n4859), .Z(n4858) );
  XOR2_X2 U3655 ( .A(w_d[80]), .B(w_d[432]), .Z(n4857) );
  NAND2_X2 U3656 ( .A1(n4860), .A2(n4861), .ZN(w_d[80]) );
  NAND2_X2 U3657 ( .A1(w_q[48]), .A2(n7219), .ZN(n4861) );
  NAND2_X2 U3658 ( .A1(w_q[80]), .A2(n7236), .ZN(n4860) );
  NAND2_X2 U3659 ( .A1(n4849), .A2(n7180), .ZN(n4854) );
  NAND2_X2 U3660 ( .A1(n4862), .A2(n4863), .ZN(n4849) );
  NAND2_X2 U3661 ( .A1(w_q[465]), .A2(n7223), .ZN(n4863) );
  NAND2_X2 U3662 ( .A1(w[17]), .A2(n7233), .ZN(n4862) );
  NAND2_X2 U3663 ( .A1(n4864), .A2(n4865), .ZN(w_d[496]) );
  NAND2_X2 U3664 ( .A1(n7178), .A2(n4866), .ZN(n4865) );
  XOR2_X2 U3665 ( .A(n4867), .B(n4868), .Z(n4866) );
  XOR2_X2 U3666 ( .A(w_d[239]), .B(n4869), .Z(n4868) );
  XOR2_X2 U3667 ( .A(w_d[79]), .B(w_d[431]), .Z(n4867) );
  NAND2_X2 U3668 ( .A1(n4870), .A2(n4871), .ZN(w_d[79]) );
  NAND2_X2 U3669 ( .A1(w_q[47]), .A2(n7226), .ZN(n4871) );
  NAND2_X2 U3670 ( .A1(w_q[79]), .A2(n7231), .ZN(n4870) );
  NAND2_X2 U3671 ( .A1(n4859), .A2(n7180), .ZN(n4864) );
  NAND2_X2 U3672 ( .A1(n4872), .A2(n4873), .ZN(n4859) );
  NAND2_X2 U3673 ( .A1(w_q[464]), .A2(n7222), .ZN(n4873) );
  NAND2_X2 U3674 ( .A1(w[16]), .A2(n7234), .ZN(n4872) );
  NAND2_X2 U3675 ( .A1(n4874), .A2(n4875), .ZN(w_d[495]) );
  NAND2_X2 U3676 ( .A1(n7178), .A2(n4876), .ZN(n4875) );
  XOR2_X2 U3677 ( .A(n4877), .B(n4878), .Z(n4876) );
  XOR2_X2 U3678 ( .A(w_d[238]), .B(n4879), .Z(n4878) );
  XOR2_X2 U3679 ( .A(w_d[78]), .B(w_d[430]), .Z(n4877) );
  NAND2_X2 U3680 ( .A1(n4880), .A2(n4881), .ZN(w_d[78]) );
  NAND2_X2 U3681 ( .A1(w_q[46]), .A2(n7220), .ZN(n4881) );
  NAND2_X2 U3682 ( .A1(w_q[78]), .A2(n7235), .ZN(n4880) );
  NAND2_X2 U3683 ( .A1(n4869), .A2(n7180), .ZN(n4874) );
  NAND2_X2 U3684 ( .A1(n4882), .A2(n4883), .ZN(n4869) );
  NAND2_X2 U3685 ( .A1(w_q[463]), .A2(n7224), .ZN(n4883) );
  NAND2_X2 U3686 ( .A1(w[15]), .A2(n7234), .ZN(n4882) );
  NAND2_X2 U3687 ( .A1(n4884), .A2(n4885), .ZN(w_d[494]) );
  NAND2_X2 U3688 ( .A1(n7178), .A2(n4886), .ZN(n4885) );
  XOR2_X2 U3689 ( .A(n4887), .B(n4888), .Z(n4886) );
  XOR2_X2 U3690 ( .A(w_d[237]), .B(n4889), .Z(n4888) );
  XOR2_X2 U3691 ( .A(w_d[77]), .B(w_d[429]), .Z(n4887) );
  NAND2_X2 U3692 ( .A1(n4890), .A2(n4891), .ZN(w_d[77]) );
  NAND2_X2 U3693 ( .A1(w_q[45]), .A2(n7221), .ZN(n4891) );
  NAND2_X2 U3694 ( .A1(w_q[77]), .A2(n7236), .ZN(n4890) );
  NAND2_X2 U3695 ( .A1(n4879), .A2(n7180), .ZN(n4884) );
  NAND2_X2 U3696 ( .A1(n4892), .A2(n4893), .ZN(n4879) );
  NAND2_X2 U3697 ( .A1(w_q[462]), .A2(n7223), .ZN(n4893) );
  NAND2_X2 U3698 ( .A1(w[14]), .A2(n7232), .ZN(n4892) );
  NAND2_X2 U3699 ( .A1(n4894), .A2(n4895), .ZN(w_d[493]) );
  NAND2_X2 U3700 ( .A1(n7178), .A2(n4896), .ZN(n4895) );
  XOR2_X2 U3701 ( .A(n4897), .B(n4898), .Z(n4896) );
  XOR2_X2 U3702 ( .A(w_d[236]), .B(n4899), .Z(n4898) );
  XOR2_X2 U3703 ( .A(w_d[76]), .B(w_d[428]), .Z(n4897) );
  NAND2_X2 U3704 ( .A1(n4900), .A2(n4901), .ZN(w_d[76]) );
  NAND2_X2 U3705 ( .A1(w_q[44]), .A2(n7223), .ZN(n4901) );
  NAND2_X2 U3706 ( .A1(w_q[76]), .A2(n7238), .ZN(n4900) );
  NAND2_X2 U3707 ( .A1(n4889), .A2(n7180), .ZN(n4894) );
  NAND2_X2 U3708 ( .A1(n4902), .A2(n4903), .ZN(n4889) );
  NAND2_X2 U3709 ( .A1(w_q[461]), .A2(n7222), .ZN(n4903) );
  NAND2_X2 U3710 ( .A1(w[13]), .A2(n7235), .ZN(n4902) );
  NAND2_X2 U3711 ( .A1(n4904), .A2(n4905), .ZN(w_d[492]) );
  NAND2_X2 U3712 ( .A1(n7178), .A2(n4906), .ZN(n4905) );
  XOR2_X2 U3713 ( .A(n4907), .B(n4908), .Z(n4906) );
  XOR2_X2 U3714 ( .A(w_d[235]), .B(n4909), .Z(n4908) );
  XOR2_X2 U3715 ( .A(w_d[75]), .B(w_d[427]), .Z(n4907) );
  NAND2_X2 U3716 ( .A1(n4910), .A2(n4911), .ZN(w_d[75]) );
  NAND2_X2 U3717 ( .A1(w_q[43]), .A2(n7222), .ZN(n4911) );
  NAND2_X2 U3718 ( .A1(w_q[75]), .A2(n7231), .ZN(n4910) );
  NAND2_X2 U3719 ( .A1(n4899), .A2(n7180), .ZN(n4904) );
  NAND2_X2 U3720 ( .A1(n4912), .A2(n4913), .ZN(n4899) );
  NAND2_X2 U3721 ( .A1(w_q[460]), .A2(n7225), .ZN(n4913) );
  NAND2_X2 U3722 ( .A1(w[12]), .A2(n7230), .ZN(n4912) );
  NAND2_X2 U3723 ( .A1(n4914), .A2(n4915), .ZN(w_d[491]) );
  NAND2_X2 U3724 ( .A1(n7178), .A2(n4916), .ZN(n4915) );
  XOR2_X2 U3725 ( .A(n4917), .B(n4918), .Z(n4916) );
  XOR2_X2 U3726 ( .A(w_d[234]), .B(n4919), .Z(n4918) );
  XOR2_X2 U3727 ( .A(w_d[74]), .B(w_d[426]), .Z(n4917) );
  NAND2_X2 U3728 ( .A1(n4920), .A2(n4921), .ZN(w_d[74]) );
  NAND2_X2 U3729 ( .A1(w_q[42]), .A2(n7225), .ZN(n4921) );
  NAND2_X2 U3730 ( .A1(w_q[74]), .A2(n7232), .ZN(n4920) );
  NAND2_X2 U3731 ( .A1(n4909), .A2(n7180), .ZN(n4914) );
  NAND2_X2 U3732 ( .A1(n4922), .A2(n4923), .ZN(n4909) );
  NAND2_X2 U3733 ( .A1(w_q[459]), .A2(n7221), .ZN(n4923) );
  NAND2_X2 U3735 ( .A1(n4924), .A2(n4925), .ZN(w_d[490]) );
  NAND2_X2 U3736 ( .A1(n7177), .A2(n4926), .ZN(n4925) );
  XOR2_X2 U3737 ( .A(n4927), .B(n4928), .Z(n4926) );
  XOR2_X2 U3738 ( .A(w_d[233]), .B(n4929), .Z(n4928) );
  XOR2_X2 U3739 ( .A(w_d[73]), .B(w_d[425]), .Z(n4927) );
  NAND2_X2 U3740 ( .A1(n4930), .A2(n4931), .ZN(w_d[73]) );
  NAND2_X2 U3741 ( .A1(w_q[41]), .A2(n7219), .ZN(n4931) );
  NAND2_X2 U3742 ( .A1(w_q[73]), .A2(n7235), .ZN(n4930) );
  NAND2_X2 U3743 ( .A1(n4919), .A2(n7180), .ZN(n4924) );
  NAND2_X2 U3744 ( .A1(n4932), .A2(n4933), .ZN(n4919) );
  NAND2_X2 U3745 ( .A1(w_q[458]), .A2(n7224), .ZN(n4933) );
  NAND2_X2 U3746 ( .A1(w[10]), .A2(n7234), .ZN(n4932) );
  NAND2_X2 U3747 ( .A1(n4934), .A2(n4935), .ZN(w_d[48]) );
  NAND2_X2 U3748 ( .A1(w_q[16]), .A2(n7212), .ZN(n4935) );
  NAND2_X2 U3749 ( .A1(w_q[48]), .A2(n7273), .ZN(n4934) );
  NAND2_X2 U3750 ( .A1(n4936), .A2(n4937), .ZN(w_d[489]) );
  NAND2_X2 U3751 ( .A1(n7177), .A2(n4938), .ZN(n4937) );
  XOR2_X2 U3752 ( .A(n4939), .B(n4940), .Z(n4938) );
  XOR2_X2 U3753 ( .A(w_d[232]), .B(n4941), .Z(n4940) );
  XOR2_X2 U3754 ( .A(w_d[72]), .B(w_d[424]), .Z(n4939) );
  NAND2_X2 U3755 ( .A1(n4942), .A2(n4943), .ZN(w_d[72]) );
  NAND2_X2 U3756 ( .A1(w_q[40]), .A2(n7226), .ZN(n4943) );
  NAND2_X2 U3757 ( .A1(w_q[72]), .A2(n7236), .ZN(n4942) );
  NAND2_X2 U3758 ( .A1(n4929), .A2(n7180), .ZN(n4936) );
  NAND2_X2 U3759 ( .A1(n4944), .A2(n4945), .ZN(n4929) );
  NAND2_X2 U3760 ( .A1(w_q[457]), .A2(n7221), .ZN(n4945) );
  NAND2_X2 U3761 ( .A1(w[9]), .A2(n7233), .ZN(n4944) );
  NAND2_X2 U3762 ( .A1(n4946), .A2(n4947), .ZN(w_d[488]) );
  NAND2_X2 U3763 ( .A1(n7177), .A2(n4948), .ZN(n4947) );
  XOR2_X2 U3764 ( .A(n4949), .B(n4950), .Z(n4948) );
  XOR2_X2 U3765 ( .A(w_d[231]), .B(n4951), .Z(n4950) );
  XOR2_X2 U3766 ( .A(w_d[71]), .B(w_d[423]), .Z(n4949) );
  NAND2_X2 U3767 ( .A1(n4952), .A2(n4953), .ZN(w_d[71]) );
  NAND2_X2 U3768 ( .A1(w_q[39]), .A2(n7220), .ZN(n4953) );
  NAND2_X2 U3769 ( .A1(w_q[71]), .A2(n7231), .ZN(n4952) );
  NAND2_X2 U3770 ( .A1(n4941), .A2(n7180), .ZN(n4946) );
  NAND2_X2 U3771 ( .A1(n4954), .A2(n4955), .ZN(n4941) );
  NAND2_X2 U3772 ( .A1(w_q[456]), .A2(n7224), .ZN(n4955) );
  NAND2_X2 U3773 ( .A1(w[8]), .A2(n7230), .ZN(n4954) );
  NAND2_X2 U3774 ( .A1(n4956), .A2(n4957), .ZN(w_d[487]) );
  NAND2_X2 U3775 ( .A1(n7177), .A2(n4958), .ZN(n4957) );
  XOR2_X2 U3776 ( .A(n4959), .B(n4960), .Z(n4958) );
  XOR2_X2 U3777 ( .A(w_d[230]), .B(n4961), .Z(n4960) );
  XOR2_X2 U3778 ( .A(w_d[70]), .B(w_d[422]), .Z(n4959) );
  NAND2_X2 U3779 ( .A1(n4962), .A2(n4963), .ZN(w_d[70]) );
  NAND2_X2 U3780 ( .A1(w_q[38]), .A2(n7219), .ZN(n4963) );
  NAND2_X2 U3781 ( .A1(w_q[70]), .A2(n7236), .ZN(n4962) );
  NAND2_X2 U3782 ( .A1(n4951), .A2(n7180), .ZN(n4956) );
  NAND2_X2 U3783 ( .A1(n4964), .A2(n4965), .ZN(n4951) );
  NAND2_X2 U3784 ( .A1(w_q[455]), .A2(n7225), .ZN(n4965) );
  NAND2_X2 U3785 ( .A1(w[7]), .A2(n7233), .ZN(n4964) );
  NAND2_X2 U3786 ( .A1(n4966), .A2(n4967), .ZN(w_d[486]) );
  NAND2_X2 U3787 ( .A1(n7177), .A2(n4968), .ZN(n4967) );
  XOR2_X2 U3788 ( .A(n4969), .B(n4970), .Z(n4968) );
  XOR2_X2 U3789 ( .A(w_d[229]), .B(n4971), .Z(n4970) );
  XOR2_X2 U3790 ( .A(w_d[69]), .B(w_d[421]), .Z(n4969) );
  NAND2_X2 U3791 ( .A1(n4972), .A2(n4973), .ZN(w_d[69]) );
  NAND2_X2 U3792 ( .A1(w_q[37]), .A2(n7221), .ZN(n4973) );
  NAND2_X2 U3793 ( .A1(w_q[69]), .A2(n7238), .ZN(n4972) );
  NAND2_X2 U3794 ( .A1(n4961), .A2(n7180), .ZN(n4966) );
  NAND2_X2 U3795 ( .A1(n4974), .A2(n4975), .ZN(n4961) );
  NAND2_X2 U3796 ( .A1(w_q[454]), .A2(n7223), .ZN(n4975) );
  NAND2_X2 U3797 ( .A1(w[6]), .A2(n7234), .ZN(n4974) );
  NAND2_X2 U3798 ( .A1(n4976), .A2(n4977), .ZN(w_d[485]) );
  NAND2_X2 U3799 ( .A1(n7177), .A2(n4978), .ZN(n4977) );
  XOR2_X2 U3800 ( .A(n4979), .B(n4980), .Z(n4978) );
  XOR2_X2 U3801 ( .A(w_d[228]), .B(n4981), .Z(n4980) );
  XOR2_X2 U3802 ( .A(w_d[68]), .B(w_d[420]), .Z(n4979) );
  NAND2_X2 U3803 ( .A1(n4982), .A2(n4983), .ZN(w_d[68]) );
  NAND2_X2 U3804 ( .A1(w_q[36]), .A2(n7224), .ZN(n4983) );
  NAND2_X2 U3805 ( .A1(w_q[68]), .A2(n7230), .ZN(n4982) );
  NAND2_X2 U3806 ( .A1(n4971), .A2(n7180), .ZN(n4976) );
  NAND2_X2 U3807 ( .A1(n4984), .A2(n4985), .ZN(n4971) );
  NAND2_X2 U3808 ( .A1(w_q[453]), .A2(n7222), .ZN(n4985) );
  NAND2_X2 U3809 ( .A1(w[5]), .A2(n7232), .ZN(n4984) );
  NAND2_X2 U3810 ( .A1(n4986), .A2(n4987), .ZN(w_d[484]) );
  NAND2_X2 U3811 ( .A1(n7177), .A2(n4988), .ZN(n4987) );
  XOR2_X2 U3812 ( .A(n4989), .B(n4990), .Z(n4988) );
  XOR2_X2 U3813 ( .A(w_d[227]), .B(n4991), .Z(n4990) );
  XOR2_X2 U3814 ( .A(w_d[67]), .B(w_d[419]), .Z(n4989) );
  NAND2_X2 U3815 ( .A1(n4992), .A2(n4993), .ZN(w_d[67]) );
  NAND2_X2 U3816 ( .A1(w_q[35]), .A2(n7217), .ZN(n4993) );
  NAND2_X2 U3817 ( .A1(w_q[67]), .A2(n7232), .ZN(n4992) );
  NAND2_X2 U3818 ( .A1(n4981), .A2(n7180), .ZN(n4986) );
  NAND2_X2 U3819 ( .A1(n4994), .A2(n4995), .ZN(n4981) );
  NAND2_X2 U3820 ( .A1(w_q[452]), .A2(n7217), .ZN(n4995) );
  NAND2_X2 U3821 ( .A1(w[4]), .A2(n7233), .ZN(n4994) );
  NAND2_X2 U3822 ( .A1(n4996), .A2(n4997), .ZN(w_d[483]) );
  NAND2_X2 U3823 ( .A1(n7177), .A2(n4998), .ZN(n4997) );
  XOR2_X2 U3824 ( .A(n4999), .B(n5000), .Z(n4998) );
  XOR2_X2 U3825 ( .A(w_d[226]), .B(n5001), .Z(n5000) );
  XOR2_X2 U3826 ( .A(w_d[66]), .B(w_d[418]), .Z(n4999) );
  NAND2_X2 U3827 ( .A1(n5002), .A2(n5003), .ZN(w_d[66]) );
  NAND2_X2 U3828 ( .A1(w_q[34]), .A2(n7217), .ZN(n5003) );
  NAND2_X2 U3829 ( .A1(w_q[66]), .A2(n7235), .ZN(n5002) );
  NAND2_X2 U3830 ( .A1(n4991), .A2(n7180), .ZN(n4996) );
  NAND2_X2 U3831 ( .A1(n5004), .A2(n5005), .ZN(n4991) );
  NAND2_X2 U3832 ( .A1(w_q[451]), .A2(n7217), .ZN(n5005) );
  NAND2_X2 U3833 ( .A1(w[3]), .A2(n7231), .ZN(n5004) );
  NAND2_X2 U3834 ( .A1(n5006), .A2(n5007), .ZN(w_d[482]) );
  NAND2_X2 U3835 ( .A1(n7177), .A2(n5008), .ZN(n5007) );
  XOR2_X2 U3836 ( .A(n5009), .B(n5010), .Z(n5008) );
  XOR2_X2 U3837 ( .A(w_d[225]), .B(n5011), .Z(n5010) );
  XOR2_X2 U3838 ( .A(w_d[65]), .B(w_d[417]), .Z(n5009) );
  NAND2_X2 U3839 ( .A1(n5012), .A2(n5013), .ZN(w_d[65]) );
  NAND2_X2 U3840 ( .A1(w_q[33]), .A2(n7217), .ZN(n5013) );
  NAND2_X2 U3841 ( .A1(w_q[65]), .A2(n7275), .ZN(n5012) );
  NAND2_X2 U3842 ( .A1(n5001), .A2(n7180), .ZN(n5006) );
  NAND2_X2 U3843 ( .A1(n5014), .A2(n5015), .ZN(n5001) );
  NAND2_X2 U3844 ( .A1(w_q[450]), .A2(n7217), .ZN(n5015) );
  NAND2_X2 U3845 ( .A1(w[2]), .A2(n7275), .ZN(n5014) );
  NAND2_X2 U3846 ( .A1(n5016), .A2(n5017), .ZN(w_d[481]) );
  NAND2_X2 U3847 ( .A1(n7177), .A2(n5018), .ZN(n5017) );
  XOR2_X2 U3848 ( .A(n5019), .B(n5020), .Z(n5018) );
  XOR2_X2 U3849 ( .A(w_d[224]), .B(n5021), .Z(n5020) );
  XOR2_X2 U3850 ( .A(w_d[64]), .B(w_d[416]), .Z(n5019) );
  NAND2_X2 U3851 ( .A1(n5022), .A2(n5023), .ZN(w_d[64]) );
  NAND2_X2 U3852 ( .A1(w_q[32]), .A2(n7225), .ZN(n5023) );
  NAND2_X2 U3853 ( .A1(w_q[64]), .A2(n7275), .ZN(n5022) );
  NAND2_X2 U3854 ( .A1(n5011), .A2(n7180), .ZN(n5016) );
  NAND2_X2 U3855 ( .A1(n5024), .A2(n5025), .ZN(n5011) );
  NAND2_X2 U3856 ( .A1(w_q[449]), .A2(n7217), .ZN(n5025) );
  NAND2_X2 U3857 ( .A1(w[1]), .A2(n7275), .ZN(n5024) );
  NAND2_X2 U3858 ( .A1(n5026), .A2(n5027), .ZN(w_d[480]) );
  NAND2_X2 U3859 ( .A1(n5021), .A2(n7180), .ZN(n5027) );
  NAND2_X2 U3860 ( .A1(n5028), .A2(n5029), .ZN(n5021) );
  NAND2_X2 U3861 ( .A1(w_q[448]), .A2(n7217), .ZN(n5029) );
  NAND2_X2 U3862 ( .A1(w[0]), .A2(n7275), .ZN(n5028) );
  NAND2_X2 U3863 ( .A1(n7177), .A2(n5030), .ZN(n5026) );
  XOR2_X2 U3864 ( .A(n5031), .B(n5032), .Z(n5030) );
  XOR2_X2 U3865 ( .A(w_d[447]), .B(w_d[255]), .Z(n5032) );
  XOR2_X2 U3866 ( .A(w_d[95]), .B(n4715), .Z(n5031) );
  NAND2_X2 U3867 ( .A1(n5033), .A2(n5034), .ZN(n4715) );
  NAND2_X2 U3868 ( .A1(w_q[479]), .A2(n7223), .ZN(n5034) );
  NAND2_X2 U3869 ( .A1(w[31]), .A2(n7275), .ZN(n5033) );
  NAND2_X2 U3870 ( .A1(n5035), .A2(n5036), .ZN(w_d[95]) );
  NAND2_X2 U3871 ( .A1(w_q[63]), .A2(n7222), .ZN(n5036) );
  NAND2_X2 U3872 ( .A1(w_q[95]), .A2(n7275), .ZN(n5035) );
  NAND2_X2 U3875 ( .A1(n5039), .A2(n5040), .ZN(w_d[47]) );
  NAND2_X2 U3876 ( .A1(w_q[15]), .A2(n7214), .ZN(n5040) );
  NAND2_X2 U3877 ( .A1(w_q[47]), .A2(n7275), .ZN(n5039) );
  NAND2_X2 U3878 ( .A1(n5041), .A2(n5042), .ZN(w_d[479]) );
  NAND2_X2 U3879 ( .A1(w_q[447]), .A2(n7214), .ZN(n5042) );
  NAND2_X2 U3880 ( .A1(w_q[479]), .A2(n7275), .ZN(n5041) );
  NAND2_X2 U3881 ( .A1(n5043), .A2(n5044), .ZN(w_d[478]) );
  NAND2_X2 U3882 ( .A1(w_q[446]), .A2(n7214), .ZN(n5044) );
  NAND2_X2 U3883 ( .A1(w_q[478]), .A2(n7275), .ZN(n5043) );
  NAND2_X2 U3884 ( .A1(n5045), .A2(n5046), .ZN(w_d[477]) );
  NAND2_X2 U3885 ( .A1(w_q[445]), .A2(n7214), .ZN(n5046) );
  NAND2_X2 U3886 ( .A1(w_q[477]), .A2(n7275), .ZN(n5045) );
  NAND2_X2 U3887 ( .A1(n5047), .A2(n5048), .ZN(w_d[476]) );
  NAND2_X2 U3888 ( .A1(w_q[444]), .A2(n7214), .ZN(n5048) );
  NAND2_X2 U3889 ( .A1(w_q[476]), .A2(n7274), .ZN(n5047) );
  NAND2_X2 U3890 ( .A1(n5049), .A2(n5050), .ZN(w_d[475]) );
  NAND2_X2 U3891 ( .A1(w_q[443]), .A2(n7214), .ZN(n5050) );
  NAND2_X2 U3892 ( .A1(w_q[475]), .A2(n7274), .ZN(n5049) );
  NAND2_X2 U3893 ( .A1(n5051), .A2(n5052), .ZN(w_d[474]) );
  NAND2_X2 U3894 ( .A1(w_q[442]), .A2(n7214), .ZN(n5052) );
  NAND2_X2 U3895 ( .A1(w_q[474]), .A2(n7274), .ZN(n5051) );
  NAND2_X2 U3896 ( .A1(n5053), .A2(n5054), .ZN(w_d[473]) );
  NAND2_X2 U3897 ( .A1(w_q[441]), .A2(n7214), .ZN(n5054) );
  NAND2_X2 U3898 ( .A1(w_q[473]), .A2(n7274), .ZN(n5053) );
  NAND2_X2 U3899 ( .A1(n5055), .A2(n5056), .ZN(w_d[472]) );
  NAND2_X2 U3900 ( .A1(w_q[440]), .A2(n7214), .ZN(n5056) );
  NAND2_X2 U3901 ( .A1(w_q[472]), .A2(n7274), .ZN(n5055) );
  NAND2_X2 U3902 ( .A1(n5057), .A2(n5058), .ZN(w_d[471]) );
  NAND2_X2 U3903 ( .A1(w_q[439]), .A2(n7214), .ZN(n5058) );
  NAND2_X2 U3904 ( .A1(w_q[471]), .A2(n7274), .ZN(n5057) );
  NAND2_X2 U3905 ( .A1(n5059), .A2(n5060), .ZN(w_d[470]) );
  NAND2_X2 U3906 ( .A1(w_q[438]), .A2(n7214), .ZN(n5060) );
  NAND2_X2 U3907 ( .A1(w_q[470]), .A2(n7274), .ZN(n5059) );
  NAND2_X2 U3908 ( .A1(n5061), .A2(n5062), .ZN(w_d[46]) );
  NAND2_X2 U3909 ( .A1(w_q[14]), .A2(n7213), .ZN(n5062) );
  NAND2_X2 U3910 ( .A1(w_q[46]), .A2(n7274), .ZN(n5061) );
  NAND2_X2 U3911 ( .A1(n5063), .A2(n5064), .ZN(w_d[469]) );
  NAND2_X2 U3912 ( .A1(w_q[437]), .A2(n7213), .ZN(n5064) );
  NAND2_X2 U3913 ( .A1(w_q[469]), .A2(n7274), .ZN(n5063) );
  NAND2_X2 U3914 ( .A1(n5065), .A2(n5066), .ZN(w_d[468]) );
  NAND2_X2 U3915 ( .A1(w_q[436]), .A2(n7213), .ZN(n5066) );
  NAND2_X2 U3916 ( .A1(w_q[468]), .A2(n7274), .ZN(n5065) );
  NAND2_X2 U3917 ( .A1(n5067), .A2(n5068), .ZN(w_d[467]) );
  NAND2_X2 U3918 ( .A1(w_q[435]), .A2(n7213), .ZN(n5068) );
  NAND2_X2 U3919 ( .A1(w_q[467]), .A2(n7274), .ZN(n5067) );
  NAND2_X2 U3920 ( .A1(n5069), .A2(n5070), .ZN(w_d[466]) );
  NAND2_X2 U3921 ( .A1(w_q[434]), .A2(n7213), .ZN(n5070) );
  NAND2_X2 U3922 ( .A1(w_q[466]), .A2(n7273), .ZN(n5069) );
  NAND2_X2 U3923 ( .A1(n5071), .A2(n5072), .ZN(w_d[465]) );
  NAND2_X2 U3924 ( .A1(w_q[433]), .A2(n7213), .ZN(n5072) );
  NAND2_X2 U3925 ( .A1(w_q[465]), .A2(n7273), .ZN(n5071) );
  NAND2_X2 U3926 ( .A1(n5073), .A2(n5074), .ZN(w_d[464]) );
  NAND2_X2 U3927 ( .A1(w_q[432]), .A2(n7213), .ZN(n5074) );
  NAND2_X2 U3928 ( .A1(w_q[464]), .A2(n7273), .ZN(n5073) );
  NAND2_X2 U3929 ( .A1(n5075), .A2(n5076), .ZN(w_d[463]) );
  NAND2_X2 U3930 ( .A1(w_q[431]), .A2(n7213), .ZN(n5076) );
  NAND2_X2 U3931 ( .A1(w_q[463]), .A2(n7273), .ZN(n5075) );
  NAND2_X2 U3932 ( .A1(n5077), .A2(n5078), .ZN(w_d[462]) );
  NAND2_X2 U3933 ( .A1(w_q[430]), .A2(n7213), .ZN(n5078) );
  NAND2_X2 U3934 ( .A1(w_q[462]), .A2(n7273), .ZN(n5077) );
  NAND2_X2 U3935 ( .A1(n5079), .A2(n5080), .ZN(w_d[461]) );
  NAND2_X2 U3936 ( .A1(w_q[429]), .A2(n7213), .ZN(n5080) );
  NAND2_X2 U3937 ( .A1(w_q[461]), .A2(n7273), .ZN(n5079) );
  NAND2_X2 U3938 ( .A1(n5081), .A2(n5082), .ZN(w_d[460]) );
  NAND2_X2 U3939 ( .A1(w_q[428]), .A2(n7213), .ZN(n5082) );
  NAND2_X2 U3940 ( .A1(w_q[460]), .A2(n7273), .ZN(n5081) );
  NAND2_X2 U3941 ( .A1(n5083), .A2(n5084), .ZN(w_d[45]) );
  NAND2_X2 U3942 ( .A1(w_q[13]), .A2(n7212), .ZN(n5084) );
  NAND2_X2 U3943 ( .A1(w_q[45]), .A2(n7273), .ZN(n5083) );
  NAND2_X2 U3944 ( .A1(n5085), .A2(n5086), .ZN(w_d[459]) );
  NAND2_X2 U3945 ( .A1(w_q[427]), .A2(n7212), .ZN(n5086) );
  NAND2_X2 U3946 ( .A1(w_q[459]), .A2(n7273), .ZN(n5085) );
  NAND2_X2 U3947 ( .A1(n5087), .A2(n5088), .ZN(w_d[458]) );
  NAND2_X2 U3948 ( .A1(w_q[426]), .A2(n7212), .ZN(n5088) );
  NAND2_X2 U3949 ( .A1(w_q[458]), .A2(n7273), .ZN(n5087) );
  NAND2_X2 U3950 ( .A1(n5089), .A2(n5090), .ZN(w_d[457]) );
  NAND2_X2 U3951 ( .A1(w_q[425]), .A2(n7212), .ZN(n5090) );
  NAND2_X2 U3952 ( .A1(w_q[457]), .A2(n7273), .ZN(n5089) );
  NAND2_X2 U3953 ( .A1(n5091), .A2(n5092), .ZN(w_d[456]) );
  NAND2_X2 U3954 ( .A1(w_q[424]), .A2(n7212), .ZN(n5092) );
  NAND2_X2 U3955 ( .A1(w_q[456]), .A2(n7272), .ZN(n5091) );
  NAND2_X2 U3956 ( .A1(n5093), .A2(n5094), .ZN(w_d[455]) );
  NAND2_X2 U3957 ( .A1(w_q[423]), .A2(n7212), .ZN(n5094) );
  NAND2_X2 U3958 ( .A1(w_q[455]), .A2(n7272), .ZN(n5093) );
  NAND2_X2 U3959 ( .A1(n5095), .A2(n5096), .ZN(w_d[454]) );
  NAND2_X2 U3960 ( .A1(w_q[422]), .A2(n7212), .ZN(n5096) );
  NAND2_X2 U3961 ( .A1(w_q[454]), .A2(n7272), .ZN(n5095) );
  NAND2_X2 U3962 ( .A1(n5097), .A2(n5098), .ZN(w_d[453]) );
  NAND2_X2 U3963 ( .A1(w_q[421]), .A2(n7212), .ZN(n5098) );
  NAND2_X2 U3964 ( .A1(w_q[453]), .A2(n7272), .ZN(n5097) );
  NAND2_X2 U3965 ( .A1(n5099), .A2(n5100), .ZN(w_d[452]) );
  NAND2_X2 U3966 ( .A1(w_q[420]), .A2(n7212), .ZN(n5100) );
  NAND2_X2 U3967 ( .A1(w_q[452]), .A2(n7272), .ZN(n5099) );
  NAND2_X2 U3968 ( .A1(n5101), .A2(n5102), .ZN(w_d[451]) );
  NAND2_X2 U3969 ( .A1(w_q[419]), .A2(n7212), .ZN(n5102) );
  NAND2_X2 U3970 ( .A1(w_q[451]), .A2(n7272), .ZN(n5101) );
  NAND2_X2 U3971 ( .A1(n5103), .A2(n5104), .ZN(w_d[450]) );
  NAND2_X2 U3972 ( .A1(w_q[418]), .A2(n7212), .ZN(n5104) );
  NAND2_X2 U3973 ( .A1(w_q[450]), .A2(n7272), .ZN(n5103) );
  NAND2_X2 U3974 ( .A1(n5105), .A2(n5106), .ZN(w_d[44]) );
  NAND2_X2 U3975 ( .A1(w_q[12]), .A2(n7216), .ZN(n5106) );
  NAND2_X2 U3976 ( .A1(w_q[44]), .A2(n7272), .ZN(n5105) );
  NAND2_X2 U3977 ( .A1(n5107), .A2(n5108), .ZN(w_d[449]) );
  NAND2_X2 U3978 ( .A1(w_q[417]), .A2(n7196), .ZN(n5108) );
  NAND2_X2 U3979 ( .A1(w_q[449]), .A2(n7272), .ZN(n5107) );
  NAND2_X2 U3980 ( .A1(n5109), .A2(n5110), .ZN(w_d[448]) );
  NAND2_X2 U3981 ( .A1(w_q[416]), .A2(n7197), .ZN(n5110) );
  NAND2_X2 U3982 ( .A1(w_q[448]), .A2(n7272), .ZN(n5109) );
  NAND2_X2 U3983 ( .A1(n5111), .A2(n5112), .ZN(w_d[447]) );
  NAND2_X2 U3984 ( .A1(w_q[415]), .A2(n7218), .ZN(n5112) );
  NAND2_X2 U3985 ( .A1(w_q[447]), .A2(n7272), .ZN(n5111) );
  NAND2_X2 U3986 ( .A1(n5113), .A2(n5114), .ZN(w_d[446]) );
  NAND2_X2 U3987 ( .A1(w_q[414]), .A2(n7218), .ZN(n5114) );
  NAND2_X2 U3988 ( .A1(w_q[446]), .A2(n7271), .ZN(n5113) );
  NAND2_X2 U3989 ( .A1(n5115), .A2(n5116), .ZN(w_d[445]) );
  NAND2_X2 U3990 ( .A1(w_q[413]), .A2(n7218), .ZN(n5116) );
  NAND2_X2 U3991 ( .A1(w_q[445]), .A2(n7271), .ZN(n5115) );
  NAND2_X2 U3992 ( .A1(n5117), .A2(n5118), .ZN(w_d[444]) );
  NAND2_X2 U3993 ( .A1(w_q[412]), .A2(n7218), .ZN(n5118) );
  NAND2_X2 U3994 ( .A1(w_q[444]), .A2(n7271), .ZN(n5117) );
  NAND2_X2 U3995 ( .A1(n5119), .A2(n5120), .ZN(w_d[443]) );
  NAND2_X2 U3996 ( .A1(w_q[411]), .A2(n7218), .ZN(n5120) );
  NAND2_X2 U3997 ( .A1(w_q[443]), .A2(n7271), .ZN(n5119) );
  NAND2_X2 U3998 ( .A1(n5121), .A2(n5122), .ZN(w_d[442]) );
  NAND2_X2 U3999 ( .A1(w_q[410]), .A2(n7218), .ZN(n5122) );
  NAND2_X2 U4000 ( .A1(w_q[442]), .A2(n7271), .ZN(n5121) );
  NAND2_X2 U4001 ( .A1(n5123), .A2(n5124), .ZN(w_d[441]) );
  NAND2_X2 U4002 ( .A1(w_q[409]), .A2(n7218), .ZN(n5124) );
  NAND2_X2 U4003 ( .A1(w_q[441]), .A2(n7271), .ZN(n5123) );
  NAND2_X2 U4004 ( .A1(n5125), .A2(n5126), .ZN(w_d[440]) );
  NAND2_X2 U4005 ( .A1(w_q[408]), .A2(n7218), .ZN(n5126) );
  NAND2_X2 U4006 ( .A1(w_q[440]), .A2(n7271), .ZN(n5125) );
  NAND2_X2 U4007 ( .A1(n5127), .A2(n5128), .ZN(w_d[43]) );
  NAND2_X2 U4008 ( .A1(w_q[11]), .A2(n7216), .ZN(n5128) );
  NAND2_X2 U4009 ( .A1(w_q[43]), .A2(n7271), .ZN(n5127) );
  NAND2_X2 U4010 ( .A1(n5129), .A2(n5130), .ZN(w_d[439]) );
  NAND2_X2 U4011 ( .A1(w_q[407]), .A2(n7225), .ZN(n5130) );
  NAND2_X2 U4012 ( .A1(w_q[439]), .A2(n7271), .ZN(n5129) );
  NAND2_X2 U4013 ( .A1(n5131), .A2(n5132), .ZN(w_d[438]) );
  NAND2_X2 U4014 ( .A1(w_q[406]), .A2(n7223), .ZN(n5132) );
  NAND2_X2 U4015 ( .A1(w_q[438]), .A2(n7271), .ZN(n5131) );
  NAND2_X2 U4016 ( .A1(n5133), .A2(n5134), .ZN(w_d[437]) );
  NAND2_X2 U4017 ( .A1(w_q[405]), .A2(n7222), .ZN(n5134) );
  NAND2_X2 U4018 ( .A1(w_q[437]), .A2(n7271), .ZN(n5133) );
  NAND2_X2 U4019 ( .A1(n5135), .A2(n5136), .ZN(w_d[436]) );
  NAND2_X2 U4020 ( .A1(w_q[404]), .A2(n7226), .ZN(n5136) );
  NAND2_X2 U4021 ( .A1(w_q[436]), .A2(n7270), .ZN(n5135) );
  NAND2_X2 U4022 ( .A1(n5137), .A2(n5138), .ZN(w_d[435]) );
  NAND2_X2 U4023 ( .A1(w_q[403]), .A2(n7220), .ZN(n5138) );
  NAND2_X2 U4024 ( .A1(w_q[435]), .A2(n7270), .ZN(n5137) );
  NAND2_X2 U4025 ( .A1(n5139), .A2(n5140), .ZN(w_d[434]) );
  NAND2_X2 U4026 ( .A1(w_q[402]), .A2(n7219), .ZN(n5140) );
  NAND2_X2 U4027 ( .A1(w_q[434]), .A2(n7270), .ZN(n5139) );
  NAND2_X2 U4028 ( .A1(n5141), .A2(n5142), .ZN(w_d[433]) );
  NAND2_X2 U4029 ( .A1(w_q[401]), .A2(n7218), .ZN(n5142) );
  NAND2_X2 U4030 ( .A1(w_q[433]), .A2(n7270), .ZN(n5141) );
  NAND2_X2 U4031 ( .A1(n5143), .A2(n5144), .ZN(w_d[432]) );
  NAND2_X2 U4032 ( .A1(w_q[400]), .A2(n7217), .ZN(n5144) );
  NAND2_X2 U4033 ( .A1(w_q[432]), .A2(n7270), .ZN(n5143) );
  NAND2_X2 U4034 ( .A1(n5145), .A2(n5146), .ZN(w_d[431]) );
  NAND2_X2 U4035 ( .A1(w_q[399]), .A2(n7221), .ZN(n5146) );
  NAND2_X2 U4036 ( .A1(w_q[431]), .A2(n7270), .ZN(n5145) );
  NAND2_X2 U4037 ( .A1(n5147), .A2(n5148), .ZN(w_d[430]) );
  NAND2_X2 U4038 ( .A1(w_q[398]), .A2(n7224), .ZN(n5148) );
  NAND2_X2 U4039 ( .A1(w_q[430]), .A2(n7270), .ZN(n5147) );
  NAND2_X2 U4040 ( .A1(n5149), .A2(n5150), .ZN(w_d[42]) );
  NAND2_X2 U4041 ( .A1(w_q[10]), .A2(n7211), .ZN(n5150) );
  NAND2_X2 U4042 ( .A1(w_q[42]), .A2(n7270), .ZN(n5149) );
  NAND2_X2 U4043 ( .A1(n5151), .A2(n5152), .ZN(w_d[429]) );
  NAND2_X2 U4044 ( .A1(w_q[397]), .A2(n7211), .ZN(n5152) );
  NAND2_X2 U4045 ( .A1(w_q[429]), .A2(n7270), .ZN(n5151) );
  NAND2_X2 U4046 ( .A1(n5153), .A2(n5154), .ZN(w_d[428]) );
  NAND2_X2 U4047 ( .A1(w_q[396]), .A2(n7211), .ZN(n5154) );
  NAND2_X2 U4048 ( .A1(w_q[428]), .A2(n7270), .ZN(n5153) );
  NAND2_X2 U4049 ( .A1(n5155), .A2(n5156), .ZN(w_d[427]) );
  NAND2_X2 U4050 ( .A1(w_q[395]), .A2(n7211), .ZN(n5156) );
  NAND2_X2 U4051 ( .A1(w_q[427]), .A2(n7270), .ZN(n5155) );
  NAND2_X2 U4052 ( .A1(n5157), .A2(n5158), .ZN(w_d[426]) );
  NAND2_X2 U4053 ( .A1(w_q[394]), .A2(n7211), .ZN(n5158) );
  NAND2_X2 U4054 ( .A1(w_q[426]), .A2(n7269), .ZN(n5157) );
  NAND2_X2 U4055 ( .A1(n5159), .A2(n5160), .ZN(w_d[425]) );
  NAND2_X2 U4056 ( .A1(w_q[393]), .A2(n7211), .ZN(n5160) );
  NAND2_X2 U4057 ( .A1(w_q[425]), .A2(n7269), .ZN(n5159) );
  NAND2_X2 U4058 ( .A1(n5161), .A2(n5162), .ZN(w_d[424]) );
  NAND2_X2 U4059 ( .A1(w_q[392]), .A2(n7211), .ZN(n5162) );
  NAND2_X2 U4060 ( .A1(w_q[424]), .A2(n7269), .ZN(n5161) );
  NAND2_X2 U4061 ( .A1(n5163), .A2(n5164), .ZN(w_d[423]) );
  NAND2_X2 U4062 ( .A1(w_q[391]), .A2(n7211), .ZN(n5164) );
  NAND2_X2 U4063 ( .A1(w_q[423]), .A2(n7269), .ZN(n5163) );
  NAND2_X2 U4064 ( .A1(n5165), .A2(n5166), .ZN(w_d[422]) );
  NAND2_X2 U4065 ( .A1(w_q[390]), .A2(n7211), .ZN(n5166) );
  NAND2_X2 U4066 ( .A1(w_q[422]), .A2(n7269), .ZN(n5165) );
  NAND2_X2 U4067 ( .A1(n5167), .A2(n5168), .ZN(w_d[421]) );
  NAND2_X2 U4068 ( .A1(w_q[389]), .A2(n7211), .ZN(n5168) );
  NAND2_X2 U4069 ( .A1(w_q[421]), .A2(n7269), .ZN(n5167) );
  NAND2_X2 U4070 ( .A1(n5169), .A2(n5170), .ZN(w_d[420]) );
  NAND2_X2 U4071 ( .A1(w_q[388]), .A2(n7211), .ZN(n5170) );
  NAND2_X2 U4072 ( .A1(w_q[420]), .A2(n7269), .ZN(n5169) );
  NAND2_X2 U4073 ( .A1(n5171), .A2(n5172), .ZN(w_d[41]) );
  NAND2_X2 U4074 ( .A1(w_q[9]), .A2(n7210), .ZN(n5172) );
  NAND2_X2 U4075 ( .A1(w_q[41]), .A2(n7269), .ZN(n5171) );
  NAND2_X2 U4076 ( .A1(n5173), .A2(n5174), .ZN(w_d[419]) );
  NAND2_X2 U4077 ( .A1(w_q[387]), .A2(n7210), .ZN(n5174) );
  NAND2_X2 U4078 ( .A1(w_q[419]), .A2(n7269), .ZN(n5173) );
  NAND2_X2 U4079 ( .A1(n5175), .A2(n5176), .ZN(w_d[418]) );
  NAND2_X2 U4080 ( .A1(w_q[386]), .A2(n7210), .ZN(n5176) );
  NAND2_X2 U4081 ( .A1(w_q[418]), .A2(n7269), .ZN(n5175) );
  NAND2_X2 U4082 ( .A1(n5177), .A2(n5178), .ZN(w_d[417]) );
  NAND2_X2 U4083 ( .A1(w_q[385]), .A2(n7210), .ZN(n5178) );
  NAND2_X2 U4084 ( .A1(w_q[417]), .A2(n7269), .ZN(n5177) );
  NAND2_X2 U4085 ( .A1(n5179), .A2(n5180), .ZN(w_d[416]) );
  NAND2_X2 U4086 ( .A1(w_q[384]), .A2(n7210), .ZN(n5180) );
  NAND2_X2 U4087 ( .A1(w_q[416]), .A2(n7268), .ZN(n5179) );
  NAND2_X2 U4088 ( .A1(n5181), .A2(n5182), .ZN(w_d[415]) );
  NAND2_X2 U4089 ( .A1(w_q[383]), .A2(n7210), .ZN(n5182) );
  NAND2_X2 U4090 ( .A1(w_q[415]), .A2(n7268), .ZN(n5181) );
  NAND2_X2 U4091 ( .A1(n5183), .A2(n5184), .ZN(w_d[414]) );
  NAND2_X2 U4092 ( .A1(w_q[382]), .A2(n7210), .ZN(n5184) );
  NAND2_X2 U4093 ( .A1(w_q[414]), .A2(n7268), .ZN(n5183) );
  NAND2_X2 U4094 ( .A1(n5185), .A2(n5186), .ZN(w_d[413]) );
  NAND2_X2 U4095 ( .A1(w_q[381]), .A2(n7210), .ZN(n5186) );
  NAND2_X2 U4096 ( .A1(w_q[413]), .A2(n7268), .ZN(n5185) );
  NAND2_X2 U4097 ( .A1(n5187), .A2(n5188), .ZN(w_d[412]) );
  NAND2_X2 U4098 ( .A1(w_q[380]), .A2(n7210), .ZN(n5188) );
  NAND2_X2 U4099 ( .A1(w_q[412]), .A2(n7268), .ZN(n5187) );
  NAND2_X2 U4100 ( .A1(n5189), .A2(n5190), .ZN(w_d[411]) );
  NAND2_X2 U4101 ( .A1(w_q[379]), .A2(n7210), .ZN(n5190) );
  NAND2_X2 U4102 ( .A1(w_q[411]), .A2(n7268), .ZN(n5189) );
  NAND2_X2 U4103 ( .A1(n5191), .A2(n5192), .ZN(w_d[410]) );
  NAND2_X2 U4104 ( .A1(w_q[378]), .A2(n7210), .ZN(n5192) );
  NAND2_X2 U4105 ( .A1(w_q[410]), .A2(n7268), .ZN(n5191) );
  NAND2_X2 U4106 ( .A1(n5193), .A2(n5194), .ZN(w_d[40]) );
  NAND2_X2 U4107 ( .A1(w_q[8]), .A2(n7209), .ZN(n5194) );
  NAND2_X2 U4108 ( .A1(w_q[40]), .A2(n7268), .ZN(n5193) );
  NAND2_X2 U4109 ( .A1(n5195), .A2(n5196), .ZN(w_d[409]) );
  NAND2_X2 U4110 ( .A1(w_q[377]), .A2(n7209), .ZN(n5196) );
  NAND2_X2 U4111 ( .A1(w_q[409]), .A2(n7268), .ZN(n5195) );
  NAND2_X2 U4112 ( .A1(n5197), .A2(n5198), .ZN(w_d[408]) );
  NAND2_X2 U4113 ( .A1(w_q[376]), .A2(n7209), .ZN(n5198) );
  NAND2_X2 U4114 ( .A1(w_q[408]), .A2(n7268), .ZN(n5197) );
  NAND2_X2 U4115 ( .A1(n5199), .A2(n5200), .ZN(w_d[407]) );
  NAND2_X2 U4116 ( .A1(w_q[375]), .A2(n7209), .ZN(n5200) );
  NAND2_X2 U4117 ( .A1(w_q[407]), .A2(n7268), .ZN(n5199) );
  NAND2_X2 U4118 ( .A1(n5201), .A2(n5202), .ZN(w_d[406]) );
  NAND2_X2 U4119 ( .A1(w_q[374]), .A2(n7209), .ZN(n5202) );
  NAND2_X2 U4120 ( .A1(w_q[406]), .A2(n7267), .ZN(n5201) );
  NAND2_X2 U4121 ( .A1(n5203), .A2(n5204), .ZN(w_d[405]) );
  NAND2_X2 U4122 ( .A1(w_q[373]), .A2(n7209), .ZN(n5204) );
  NAND2_X2 U4123 ( .A1(w_q[405]), .A2(n7267), .ZN(n5203) );
  NAND2_X2 U4124 ( .A1(n5205), .A2(n5206), .ZN(w_d[404]) );
  NAND2_X2 U4125 ( .A1(w_q[372]), .A2(n7209), .ZN(n5206) );
  NAND2_X2 U4126 ( .A1(w_q[404]), .A2(n7267), .ZN(n5205) );
  NAND2_X2 U4127 ( .A1(n5207), .A2(n5208), .ZN(w_d[403]) );
  NAND2_X2 U4128 ( .A1(w_q[371]), .A2(n7209), .ZN(n5208) );
  NAND2_X2 U4129 ( .A1(w_q[403]), .A2(n7267), .ZN(n5207) );
  NAND2_X2 U4130 ( .A1(n5209), .A2(n5210), .ZN(w_d[402]) );
  NAND2_X2 U4131 ( .A1(w_q[370]), .A2(n7209), .ZN(n5210) );
  NAND2_X2 U4132 ( .A1(w_q[402]), .A2(n7267), .ZN(n5209) );
  NAND2_X2 U4133 ( .A1(n5211), .A2(n5212), .ZN(w_d[401]) );
  NAND2_X2 U4134 ( .A1(w_q[369]), .A2(n7209), .ZN(n5212) );
  NAND2_X2 U4135 ( .A1(w_q[401]), .A2(n7267), .ZN(n5211) );
  NAND2_X2 U4136 ( .A1(n5213), .A2(n5214), .ZN(w_d[400]) );
  NAND2_X2 U4137 ( .A1(w_q[368]), .A2(n7209), .ZN(n5214) );
  NAND2_X2 U4138 ( .A1(w_q[400]), .A2(n7267), .ZN(n5213) );
  NAND2_X2 U4140 ( .A1(w[3]), .A2(n7159), .ZN(n5217) );
  NAND2_X2 U4141 ( .A1(w_q[3]), .A2(n7267), .ZN(n5216) );
  NAND2_X2 U4143 ( .A1(n5218), .A2(n5219), .ZN(w_d[39]) );
  NAND2_X2 U4144 ( .A1(w_q[7]), .A2(n7208), .ZN(n5219) );
  NAND2_X2 U4145 ( .A1(w_q[39]), .A2(n7267), .ZN(n5218) );
  NAND2_X2 U4146 ( .A1(n5220), .A2(n5221), .ZN(w_d[399]) );
  NAND2_X2 U4147 ( .A1(w_q[367]), .A2(n7208), .ZN(n5221) );
  NAND2_X2 U4148 ( .A1(w_q[399]), .A2(n7267), .ZN(n5220) );
  NAND2_X2 U4149 ( .A1(n5222), .A2(n5223), .ZN(w_d[398]) );
  NAND2_X2 U4150 ( .A1(w_q[366]), .A2(n7208), .ZN(n5223) );
  NAND2_X2 U4151 ( .A1(w_q[398]), .A2(n7267), .ZN(n5222) );
  NAND2_X2 U4152 ( .A1(n5224), .A2(n5225), .ZN(w_d[397]) );
  NAND2_X2 U4153 ( .A1(w_q[365]), .A2(n7208), .ZN(n5225) );
  NAND2_X2 U4154 ( .A1(w_q[397]), .A2(n7266), .ZN(n5224) );
  NAND2_X2 U4155 ( .A1(n5226), .A2(n5227), .ZN(w_d[396]) );
  NAND2_X2 U4156 ( .A1(w_q[364]), .A2(n7208), .ZN(n5227) );
  NAND2_X2 U4157 ( .A1(w_q[396]), .A2(n7266), .ZN(n5226) );
  NAND2_X2 U4158 ( .A1(n5228), .A2(n5229), .ZN(w_d[395]) );
  NAND2_X2 U4159 ( .A1(w_q[363]), .A2(n7208), .ZN(n5229) );
  NAND2_X2 U4160 ( .A1(w_q[395]), .A2(n7266), .ZN(n5228) );
  NAND2_X2 U4161 ( .A1(n5230), .A2(n5231), .ZN(w_d[394]) );
  NAND2_X2 U4162 ( .A1(w_q[362]), .A2(n7208), .ZN(n5231) );
  NAND2_X2 U4163 ( .A1(w_q[394]), .A2(n7266), .ZN(n5230) );
  NAND2_X2 U4164 ( .A1(n5232), .A2(n5233), .ZN(w_d[393]) );
  NAND2_X2 U4165 ( .A1(w_q[361]), .A2(n7208), .ZN(n5233) );
  NAND2_X2 U4166 ( .A1(w_q[393]), .A2(n7266), .ZN(n5232) );
  NAND2_X2 U4167 ( .A1(n5234), .A2(n5235), .ZN(w_d[392]) );
  NAND2_X2 U4168 ( .A1(w_q[360]), .A2(n7208), .ZN(n5235) );
  NAND2_X2 U4169 ( .A1(w_q[392]), .A2(n7266), .ZN(n5234) );
  NAND2_X2 U4170 ( .A1(n5236), .A2(n5237), .ZN(w_d[391]) );
  NAND2_X2 U4171 ( .A1(w_q[359]), .A2(n7208), .ZN(n5237) );
  NAND2_X2 U4172 ( .A1(w_q[391]), .A2(n7266), .ZN(n5236) );
  NAND2_X2 U4173 ( .A1(n5238), .A2(n5239), .ZN(w_d[390]) );
  NAND2_X2 U4174 ( .A1(w_q[358]), .A2(n7208), .ZN(n5239) );
  NAND2_X2 U4175 ( .A1(w_q[390]), .A2(n7266), .ZN(n5238) );
  NAND2_X2 U4176 ( .A1(n5240), .A2(n5241), .ZN(w_d[38]) );
  NAND2_X2 U4177 ( .A1(w_q[6]), .A2(n7207), .ZN(n5241) );
  NAND2_X2 U4178 ( .A1(w_q[38]), .A2(n7266), .ZN(n5240) );
  NAND2_X2 U4179 ( .A1(n5242), .A2(n5243), .ZN(w_d[389]) );
  NAND2_X2 U4180 ( .A1(w_q[357]), .A2(n7207), .ZN(n5243) );
  NAND2_X2 U4181 ( .A1(w_q[389]), .A2(n7266), .ZN(n5242) );
  NAND2_X2 U4182 ( .A1(n5244), .A2(n5245), .ZN(w_d[388]) );
  NAND2_X2 U4183 ( .A1(w_q[356]), .A2(n7207), .ZN(n5245) );
  NAND2_X2 U4184 ( .A1(w_q[388]), .A2(n7266), .ZN(n5244) );
  NAND2_X2 U4185 ( .A1(n5246), .A2(n5247), .ZN(w_d[387]) );
  NAND2_X2 U4186 ( .A1(w_q[355]), .A2(n7207), .ZN(n5247) );
  NAND2_X2 U4187 ( .A1(w_q[387]), .A2(n7265), .ZN(n5246) );
  NAND2_X2 U4188 ( .A1(n5248), .A2(n5249), .ZN(w_d[386]) );
  NAND2_X2 U4189 ( .A1(w_q[354]), .A2(n7207), .ZN(n5249) );
  NAND2_X2 U4190 ( .A1(w_q[386]), .A2(n7265), .ZN(n5248) );
  NAND2_X2 U4191 ( .A1(n5250), .A2(n5251), .ZN(w_d[385]) );
  NAND2_X2 U4192 ( .A1(w_q[353]), .A2(n7207), .ZN(n5251) );
  NAND2_X2 U4193 ( .A1(w_q[385]), .A2(n7265), .ZN(n5250) );
  NAND2_X2 U4194 ( .A1(n5252), .A2(n5253), .ZN(w_d[384]) );
  NAND2_X2 U4195 ( .A1(w_q[352]), .A2(n7207), .ZN(n5253) );
  NAND2_X2 U4196 ( .A1(w_q[384]), .A2(n7265), .ZN(n5252) );
  NAND2_X2 U4197 ( .A1(n5254), .A2(n5255), .ZN(w_d[383]) );
  NAND2_X2 U4198 ( .A1(w_q[351]), .A2(n7207), .ZN(n5255) );
  NAND2_X2 U4199 ( .A1(w_q[383]), .A2(n7265), .ZN(n5254) );
  NAND2_X2 U4200 ( .A1(n5256), .A2(n5257), .ZN(w_d[382]) );
  NAND2_X2 U4201 ( .A1(w_q[350]), .A2(n7207), .ZN(n5257) );
  NAND2_X2 U4202 ( .A1(w_q[382]), .A2(n7265), .ZN(n5256) );
  NAND2_X2 U4203 ( .A1(n5258), .A2(n5259), .ZN(w_d[381]) );
  NAND2_X2 U4204 ( .A1(w_q[349]), .A2(n7207), .ZN(n5259) );
  NAND2_X2 U4205 ( .A1(w_q[381]), .A2(n7265), .ZN(n5258) );
  NAND2_X2 U4206 ( .A1(n5260), .A2(n5261), .ZN(w_d[380]) );
  NAND2_X2 U4207 ( .A1(w_q[348]), .A2(n7207), .ZN(n5261) );
  NAND2_X2 U4208 ( .A1(w_q[380]), .A2(n7265), .ZN(n5260) );
  NAND2_X2 U4209 ( .A1(n5262), .A2(n5263), .ZN(w_d[37]) );
  NAND2_X2 U4210 ( .A1(w_q[5]), .A2(n7206), .ZN(n5263) );
  NAND2_X2 U4211 ( .A1(w_q[37]), .A2(n7265), .ZN(n5262) );
  NAND2_X2 U4212 ( .A1(n5264), .A2(n5265), .ZN(w_d[379]) );
  NAND2_X2 U4213 ( .A1(w_q[347]), .A2(n7206), .ZN(n5265) );
  NAND2_X2 U4214 ( .A1(w_q[379]), .A2(n7265), .ZN(n5264) );
  NAND2_X2 U4215 ( .A1(n5266), .A2(n5267), .ZN(w_d[378]) );
  NAND2_X2 U4216 ( .A1(w_q[346]), .A2(n7206), .ZN(n5267) );
  NAND2_X2 U4217 ( .A1(w_q[378]), .A2(n7265), .ZN(n5266) );
  NAND2_X2 U4218 ( .A1(n5268), .A2(n5269), .ZN(w_d[377]) );
  NAND2_X2 U4219 ( .A1(w_q[345]), .A2(n7206), .ZN(n5269) );
  NAND2_X2 U4220 ( .A1(w_q[377]), .A2(n7264), .ZN(n5268) );
  NAND2_X2 U4221 ( .A1(n5270), .A2(n5271), .ZN(w_d[376]) );
  NAND2_X2 U4222 ( .A1(w_q[344]), .A2(n7206), .ZN(n5271) );
  NAND2_X2 U4223 ( .A1(w_q[376]), .A2(n7264), .ZN(n5270) );
  NAND2_X2 U4224 ( .A1(n5272), .A2(n5273), .ZN(w_d[375]) );
  NAND2_X2 U4225 ( .A1(w_q[343]), .A2(n7206), .ZN(n5273) );
  NAND2_X2 U4226 ( .A1(w_q[375]), .A2(n7264), .ZN(n5272) );
  NAND2_X2 U4227 ( .A1(n5274), .A2(n5275), .ZN(w_d[374]) );
  NAND2_X2 U4228 ( .A1(w_q[342]), .A2(n7206), .ZN(n5275) );
  NAND2_X2 U4229 ( .A1(w_q[374]), .A2(n7264), .ZN(n5274) );
  NAND2_X2 U4230 ( .A1(n5276), .A2(n5277), .ZN(w_d[373]) );
  NAND2_X2 U4231 ( .A1(w_q[341]), .A2(n7206), .ZN(n5277) );
  NAND2_X2 U4232 ( .A1(w_q[373]), .A2(n7264), .ZN(n5276) );
  NAND2_X2 U4233 ( .A1(n5278), .A2(n5279), .ZN(w_d[372]) );
  NAND2_X2 U4234 ( .A1(w_q[340]), .A2(n7206), .ZN(n5279) );
  NAND2_X2 U4235 ( .A1(w_q[372]), .A2(n7264), .ZN(n5278) );
  NAND2_X2 U4236 ( .A1(n5280), .A2(n5281), .ZN(w_d[371]) );
  NAND2_X2 U4237 ( .A1(w_q[339]), .A2(n7206), .ZN(n5281) );
  NAND2_X2 U4238 ( .A1(w_q[371]), .A2(n7264), .ZN(n5280) );
  NAND2_X2 U4239 ( .A1(n5282), .A2(n5283), .ZN(w_d[370]) );
  NAND2_X2 U4240 ( .A1(w_q[338]), .A2(n7206), .ZN(n5283) );
  NAND2_X2 U4241 ( .A1(w_q[370]), .A2(n7264), .ZN(n5282) );
  NAND2_X2 U4242 ( .A1(n5284), .A2(n5285), .ZN(w_d[36]) );
  NAND2_X2 U4243 ( .A1(w_q[4]), .A2(n7205), .ZN(n5285) );
  NAND2_X2 U4244 ( .A1(w_q[36]), .A2(n7264), .ZN(n5284) );
  NAND2_X2 U4245 ( .A1(n5286), .A2(n5287), .ZN(w_d[369]) );
  NAND2_X2 U4246 ( .A1(w_q[337]), .A2(n7205), .ZN(n5287) );
  NAND2_X2 U4247 ( .A1(w_q[369]), .A2(n7264), .ZN(n5286) );
  NAND2_X2 U4248 ( .A1(n5288), .A2(n5289), .ZN(w_d[368]) );
  NAND2_X2 U4249 ( .A1(w_q[336]), .A2(n7205), .ZN(n5289) );
  NAND2_X2 U4250 ( .A1(w_q[368]), .A2(n7264), .ZN(n5288) );
  NAND2_X2 U4251 ( .A1(n5290), .A2(n5291), .ZN(w_d[367]) );
  NAND2_X2 U4252 ( .A1(w_q[335]), .A2(n7205), .ZN(n5291) );
  NAND2_X2 U4253 ( .A1(w_q[367]), .A2(n7263), .ZN(n5290) );
  NAND2_X2 U4254 ( .A1(n5292), .A2(n5293), .ZN(w_d[366]) );
  NAND2_X2 U4255 ( .A1(w_q[334]), .A2(n7205), .ZN(n5293) );
  NAND2_X2 U4256 ( .A1(w_q[366]), .A2(n7263), .ZN(n5292) );
  NAND2_X2 U4257 ( .A1(n5294), .A2(n5295), .ZN(w_d[365]) );
  NAND2_X2 U4258 ( .A1(w_q[333]), .A2(n7205), .ZN(n5295) );
  NAND2_X2 U4259 ( .A1(w_q[365]), .A2(n7263), .ZN(n5294) );
  NAND2_X2 U4260 ( .A1(n5296), .A2(n5297), .ZN(w_d[364]) );
  NAND2_X2 U4261 ( .A1(w_q[332]), .A2(n7205), .ZN(n5297) );
  NAND2_X2 U4262 ( .A1(w_q[364]), .A2(n7263), .ZN(n5296) );
  NAND2_X2 U4263 ( .A1(n5298), .A2(n5299), .ZN(w_d[363]) );
  NAND2_X2 U4264 ( .A1(w_q[331]), .A2(n7205), .ZN(n5299) );
  NAND2_X2 U4265 ( .A1(w_q[363]), .A2(n7263), .ZN(n5298) );
  NAND2_X2 U4266 ( .A1(n5300), .A2(n5301), .ZN(w_d[362]) );
  NAND2_X2 U4267 ( .A1(w_q[330]), .A2(n7205), .ZN(n5301) );
  NAND2_X2 U4268 ( .A1(w_q[362]), .A2(n7263), .ZN(n5300) );
  NAND2_X2 U4269 ( .A1(n5302), .A2(n5303), .ZN(w_d[361]) );
  NAND2_X2 U4270 ( .A1(w_q[329]), .A2(n7205), .ZN(n5303) );
  NAND2_X2 U4271 ( .A1(w_q[361]), .A2(n7263), .ZN(n5302) );
  NAND2_X2 U4272 ( .A1(n5304), .A2(n5305), .ZN(w_d[360]) );
  NAND2_X2 U4273 ( .A1(w_q[328]), .A2(n7205), .ZN(n5305) );
  NAND2_X2 U4274 ( .A1(w_q[360]), .A2(n7263), .ZN(n5304) );
  NAND2_X2 U4275 ( .A1(n5306), .A2(n5307), .ZN(w_d[35]) );
  NAND2_X2 U4276 ( .A1(w_q[3]), .A2(n7204), .ZN(n5307) );
  NAND2_X2 U4277 ( .A1(w_q[35]), .A2(n7263), .ZN(n5306) );
  NAND2_X2 U4278 ( .A1(n5308), .A2(n5309), .ZN(w_d[359]) );
  NAND2_X2 U4279 ( .A1(w_q[327]), .A2(n7204), .ZN(n5309) );
  NAND2_X2 U4280 ( .A1(w_q[359]), .A2(n7263), .ZN(n5308) );
  NAND2_X2 U4281 ( .A1(n5310), .A2(n5311), .ZN(w_d[358]) );
  NAND2_X2 U4282 ( .A1(w_q[326]), .A2(n7204), .ZN(n5311) );
  NAND2_X2 U4283 ( .A1(w_q[358]), .A2(n7263), .ZN(n5310) );
  NAND2_X2 U4284 ( .A1(n5312), .A2(n5313), .ZN(w_d[357]) );
  NAND2_X2 U4285 ( .A1(w_q[325]), .A2(n7204), .ZN(n5313) );
  NAND2_X2 U4286 ( .A1(w_q[357]), .A2(n7262), .ZN(n5312) );
  NAND2_X2 U4287 ( .A1(n5314), .A2(n5315), .ZN(w_d[356]) );
  NAND2_X2 U4288 ( .A1(w_q[324]), .A2(n7204), .ZN(n5315) );
  NAND2_X2 U4289 ( .A1(w_q[356]), .A2(n7262), .ZN(n5314) );
  NAND2_X2 U4290 ( .A1(n5316), .A2(n5317), .ZN(w_d[355]) );
  NAND2_X2 U4291 ( .A1(w_q[323]), .A2(n7204), .ZN(n5317) );
  NAND2_X2 U4292 ( .A1(w_q[355]), .A2(n7262), .ZN(n5316) );
  NAND2_X2 U4293 ( .A1(n5318), .A2(n5319), .ZN(w_d[354]) );
  NAND2_X2 U4294 ( .A1(w_q[322]), .A2(n7204), .ZN(n5319) );
  NAND2_X2 U4295 ( .A1(w_q[354]), .A2(n7262), .ZN(n5318) );
  NAND2_X2 U4296 ( .A1(n5320), .A2(n5321), .ZN(w_d[353]) );
  NAND2_X2 U4297 ( .A1(w_q[321]), .A2(n7204), .ZN(n5321) );
  NAND2_X2 U4298 ( .A1(w_q[353]), .A2(n7262), .ZN(n5320) );
  NAND2_X2 U4299 ( .A1(n5322), .A2(n5323), .ZN(w_d[352]) );
  NAND2_X2 U4300 ( .A1(w_q[320]), .A2(n7204), .ZN(n5323) );
  NAND2_X2 U4301 ( .A1(w_q[352]), .A2(n7262), .ZN(n5322) );
  NAND2_X2 U4302 ( .A1(n5324), .A2(n5325), .ZN(w_d[351]) );
  NAND2_X2 U4303 ( .A1(w_q[319]), .A2(n7204), .ZN(n5325) );
  NAND2_X2 U4304 ( .A1(w_q[351]), .A2(n7262), .ZN(n5324) );
  NAND2_X2 U4305 ( .A1(n5326), .A2(n5327), .ZN(w_d[350]) );
  NAND2_X2 U4306 ( .A1(w_q[318]), .A2(n7204), .ZN(n5327) );
  NAND2_X2 U4307 ( .A1(w_q[350]), .A2(n7262), .ZN(n5326) );
  NAND2_X2 U4308 ( .A1(n5328), .A2(n5329), .ZN(w_d[34]) );
  NAND2_X2 U4309 ( .A1(w_q[2]), .A2(n7203), .ZN(n5329) );
  NAND2_X2 U4310 ( .A1(w_q[34]), .A2(n7262), .ZN(n5328) );
  NAND2_X2 U4311 ( .A1(n5330), .A2(n5331), .ZN(w_d[349]) );
  NAND2_X2 U4312 ( .A1(w_q[317]), .A2(n7203), .ZN(n5331) );
  NAND2_X2 U4313 ( .A1(w_q[349]), .A2(n7262), .ZN(n5330) );
  NAND2_X2 U4314 ( .A1(n5332), .A2(n5333), .ZN(w_d[348]) );
  NAND2_X2 U4315 ( .A1(w_q[316]), .A2(n7203), .ZN(n5333) );
  NAND2_X2 U4316 ( .A1(w_q[348]), .A2(n7262), .ZN(n5332) );
  NAND2_X2 U4317 ( .A1(n5334), .A2(n5335), .ZN(w_d[347]) );
  NAND2_X2 U4318 ( .A1(w_q[315]), .A2(n7203), .ZN(n5335) );
  NAND2_X2 U4319 ( .A1(w_q[347]), .A2(n7261), .ZN(n5334) );
  NAND2_X2 U4320 ( .A1(n5336), .A2(n5337), .ZN(w_d[346]) );
  NAND2_X2 U4321 ( .A1(w_q[314]), .A2(n7203), .ZN(n5337) );
  NAND2_X2 U4322 ( .A1(w_q[346]), .A2(n7261), .ZN(n5336) );
  NAND2_X2 U4323 ( .A1(n5338), .A2(n5339), .ZN(w_d[345]) );
  NAND2_X2 U4324 ( .A1(w_q[313]), .A2(n7203), .ZN(n5339) );
  NAND2_X2 U4325 ( .A1(w_q[345]), .A2(n7261), .ZN(n5338) );
  NAND2_X2 U4326 ( .A1(n5340), .A2(n5341), .ZN(w_d[344]) );
  NAND2_X2 U4327 ( .A1(w_q[312]), .A2(n7203), .ZN(n5341) );
  NAND2_X2 U4328 ( .A1(w_q[344]), .A2(n7261), .ZN(n5340) );
  NAND2_X2 U4329 ( .A1(n5342), .A2(n5343), .ZN(w_d[343]) );
  NAND2_X2 U4330 ( .A1(w_q[311]), .A2(n7203), .ZN(n5343) );
  NAND2_X2 U4331 ( .A1(w_q[343]), .A2(n7261), .ZN(n5342) );
  NAND2_X2 U4332 ( .A1(n5344), .A2(n5345), .ZN(w_d[342]) );
  NAND2_X2 U4333 ( .A1(w_q[310]), .A2(n7203), .ZN(n5345) );
  NAND2_X2 U4334 ( .A1(w_q[342]), .A2(n7261), .ZN(n5344) );
  NAND2_X2 U4335 ( .A1(n5346), .A2(n5347), .ZN(w_d[341]) );
  NAND2_X2 U4336 ( .A1(w_q[309]), .A2(n7203), .ZN(n5347) );
  NAND2_X2 U4337 ( .A1(w_q[341]), .A2(n7261), .ZN(n5346) );
  NAND2_X2 U4338 ( .A1(n5348), .A2(n5349), .ZN(w_d[340]) );
  NAND2_X2 U4339 ( .A1(w_q[308]), .A2(n7203), .ZN(n5349) );
  NAND2_X2 U4340 ( .A1(w_q[340]), .A2(n7261), .ZN(n5348) );
  NAND2_X2 U4341 ( .A1(n5350), .A2(n5351), .ZN(w_d[33]) );
  NAND2_X2 U4342 ( .A1(w_q[1]), .A2(n7202), .ZN(n5351) );
  NAND2_X2 U4343 ( .A1(w_q[33]), .A2(n7261), .ZN(n5350) );
  NAND2_X2 U4344 ( .A1(n5352), .A2(n5353), .ZN(w_d[339]) );
  NAND2_X2 U4345 ( .A1(w_q[307]), .A2(n7202), .ZN(n5353) );
  NAND2_X2 U4346 ( .A1(w_q[339]), .A2(n7261), .ZN(n5352) );
  NAND2_X2 U4347 ( .A1(n5354), .A2(n5355), .ZN(w_d[338]) );
  NAND2_X2 U4348 ( .A1(w_q[306]), .A2(n7202), .ZN(n5355) );
  NAND2_X2 U4349 ( .A1(w_q[338]), .A2(n7261), .ZN(n5354) );
  NAND2_X2 U4350 ( .A1(n5356), .A2(n5357), .ZN(w_d[337]) );
  NAND2_X2 U4351 ( .A1(w_q[305]), .A2(n7202), .ZN(n5357) );
  NAND2_X2 U4352 ( .A1(w_q[337]), .A2(n7260), .ZN(n5356) );
  NAND2_X2 U4353 ( .A1(n5358), .A2(n5359), .ZN(w_d[336]) );
  NAND2_X2 U4354 ( .A1(w_q[304]), .A2(n7202), .ZN(n5359) );
  NAND2_X2 U4355 ( .A1(w_q[336]), .A2(n7260), .ZN(n5358) );
  NAND2_X2 U4356 ( .A1(n5360), .A2(n5361), .ZN(w_d[335]) );
  NAND2_X2 U4357 ( .A1(w_q[303]), .A2(n7202), .ZN(n5361) );
  NAND2_X2 U4358 ( .A1(w_q[335]), .A2(n7260), .ZN(n5360) );
  NAND2_X2 U4359 ( .A1(n5362), .A2(n5363), .ZN(w_d[334]) );
  NAND2_X2 U4360 ( .A1(w_q[302]), .A2(n7202), .ZN(n5363) );
  NAND2_X2 U4361 ( .A1(w_q[334]), .A2(n7260), .ZN(n5362) );
  NAND2_X2 U4362 ( .A1(n5364), .A2(n5365), .ZN(w_d[333]) );
  NAND2_X2 U4363 ( .A1(w_q[301]), .A2(n7202), .ZN(n5365) );
  NAND2_X2 U4364 ( .A1(w_q[333]), .A2(n7260), .ZN(n5364) );
  NAND2_X2 U4365 ( .A1(n5366), .A2(n5367), .ZN(w_d[332]) );
  NAND2_X2 U4366 ( .A1(w_q[300]), .A2(n7202), .ZN(n5367) );
  NAND2_X2 U4367 ( .A1(w_q[332]), .A2(n7260), .ZN(n5366) );
  NAND2_X2 U4368 ( .A1(n5368), .A2(n5369), .ZN(w_d[331]) );
  NAND2_X2 U4369 ( .A1(w_q[299]), .A2(n7202), .ZN(n5369) );
  NAND2_X2 U4370 ( .A1(w_q[331]), .A2(n7260), .ZN(n5368) );
  NAND2_X2 U4371 ( .A1(n5370), .A2(n5371), .ZN(w_d[330]) );
  NAND2_X2 U4372 ( .A1(w_q[298]), .A2(n7202), .ZN(n5371) );
  NAND2_X2 U4373 ( .A1(w_q[330]), .A2(n7260), .ZN(n5370) );
  NAND2_X2 U4374 ( .A1(n5372), .A2(n5373), .ZN(w_d[32]) );
  NAND2_X2 U4375 ( .A1(w_q[0]), .A2(n7201), .ZN(n5373) );
  NAND2_X2 U4376 ( .A1(w_q[32]), .A2(n7260), .ZN(n5372) );
  NAND2_X2 U4377 ( .A1(n5374), .A2(n5375), .ZN(w_d[329]) );
  NAND2_X2 U4378 ( .A1(w_q[297]), .A2(n7201), .ZN(n5375) );
  NAND2_X2 U4379 ( .A1(w_q[329]), .A2(n7260), .ZN(n5374) );
  NAND2_X2 U4380 ( .A1(n5376), .A2(n5377), .ZN(w_d[328]) );
  NAND2_X2 U4381 ( .A1(w_q[296]), .A2(n7201), .ZN(n5377) );
  NAND2_X2 U4382 ( .A1(w_q[328]), .A2(n7260), .ZN(n5376) );
  NAND2_X2 U4383 ( .A1(n5378), .A2(n5379), .ZN(w_d[327]) );
  NAND2_X2 U4384 ( .A1(w_q[295]), .A2(n7201), .ZN(n5379) );
  NAND2_X2 U4385 ( .A1(w_q[327]), .A2(n7259), .ZN(n5378) );
  NAND2_X2 U4386 ( .A1(n5380), .A2(n5381), .ZN(w_d[326]) );
  NAND2_X2 U4387 ( .A1(w_q[294]), .A2(n7201), .ZN(n5381) );
  NAND2_X2 U4388 ( .A1(w_q[326]), .A2(n7259), .ZN(n5380) );
  NAND2_X2 U4389 ( .A1(n5382), .A2(n5383), .ZN(w_d[325]) );
  NAND2_X2 U4390 ( .A1(w_q[293]), .A2(n7201), .ZN(n5383) );
  NAND2_X2 U4391 ( .A1(w_q[325]), .A2(n7259), .ZN(n5382) );
  NAND2_X2 U4392 ( .A1(n5384), .A2(n5385), .ZN(w_d[324]) );
  NAND2_X2 U4393 ( .A1(w_q[292]), .A2(n7201), .ZN(n5385) );
  NAND2_X2 U4394 ( .A1(w_q[324]), .A2(n7259), .ZN(n5384) );
  NAND2_X2 U4395 ( .A1(n5386), .A2(n5387), .ZN(w_d[323]) );
  NAND2_X2 U4396 ( .A1(w_q[291]), .A2(n7201), .ZN(n5387) );
  NAND2_X2 U4397 ( .A1(w_q[323]), .A2(n7259), .ZN(n5386) );
  NAND2_X2 U4398 ( .A1(n5388), .A2(n5389), .ZN(w_d[322]) );
  NAND2_X2 U4399 ( .A1(w_q[290]), .A2(n7201), .ZN(n5389) );
  NAND2_X2 U4400 ( .A1(w_q[322]), .A2(n7259), .ZN(n5388) );
  NAND2_X2 U4401 ( .A1(n5390), .A2(n5391), .ZN(w_d[321]) );
  NAND2_X2 U4402 ( .A1(w_q[289]), .A2(n7201), .ZN(n5391) );
  NAND2_X2 U4403 ( .A1(w_q[321]), .A2(n7259), .ZN(n5390) );
  NAND2_X2 U4404 ( .A1(n5392), .A2(n5393), .ZN(w_d[320]) );
  NAND2_X2 U4405 ( .A1(w_q[288]), .A2(n7201), .ZN(n5393) );
  NAND2_X2 U4406 ( .A1(w_q[320]), .A2(n7259), .ZN(n5392) );
  NAND2_X2 U4408 ( .A1(w[31]), .A2(n7159), .ZN(n5396) );
  NAND2_X2 U4409 ( .A1(w_q[31]), .A2(n7259), .ZN(n5395) );
  NAND2_X2 U4411 ( .A1(n5397), .A2(n5398), .ZN(w_d[319]) );
  NAND2_X2 U4412 ( .A1(w_q[287]), .A2(n7200), .ZN(n5398) );
  NAND2_X2 U4413 ( .A1(w_q[319]), .A2(n7259), .ZN(n5397) );
  NAND2_X2 U4414 ( .A1(n5399), .A2(n5400), .ZN(w_d[318]) );
  NAND2_X2 U4415 ( .A1(w_q[286]), .A2(n7200), .ZN(n5400) );
  NAND2_X2 U4416 ( .A1(w_q[318]), .A2(n7259), .ZN(n5399) );
  NAND2_X2 U4417 ( .A1(n5401), .A2(n5402), .ZN(w_d[317]) );
  NAND2_X2 U4418 ( .A1(w_q[285]), .A2(n7200), .ZN(n5402) );
  NAND2_X2 U4419 ( .A1(w_q[317]), .A2(n7258), .ZN(n5401) );
  NAND2_X2 U4420 ( .A1(n5403), .A2(n5404), .ZN(w_d[316]) );
  NAND2_X2 U4421 ( .A1(w_q[284]), .A2(n7200), .ZN(n5404) );
  NAND2_X2 U4422 ( .A1(w_q[316]), .A2(n7258), .ZN(n5403) );
  NAND2_X2 U4423 ( .A1(n5405), .A2(n5406), .ZN(w_d[315]) );
  NAND2_X2 U4424 ( .A1(w_q[283]), .A2(n7200), .ZN(n5406) );
  NAND2_X2 U4425 ( .A1(w_q[315]), .A2(n7258), .ZN(n5405) );
  NAND2_X2 U4426 ( .A1(n5407), .A2(n5408), .ZN(w_d[314]) );
  NAND2_X2 U4427 ( .A1(w_q[282]), .A2(n7200), .ZN(n5408) );
  NAND2_X2 U4428 ( .A1(w_q[314]), .A2(n7258), .ZN(n5407) );
  NAND2_X2 U4429 ( .A1(n5409), .A2(n5410), .ZN(w_d[313]) );
  NAND2_X2 U4430 ( .A1(w_q[281]), .A2(n7200), .ZN(n5410) );
  NAND2_X2 U4431 ( .A1(w_q[313]), .A2(n7258), .ZN(n5409) );
  NAND2_X2 U4432 ( .A1(n5411), .A2(n5412), .ZN(w_d[312]) );
  NAND2_X2 U4433 ( .A1(w_q[280]), .A2(n7200), .ZN(n5412) );
  NAND2_X2 U4434 ( .A1(w_q[312]), .A2(n7258), .ZN(n5411) );
  NAND2_X2 U4435 ( .A1(n5413), .A2(n5414), .ZN(w_d[311]) );
  NAND2_X2 U4436 ( .A1(w_q[279]), .A2(n7200), .ZN(n5414) );
  NAND2_X2 U4437 ( .A1(w_q[311]), .A2(n7258), .ZN(n5413) );
  NAND2_X2 U4438 ( .A1(n5415), .A2(n5416), .ZN(w_d[310]) );
  NAND2_X2 U4439 ( .A1(w_q[278]), .A2(n7200), .ZN(n5416) );
  NAND2_X2 U4440 ( .A1(w_q[310]), .A2(n7258), .ZN(n5415) );
  NAND2_X2 U4442 ( .A1(w[30]), .A2(n7159), .ZN(n5419) );
  NAND2_X2 U4443 ( .A1(w_q[30]), .A2(n7258), .ZN(n5418) );
  NAND2_X2 U4445 ( .A1(n5420), .A2(n5421), .ZN(w_d[309]) );
  NAND2_X2 U4446 ( .A1(w_q[277]), .A2(n7200), .ZN(n5421) );
  NAND2_X2 U4447 ( .A1(w_q[309]), .A2(n7258), .ZN(n5420) );
  NAND2_X2 U4448 ( .A1(n5422), .A2(n5423), .ZN(w_d[308]) );
  NAND2_X2 U4449 ( .A1(w_q[276]), .A2(n7199), .ZN(n5423) );
  NAND2_X2 U4450 ( .A1(w_q[308]), .A2(n7258), .ZN(n5422) );
  NAND2_X2 U4451 ( .A1(n5424), .A2(n5425), .ZN(w_d[307]) );
  NAND2_X2 U4452 ( .A1(w_q[275]), .A2(n7199), .ZN(n5425) );
  NAND2_X2 U4453 ( .A1(w_q[307]), .A2(n7257), .ZN(n5424) );
  NAND2_X2 U4454 ( .A1(n5426), .A2(n5427), .ZN(w_d[306]) );
  NAND2_X2 U4455 ( .A1(w_q[274]), .A2(n7199), .ZN(n5427) );
  NAND2_X2 U4456 ( .A1(w_q[306]), .A2(n7257), .ZN(n5426) );
  NAND2_X2 U4457 ( .A1(n5428), .A2(n5429), .ZN(w_d[305]) );
  NAND2_X2 U4458 ( .A1(w_q[273]), .A2(n7199), .ZN(n5429) );
  NAND2_X2 U4459 ( .A1(w_q[305]), .A2(n7257), .ZN(n5428) );
  NAND2_X2 U4460 ( .A1(n5430), .A2(n5431), .ZN(w_d[304]) );
  NAND2_X2 U4461 ( .A1(w_q[272]), .A2(n7199), .ZN(n5431) );
  NAND2_X2 U4462 ( .A1(w_q[304]), .A2(n7257), .ZN(n5430) );
  NAND2_X2 U4463 ( .A1(n5432), .A2(n5433), .ZN(w_d[303]) );
  NAND2_X2 U4464 ( .A1(w_q[271]), .A2(n7199), .ZN(n5433) );
  NAND2_X2 U4465 ( .A1(w_q[303]), .A2(n7257), .ZN(n5432) );
  NAND2_X2 U4466 ( .A1(n5434), .A2(n5435), .ZN(w_d[302]) );
  NAND2_X2 U4467 ( .A1(w_q[270]), .A2(n7199), .ZN(n5435) );
  NAND2_X2 U4468 ( .A1(w_q[302]), .A2(n7257), .ZN(n5434) );
  NAND2_X2 U4469 ( .A1(n5436), .A2(n5437), .ZN(w_d[301]) );
  NAND2_X2 U4470 ( .A1(w_q[269]), .A2(n7199), .ZN(n5437) );
  NAND2_X2 U4471 ( .A1(w_q[301]), .A2(n7257), .ZN(n5436) );
  NAND2_X2 U4472 ( .A1(n5438), .A2(n5439), .ZN(w_d[300]) );
  NAND2_X2 U4473 ( .A1(w_q[268]), .A2(n7199), .ZN(n5439) );
  NAND2_X2 U4474 ( .A1(w_q[300]), .A2(n7257), .ZN(n5438) );
  NAND2_X2 U4476 ( .A1(w[2]), .A2(n7159), .ZN(n5442) );
  NAND2_X2 U4477 ( .A1(w_q[2]), .A2(n7257), .ZN(n5441) );
  NAND2_X2 U4480 ( .A1(w[29]), .A2(n7159), .ZN(n5445) );
  NAND2_X2 U4481 ( .A1(w_q[29]), .A2(n7257), .ZN(n5444) );
  NAND2_X2 U4483 ( .A1(n5446), .A2(n5447), .ZN(w_d[299]) );
  NAND2_X2 U4484 ( .A1(w_q[267]), .A2(n7199), .ZN(n5447) );
  NAND2_X2 U4485 ( .A1(w_q[299]), .A2(n7257), .ZN(n5446) );
  NAND2_X2 U4486 ( .A1(n5448), .A2(n5449), .ZN(w_d[298]) );
  NAND2_X2 U4487 ( .A1(w_q[266]), .A2(n7199), .ZN(n5449) );
  NAND2_X2 U4488 ( .A1(w_q[298]), .A2(n7256), .ZN(n5448) );
  NAND2_X2 U4489 ( .A1(n5450), .A2(n5451), .ZN(w_d[297]) );
  NAND2_X2 U4490 ( .A1(w_q[265]), .A2(n7198), .ZN(n5451) );
  NAND2_X2 U4491 ( .A1(w_q[297]), .A2(n7256), .ZN(n5450) );
  NAND2_X2 U4492 ( .A1(n5452), .A2(n5453), .ZN(w_d[296]) );
  NAND2_X2 U4493 ( .A1(w_q[264]), .A2(n7198), .ZN(n5453) );
  NAND2_X2 U4494 ( .A1(w_q[296]), .A2(n7256), .ZN(n5452) );
  NAND2_X2 U4495 ( .A1(n5454), .A2(n5455), .ZN(w_d[295]) );
  NAND2_X2 U4496 ( .A1(w_q[263]), .A2(n7198), .ZN(n5455) );
  NAND2_X2 U4497 ( .A1(w_q[295]), .A2(n7256), .ZN(n5454) );
  NAND2_X2 U4498 ( .A1(n5456), .A2(n5457), .ZN(w_d[294]) );
  NAND2_X2 U4499 ( .A1(w_q[262]), .A2(n7198), .ZN(n5457) );
  NAND2_X2 U4500 ( .A1(w_q[294]), .A2(n7256), .ZN(n5456) );
  NAND2_X2 U4501 ( .A1(n5458), .A2(n5459), .ZN(w_d[293]) );
  NAND2_X2 U4502 ( .A1(w_q[261]), .A2(n7198), .ZN(n5459) );
  NAND2_X2 U4503 ( .A1(w_q[293]), .A2(n7256), .ZN(n5458) );
  NAND2_X2 U4504 ( .A1(n5460), .A2(n5461), .ZN(w_d[292]) );
  NAND2_X2 U4505 ( .A1(w_q[260]), .A2(n7198), .ZN(n5461) );
  NAND2_X2 U4506 ( .A1(w_q[292]), .A2(n7256), .ZN(n5460) );
  NAND2_X2 U4507 ( .A1(n5462), .A2(n5463), .ZN(w_d[291]) );
  NAND2_X2 U4508 ( .A1(w_q[259]), .A2(n7198), .ZN(n5463) );
  NAND2_X2 U4509 ( .A1(w_q[291]), .A2(n7256), .ZN(n5462) );
  NAND2_X2 U4510 ( .A1(n5464), .A2(n5465), .ZN(w_d[290]) );
  NAND2_X2 U4511 ( .A1(w_q[258]), .A2(n7198), .ZN(n5465) );
  NAND2_X2 U4512 ( .A1(w_q[290]), .A2(n7256), .ZN(n5464) );
  NAND2_X2 U4514 ( .A1(w[28]), .A2(n7159), .ZN(n5468) );
  NAND2_X2 U4515 ( .A1(w_q[28]), .A2(n7256), .ZN(n5467) );
  NAND2_X2 U4517 ( .A1(n5469), .A2(n5470), .ZN(w_d[289]) );
  NAND2_X2 U4518 ( .A1(w_q[257]), .A2(n7198), .ZN(n5470) );
  NAND2_X2 U4519 ( .A1(w_q[289]), .A2(n7256), .ZN(n5469) );
  NAND2_X2 U4520 ( .A1(n5471), .A2(n5472), .ZN(w_d[288]) );
  NAND2_X2 U4521 ( .A1(w_q[256]), .A2(n7198), .ZN(n5472) );
  NAND2_X2 U4522 ( .A1(w_q[288]), .A2(n7255), .ZN(n5471) );
  NAND2_X2 U4523 ( .A1(n5473), .A2(n5474), .ZN(w_d[287]) );
  NAND2_X2 U4524 ( .A1(w_q[255]), .A2(n7198), .ZN(n5474) );
  NAND2_X2 U4525 ( .A1(w_q[287]), .A2(n7255), .ZN(n5473) );
  NAND2_X2 U4526 ( .A1(n5475), .A2(n5476), .ZN(w_d[286]) );
  NAND2_X2 U4527 ( .A1(w_q[254]), .A2(n7197), .ZN(n5476) );
  NAND2_X2 U4528 ( .A1(w_q[286]), .A2(n7255), .ZN(n5475) );
  NAND2_X2 U4529 ( .A1(n5477), .A2(n5478), .ZN(w_d[285]) );
  NAND2_X2 U4530 ( .A1(w_q[253]), .A2(n7197), .ZN(n5478) );
  NAND2_X2 U4531 ( .A1(w_q[285]), .A2(n7255), .ZN(n5477) );
  NAND2_X2 U4532 ( .A1(n5479), .A2(n5480), .ZN(w_d[284]) );
  NAND2_X2 U4533 ( .A1(w_q[252]), .A2(n7197), .ZN(n5480) );
  NAND2_X2 U4534 ( .A1(w_q[284]), .A2(n7255), .ZN(n5479) );
  NAND2_X2 U4535 ( .A1(n5481), .A2(n5482), .ZN(w_d[283]) );
  NAND2_X2 U4536 ( .A1(w_q[251]), .A2(n7197), .ZN(n5482) );
  NAND2_X2 U4537 ( .A1(w_q[283]), .A2(n7255), .ZN(n5481) );
  NAND2_X2 U4538 ( .A1(n5483), .A2(n5484), .ZN(w_d[282]) );
  NAND2_X2 U4539 ( .A1(w_q[250]), .A2(n7197), .ZN(n5484) );
  NAND2_X2 U4540 ( .A1(w_q[282]), .A2(n7255), .ZN(n5483) );
  NAND2_X2 U4541 ( .A1(n5485), .A2(n5486), .ZN(w_d[281]) );
  NAND2_X2 U4542 ( .A1(w_q[249]), .A2(n7197), .ZN(n5486) );
  NAND2_X2 U4543 ( .A1(w_q[281]), .A2(n7255), .ZN(n5485) );
  NAND2_X2 U4544 ( .A1(n5487), .A2(n5488), .ZN(w_d[280]) );
  NAND2_X2 U4545 ( .A1(w_q[248]), .A2(n7197), .ZN(n5488) );
  NAND2_X2 U4546 ( .A1(w_q[280]), .A2(n7255), .ZN(n5487) );
  NAND2_X2 U4548 ( .A1(w[27]), .A2(n7159), .ZN(n5491) );
  NAND2_X2 U4549 ( .A1(w_q[27]), .A2(n7255), .ZN(n5490) );
  NAND2_X2 U4551 ( .A1(n5492), .A2(n5493), .ZN(w_d[279]) );
  NAND2_X2 U4552 ( .A1(w_q[247]), .A2(n7197), .ZN(n5493) );
  NAND2_X2 U4553 ( .A1(w_q[279]), .A2(n7255), .ZN(n5492) );
  NAND2_X2 U4554 ( .A1(n5494), .A2(n5495), .ZN(w_d[278]) );
  NAND2_X2 U4555 ( .A1(w_q[246]), .A2(n7197), .ZN(n5495) );
  NAND2_X2 U4556 ( .A1(w_q[278]), .A2(n7254), .ZN(n5494) );
  NAND2_X2 U4557 ( .A1(n5496), .A2(n5497), .ZN(w_d[277]) );
  NAND2_X2 U4558 ( .A1(w_q[245]), .A2(n7197), .ZN(n5497) );
  NAND2_X2 U4559 ( .A1(w_q[277]), .A2(n7254), .ZN(n5496) );
  NAND2_X2 U4560 ( .A1(n5498), .A2(n5499), .ZN(w_d[276]) );
  NAND2_X2 U4561 ( .A1(w_q[244]), .A2(n7197), .ZN(n5499) );
  NAND2_X2 U4562 ( .A1(w_q[276]), .A2(n7254), .ZN(n5498) );
  NAND2_X2 U4563 ( .A1(n5500), .A2(n5501), .ZN(w_d[275]) );
  NAND2_X2 U4564 ( .A1(w_q[243]), .A2(n7196), .ZN(n5501) );
  NAND2_X2 U4565 ( .A1(w_q[275]), .A2(n7254), .ZN(n5500) );
  NAND2_X2 U4566 ( .A1(n5502), .A2(n5503), .ZN(w_d[274]) );
  NAND2_X2 U4567 ( .A1(w_q[242]), .A2(n7196), .ZN(n5503) );
  NAND2_X2 U4568 ( .A1(w_q[274]), .A2(n7254), .ZN(n5502) );
  NAND2_X2 U4569 ( .A1(n5504), .A2(n5505), .ZN(w_d[273]) );
  NAND2_X2 U4570 ( .A1(w_q[241]), .A2(n7196), .ZN(n5505) );
  NAND2_X2 U4571 ( .A1(w_q[273]), .A2(n7254), .ZN(n5504) );
  NAND2_X2 U4572 ( .A1(n5506), .A2(n5507), .ZN(w_d[272]) );
  NAND2_X2 U4573 ( .A1(w_q[240]), .A2(n7196), .ZN(n5507) );
  NAND2_X2 U4574 ( .A1(w_q[272]), .A2(n7254), .ZN(n5506) );
  NAND2_X2 U4575 ( .A1(n5508), .A2(n5509), .ZN(w_d[271]) );
  NAND2_X2 U4576 ( .A1(w_q[239]), .A2(n7196), .ZN(n5509) );
  NAND2_X2 U4577 ( .A1(w_q[271]), .A2(n7254), .ZN(n5508) );
  NAND2_X2 U4578 ( .A1(n5510), .A2(n5511), .ZN(w_d[270]) );
  NAND2_X2 U4579 ( .A1(w_q[238]), .A2(n7196), .ZN(n5511) );
  NAND2_X2 U4580 ( .A1(w_q[270]), .A2(n7254), .ZN(n5510) );
  NAND2_X2 U4582 ( .A1(w[26]), .A2(n7160), .ZN(n5514) );
  NAND2_X2 U4583 ( .A1(w_q[26]), .A2(n7254), .ZN(n5513) );
  NAND2_X2 U4585 ( .A1(n5515), .A2(n5516), .ZN(w_d[269]) );
  NAND2_X2 U4586 ( .A1(w_q[237]), .A2(n7196), .ZN(n5516) );
  NAND2_X2 U4587 ( .A1(w_q[269]), .A2(n7254), .ZN(n5515) );
  NAND2_X2 U4588 ( .A1(n5517), .A2(n5518), .ZN(w_d[268]) );
  NAND2_X2 U4589 ( .A1(w_q[236]), .A2(n7196), .ZN(n5518) );
  NAND2_X2 U4590 ( .A1(w_q[268]), .A2(n7253), .ZN(n5517) );
  NAND2_X2 U4591 ( .A1(n5519), .A2(n5520), .ZN(w_d[267]) );
  NAND2_X2 U4592 ( .A1(w_q[235]), .A2(n7196), .ZN(n5520) );
  NAND2_X2 U4593 ( .A1(w_q[267]), .A2(n7253), .ZN(n5519) );
  NAND2_X2 U4594 ( .A1(n5521), .A2(n5522), .ZN(w_d[266]) );
  NAND2_X2 U4595 ( .A1(w_q[234]), .A2(n7196), .ZN(n5522) );
  NAND2_X2 U4596 ( .A1(w_q[266]), .A2(n7253), .ZN(n5521) );
  NAND2_X2 U4597 ( .A1(n5523), .A2(n5524), .ZN(w_d[265]) );
  NAND2_X2 U4598 ( .A1(w_q[233]), .A2(n7196), .ZN(n5524) );
  NAND2_X2 U4599 ( .A1(w_q[265]), .A2(n7253), .ZN(n5523) );
  NAND2_X2 U4600 ( .A1(n5525), .A2(n5526), .ZN(w_d[264]) );
  NAND2_X2 U4601 ( .A1(w_q[232]), .A2(n7195), .ZN(n5526) );
  NAND2_X2 U4602 ( .A1(w_q[264]), .A2(n7253), .ZN(n5525) );
  NAND2_X2 U4603 ( .A1(n5527), .A2(n5528), .ZN(w_d[263]) );
  NAND2_X2 U4604 ( .A1(w_q[231]), .A2(n7195), .ZN(n5528) );
  NAND2_X2 U4605 ( .A1(w_q[263]), .A2(n7253), .ZN(n5527) );
  NAND2_X2 U4606 ( .A1(n5529), .A2(n5530), .ZN(w_d[262]) );
  NAND2_X2 U4607 ( .A1(w_q[230]), .A2(n7195), .ZN(n5530) );
  NAND2_X2 U4608 ( .A1(w_q[262]), .A2(n7253), .ZN(n5529) );
  NAND2_X2 U4609 ( .A1(n5531), .A2(n5532), .ZN(w_d[261]) );
  NAND2_X2 U4610 ( .A1(w_q[229]), .A2(n7195), .ZN(n5532) );
  NAND2_X2 U4611 ( .A1(w_q[261]), .A2(n7253), .ZN(n5531) );
  NAND2_X2 U4612 ( .A1(n5533), .A2(n5534), .ZN(w_d[260]) );
  NAND2_X2 U4613 ( .A1(w_q[228]), .A2(n7195), .ZN(n5534) );
  NAND2_X2 U4614 ( .A1(w_q[260]), .A2(n7253), .ZN(n5533) );
  NAND2_X2 U4616 ( .A1(w[25]), .A2(n7160), .ZN(n5537) );
  NAND2_X2 U4617 ( .A1(w_q[25]), .A2(n7253), .ZN(n5536) );
  NAND2_X2 U4619 ( .A1(n5538), .A2(n5539), .ZN(w_d[259]) );
  NAND2_X2 U4620 ( .A1(w_q[227]), .A2(n7195), .ZN(n5539) );
  NAND2_X2 U4621 ( .A1(w_q[259]), .A2(n7253), .ZN(n5538) );
  NAND2_X2 U4622 ( .A1(n5540), .A2(n5541), .ZN(w_d[258]) );
  NAND2_X2 U4623 ( .A1(w_q[226]), .A2(n7195), .ZN(n5541) );
  NAND2_X2 U4624 ( .A1(w_q[258]), .A2(n7252), .ZN(n5540) );
  NAND2_X2 U4625 ( .A1(n5542), .A2(n5543), .ZN(w_d[257]) );
  NAND2_X2 U4626 ( .A1(w_q[225]), .A2(n7195), .ZN(n5543) );
  NAND2_X2 U4627 ( .A1(w_q[257]), .A2(n7252), .ZN(n5542) );
  NAND2_X2 U4628 ( .A1(n5544), .A2(n5545), .ZN(w_d[256]) );
  NAND2_X2 U4629 ( .A1(w_q[224]), .A2(n7195), .ZN(n5545) );
  NAND2_X2 U4630 ( .A1(w_q[256]), .A2(n7252), .ZN(n5544) );
  NAND2_X2 U4631 ( .A1(n5546), .A2(n5547), .ZN(w_d[255]) );
  NAND2_X2 U4632 ( .A1(w_q[223]), .A2(n7195), .ZN(n5547) );
  NAND2_X2 U4633 ( .A1(w_q[255]), .A2(n7252), .ZN(n5546) );
  NAND2_X2 U4634 ( .A1(n5548), .A2(n5549), .ZN(w_d[254]) );
  NAND2_X2 U4635 ( .A1(w_q[222]), .A2(n7195), .ZN(n5549) );
  NAND2_X2 U4636 ( .A1(w_q[254]), .A2(n7252), .ZN(n5548) );
  NAND2_X2 U4637 ( .A1(n5550), .A2(n5551), .ZN(w_d[253]) );
  NAND2_X2 U4638 ( .A1(w_q[221]), .A2(n7194), .ZN(n5551) );
  NAND2_X2 U4639 ( .A1(w_q[253]), .A2(n7252), .ZN(n5550) );
  NAND2_X2 U4640 ( .A1(n5552), .A2(n5553), .ZN(w_d[252]) );
  NAND2_X2 U4641 ( .A1(w_q[220]), .A2(n7194), .ZN(n5553) );
  NAND2_X2 U4642 ( .A1(w_q[252]), .A2(n7252), .ZN(n5552) );
  NAND2_X2 U4643 ( .A1(n5554), .A2(n5555), .ZN(w_d[251]) );
  NAND2_X2 U4644 ( .A1(w_q[219]), .A2(n7194), .ZN(n5555) );
  NAND2_X2 U4645 ( .A1(w_q[251]), .A2(n7252), .ZN(n5554) );
  NAND2_X2 U4646 ( .A1(n5556), .A2(n5557), .ZN(w_d[250]) );
  NAND2_X2 U4647 ( .A1(w_q[218]), .A2(n7194), .ZN(n5557) );
  NAND2_X2 U4648 ( .A1(w_q[250]), .A2(n7252), .ZN(n5556) );
  NAND2_X2 U4650 ( .A1(w[24]), .A2(n7160), .ZN(n5560) );
  NAND2_X2 U4651 ( .A1(w_q[24]), .A2(n7252), .ZN(n5559) );
  NAND2_X2 U4653 ( .A1(n5561), .A2(n5562), .ZN(w_d[249]) );
  NAND2_X2 U4654 ( .A1(w_q[217]), .A2(n7194), .ZN(n5562) );
  NAND2_X2 U4655 ( .A1(w_q[249]), .A2(n7252), .ZN(n5561) );
  NAND2_X2 U4656 ( .A1(n5563), .A2(n5564), .ZN(w_d[248]) );
  NAND2_X2 U4657 ( .A1(w_q[216]), .A2(n7194), .ZN(n5564) );
  NAND2_X2 U4658 ( .A1(w_q[248]), .A2(n7234), .ZN(n5563) );
  NAND2_X2 U4659 ( .A1(n5565), .A2(n5566), .ZN(w_d[247]) );
  NAND2_X2 U4660 ( .A1(w_q[215]), .A2(n7194), .ZN(n5566) );
  NAND2_X2 U4661 ( .A1(w_q[247]), .A2(n7233), .ZN(n5565) );
  NAND2_X2 U4662 ( .A1(n5567), .A2(n5568), .ZN(w_d[246]) );
  NAND2_X2 U4663 ( .A1(w_q[214]), .A2(n7194), .ZN(n5568) );
  NAND2_X2 U4664 ( .A1(w_q[246]), .A2(n7235), .ZN(n5567) );
  NAND2_X2 U4665 ( .A1(n5569), .A2(n5570), .ZN(w_d[245]) );
  NAND2_X2 U4666 ( .A1(w_q[213]), .A2(n7194), .ZN(n5570) );
  NAND2_X2 U4667 ( .A1(w_q[245]), .A2(n7236), .ZN(n5569) );
  NAND2_X2 U4668 ( .A1(n5571), .A2(n5572), .ZN(w_d[244]) );
  NAND2_X2 U4669 ( .A1(w_q[212]), .A2(n7194), .ZN(n5572) );
  NAND2_X2 U4670 ( .A1(w_q[244]), .A2(n7231), .ZN(n5571) );
  NAND2_X2 U4671 ( .A1(n5573), .A2(n5574), .ZN(w_d[243]) );
  NAND2_X2 U4672 ( .A1(w_q[211]), .A2(n7194), .ZN(n5574) );
  NAND2_X2 U4673 ( .A1(w_q[243]), .A2(n7234), .ZN(n5573) );
  NAND2_X2 U4674 ( .A1(n5575), .A2(n5576), .ZN(w_d[242]) );
  NAND2_X2 U4675 ( .A1(w_q[210]), .A2(n7193), .ZN(n5576) );
  NAND2_X2 U4676 ( .A1(w_q[242]), .A2(n7233), .ZN(n5575) );
  NAND2_X2 U4677 ( .A1(n5577), .A2(n5578), .ZN(w_d[241]) );
  NAND2_X2 U4678 ( .A1(w_q[209]), .A2(n7193), .ZN(n5578) );
  NAND2_X2 U4679 ( .A1(w_q[241]), .A2(n7232), .ZN(n5577) );
  NAND2_X2 U4680 ( .A1(n5579), .A2(n5580), .ZN(w_d[240]) );
  NAND2_X2 U4681 ( .A1(w_q[208]), .A2(n7193), .ZN(n5580) );
  NAND2_X2 U4682 ( .A1(w_q[240]), .A2(n7230), .ZN(n5579) );
  NAND2_X2 U4684 ( .A1(w[23]), .A2(n7160), .ZN(n5583) );
  NAND2_X2 U4685 ( .A1(w_q[23]), .A2(n7274), .ZN(n5582) );
  NAND2_X2 U4687 ( .A1(n5584), .A2(n5585), .ZN(w_d[239]) );
  NAND2_X2 U4688 ( .A1(w_q[207]), .A2(n7193), .ZN(n5585) );
  NAND2_X2 U4689 ( .A1(w_q[239]), .A2(n7231), .ZN(n5584) );
  NAND2_X2 U4690 ( .A1(n5586), .A2(n5587), .ZN(w_d[238]) );
  NAND2_X2 U4691 ( .A1(w_q[206]), .A2(n7193), .ZN(n5587) );
  NAND2_X2 U4692 ( .A1(w_q[238]), .A2(n7232), .ZN(n5586) );
  NAND2_X2 U4693 ( .A1(n5588), .A2(n5589), .ZN(w_d[237]) );
  NAND2_X2 U4694 ( .A1(w_q[205]), .A2(n7193), .ZN(n5589) );
  NAND2_X2 U4695 ( .A1(w_q[237]), .A2(n7230), .ZN(n5588) );
  NAND2_X2 U4696 ( .A1(n5590), .A2(n5591), .ZN(w_d[236]) );
  NAND2_X2 U4697 ( .A1(w_q[204]), .A2(n7193), .ZN(n5591) );
  NAND2_X2 U4698 ( .A1(w_q[236]), .A2(n7238), .ZN(n5590) );
  NAND2_X2 U4699 ( .A1(n5592), .A2(n5593), .ZN(w_d[235]) );
  NAND2_X2 U4700 ( .A1(w_q[203]), .A2(n7193), .ZN(n5593) );
  NAND2_X2 U4701 ( .A1(w_q[235]), .A2(n7231), .ZN(n5592) );
  NAND2_X2 U4702 ( .A1(n5594), .A2(n5595), .ZN(w_d[234]) );
  NAND2_X2 U4703 ( .A1(w_q[202]), .A2(n7193), .ZN(n5595) );
  NAND2_X2 U4704 ( .A1(w_q[234]), .A2(n7233), .ZN(n5594) );
  NAND2_X2 U4705 ( .A1(n5596), .A2(n5597), .ZN(w_d[233]) );
  NAND2_X2 U4706 ( .A1(w_q[201]), .A2(n7193), .ZN(n5597) );
  NAND2_X2 U4707 ( .A1(w_q[233]), .A2(n7235), .ZN(n5596) );
  NAND2_X2 U4708 ( .A1(n5598), .A2(n5599), .ZN(w_d[232]) );
  NAND2_X2 U4709 ( .A1(w_q[200]), .A2(n7193), .ZN(n5599) );
  NAND2_X2 U4710 ( .A1(w_q[232]), .A2(n7232), .ZN(n5598) );
  NAND2_X2 U4711 ( .A1(n5600), .A2(n5601), .ZN(w_d[231]) );
  NAND2_X2 U4712 ( .A1(w_q[199]), .A2(n7192), .ZN(n5601) );
  NAND2_X2 U4713 ( .A1(w_q[231]), .A2(n7230), .ZN(n5600) );
  NAND2_X2 U4714 ( .A1(n5602), .A2(n5603), .ZN(w_d[230]) );
  NAND2_X2 U4715 ( .A1(w_q[198]), .A2(n7192), .ZN(n5603) );
  NAND2_X2 U4716 ( .A1(w_q[230]), .A2(n7234), .ZN(n5602) );
  NAND2_X2 U4718 ( .A1(w[22]), .A2(n7160), .ZN(n5606) );
  NAND2_X2 U4719 ( .A1(w_q[22]), .A2(n7267), .ZN(n5605) );
  NAND2_X2 U4721 ( .A1(n5607), .A2(n5608), .ZN(w_d[229]) );
  NAND2_X2 U4722 ( .A1(w_q[197]), .A2(n7192), .ZN(n5608) );
  NAND2_X2 U4723 ( .A1(w_q[229]), .A2(n7238), .ZN(n5607) );
  NAND2_X2 U4724 ( .A1(n5609), .A2(n5610), .ZN(w_d[228]) );
  NAND2_X2 U4725 ( .A1(w_q[196]), .A2(n7192), .ZN(n5610) );
  NAND2_X2 U4726 ( .A1(w_q[228]), .A2(n7251), .ZN(n5609) );
  NAND2_X2 U4727 ( .A1(n5611), .A2(n5612), .ZN(w_d[227]) );
  NAND2_X2 U4728 ( .A1(w_q[195]), .A2(n7192), .ZN(n5612) );
  NAND2_X2 U4729 ( .A1(w_q[227]), .A2(n7251), .ZN(n5611) );
  NAND2_X2 U4730 ( .A1(n5613), .A2(n5614), .ZN(w_d[226]) );
  NAND2_X2 U4731 ( .A1(w_q[194]), .A2(n7192), .ZN(n5614) );
  NAND2_X2 U4732 ( .A1(w_q[226]), .A2(n7251), .ZN(n5613) );
  NAND2_X2 U4733 ( .A1(n5615), .A2(n5616), .ZN(w_d[225]) );
  NAND2_X2 U4734 ( .A1(w_q[193]), .A2(n7192), .ZN(n5616) );
  NAND2_X2 U4735 ( .A1(w_q[225]), .A2(n7251), .ZN(n5615) );
  NAND2_X2 U4736 ( .A1(n5617), .A2(n5618), .ZN(w_d[224]) );
  NAND2_X2 U4737 ( .A1(w_q[192]), .A2(n7192), .ZN(n5618) );
  NAND2_X2 U4738 ( .A1(w_q[224]), .A2(n7251), .ZN(n5617) );
  NAND2_X2 U4739 ( .A1(n5619), .A2(n5620), .ZN(w_d[223]) );
  NAND2_X2 U4740 ( .A1(w_q[191]), .A2(n7192), .ZN(n5620) );
  NAND2_X2 U4741 ( .A1(w_q[223]), .A2(n7251), .ZN(n5619) );
  NAND2_X2 U4742 ( .A1(n5621), .A2(n5622), .ZN(w_d[222]) );
  NAND2_X2 U4743 ( .A1(w_q[190]), .A2(n7192), .ZN(n5622) );
  NAND2_X2 U4744 ( .A1(w_q[222]), .A2(n7251), .ZN(n5621) );
  NAND2_X2 U4745 ( .A1(n5623), .A2(n5624), .ZN(w_d[221]) );
  NAND2_X2 U4746 ( .A1(w_q[189]), .A2(n7192), .ZN(n5624) );
  NAND2_X2 U4747 ( .A1(w_q[221]), .A2(n7251), .ZN(n5623) );
  NAND2_X2 U4748 ( .A1(n5625), .A2(n5626), .ZN(w_d[220]) );
  NAND2_X2 U4749 ( .A1(w_q[188]), .A2(n7191), .ZN(n5626) );
  NAND2_X2 U4750 ( .A1(w_q[220]), .A2(n7251), .ZN(n5625) );
  NAND2_X2 U4752 ( .A1(w[21]), .A2(n7160), .ZN(n5629) );
  NAND2_X2 U4753 ( .A1(w_q[21]), .A2(n7251), .ZN(n5628) );
  NAND2_X2 U4755 ( .A1(n5630), .A2(n5631), .ZN(w_d[219]) );
  NAND2_X2 U4756 ( .A1(w_q[187]), .A2(n7191), .ZN(n5631) );
  NAND2_X2 U4757 ( .A1(w_q[219]), .A2(n7251), .ZN(n5630) );
  NAND2_X2 U4758 ( .A1(n5632), .A2(n5633), .ZN(w_d[218]) );
  NAND2_X2 U4759 ( .A1(w_q[186]), .A2(n7191), .ZN(n5633) );
  NAND2_X2 U4760 ( .A1(w_q[218]), .A2(n7250), .ZN(n5632) );
  NAND2_X2 U4761 ( .A1(n5634), .A2(n5635), .ZN(w_d[217]) );
  NAND2_X2 U4762 ( .A1(w_q[185]), .A2(n7191), .ZN(n5635) );
  NAND2_X2 U4763 ( .A1(w_q[217]), .A2(n7250), .ZN(n5634) );
  NAND2_X2 U4764 ( .A1(n5636), .A2(n5637), .ZN(w_d[216]) );
  NAND2_X2 U4765 ( .A1(w_q[184]), .A2(n7191), .ZN(n5637) );
  NAND2_X2 U4766 ( .A1(w_q[216]), .A2(n7250), .ZN(n5636) );
  NAND2_X2 U4767 ( .A1(n5638), .A2(n5639), .ZN(w_d[215]) );
  NAND2_X2 U4768 ( .A1(w_q[183]), .A2(n7191), .ZN(n5639) );
  NAND2_X2 U4769 ( .A1(w_q[215]), .A2(n7250), .ZN(n5638) );
  NAND2_X2 U4770 ( .A1(n5640), .A2(n5641), .ZN(w_d[214]) );
  NAND2_X2 U4771 ( .A1(w_q[182]), .A2(n7191), .ZN(n5641) );
  NAND2_X2 U4772 ( .A1(w_q[214]), .A2(n7250), .ZN(n5640) );
  NAND2_X2 U4773 ( .A1(n5642), .A2(n5643), .ZN(w_d[213]) );
  NAND2_X2 U4774 ( .A1(w_q[181]), .A2(n7191), .ZN(n5643) );
  NAND2_X2 U4775 ( .A1(w_q[213]), .A2(n7250), .ZN(n5642) );
  NAND2_X2 U4776 ( .A1(n5644), .A2(n5645), .ZN(w_d[212]) );
  NAND2_X2 U4777 ( .A1(w_q[180]), .A2(n7191), .ZN(n5645) );
  NAND2_X2 U4778 ( .A1(w_q[212]), .A2(n7250), .ZN(n5644) );
  NAND2_X2 U4779 ( .A1(n5646), .A2(n5647), .ZN(w_d[211]) );
  NAND2_X2 U4780 ( .A1(w_q[179]), .A2(n7191), .ZN(n5647) );
  NAND2_X2 U4781 ( .A1(w_q[211]), .A2(n7250), .ZN(n5646) );
  NAND2_X2 U4782 ( .A1(n5648), .A2(n5649), .ZN(w_d[210]) );
  NAND2_X2 U4783 ( .A1(w_q[178]), .A2(n7191), .ZN(n5649) );
  NAND2_X2 U4784 ( .A1(w_q[210]), .A2(n7250), .ZN(n5648) );
  NAND2_X2 U4786 ( .A1(w[20]), .A2(n7160), .ZN(n5652) );
  NAND2_X2 U4787 ( .A1(w_q[20]), .A2(n7250), .ZN(n5651) );
  NAND2_X2 U4789 ( .A1(n5653), .A2(n5654), .ZN(w_d[209]) );
  NAND2_X2 U4790 ( .A1(w_q[177]), .A2(n7190), .ZN(n5654) );
  NAND2_X2 U4791 ( .A1(w_q[209]), .A2(n7250), .ZN(n5653) );
  NAND2_X2 U4792 ( .A1(n5655), .A2(n5656), .ZN(w_d[208]) );
  NAND2_X2 U4793 ( .A1(w_q[176]), .A2(n7190), .ZN(n5656) );
  NAND2_X2 U4794 ( .A1(w_q[208]), .A2(n7249), .ZN(n5655) );
  NAND2_X2 U4795 ( .A1(n5657), .A2(n5658), .ZN(w_d[207]) );
  NAND2_X2 U4796 ( .A1(w_q[175]), .A2(n7190), .ZN(n5658) );
  NAND2_X2 U4797 ( .A1(w_q[207]), .A2(n7249), .ZN(n5657) );
  NAND2_X2 U4798 ( .A1(n5659), .A2(n5660), .ZN(w_d[206]) );
  NAND2_X2 U4799 ( .A1(w_q[174]), .A2(n7190), .ZN(n5660) );
  NAND2_X2 U4800 ( .A1(w_q[206]), .A2(n7249), .ZN(n5659) );
  NAND2_X2 U4801 ( .A1(n5661), .A2(n5662), .ZN(w_d[205]) );
  NAND2_X2 U4802 ( .A1(w_q[173]), .A2(n7190), .ZN(n5662) );
  NAND2_X2 U4803 ( .A1(w_q[205]), .A2(n7249), .ZN(n5661) );
  NAND2_X2 U4804 ( .A1(n5663), .A2(n5664), .ZN(w_d[204]) );
  NAND2_X2 U4805 ( .A1(w_q[172]), .A2(n7190), .ZN(n5664) );
  NAND2_X2 U4806 ( .A1(w_q[204]), .A2(n7249), .ZN(n5663) );
  NAND2_X2 U4807 ( .A1(n5665), .A2(n5666), .ZN(w_d[203]) );
  NAND2_X2 U4808 ( .A1(w_q[171]), .A2(n7190), .ZN(n5666) );
  NAND2_X2 U4809 ( .A1(w_q[203]), .A2(n7249), .ZN(n5665) );
  NAND2_X2 U4810 ( .A1(n5667), .A2(n5668), .ZN(w_d[202]) );
  NAND2_X2 U4811 ( .A1(w_q[170]), .A2(n7190), .ZN(n5668) );
  NAND2_X2 U4812 ( .A1(w_q[202]), .A2(n7249), .ZN(n5667) );
  NAND2_X2 U4813 ( .A1(n5669), .A2(n5670), .ZN(w_d[201]) );
  NAND2_X2 U4814 ( .A1(w_q[169]), .A2(n7190), .ZN(n5670) );
  NAND2_X2 U4815 ( .A1(w_q[201]), .A2(n7249), .ZN(n5669) );
  NAND2_X2 U4816 ( .A1(n5671), .A2(n5672), .ZN(w_d[200]) );
  NAND2_X2 U4817 ( .A1(w_q[168]), .A2(n7190), .ZN(n5672) );
  NAND2_X2 U4818 ( .A1(w_q[200]), .A2(n7249), .ZN(n5671) );
  NAND2_X2 U4820 ( .A1(w[1]), .A2(n7160), .ZN(n5675) );
  NAND2_X2 U4821 ( .A1(w_q[1]), .A2(n7249), .ZN(n5674) );
  NAND2_X2 U4824 ( .A1(w[19]), .A2(n7160), .ZN(n5678) );
  NAND2_X2 U4825 ( .A1(w_q[19]), .A2(n7249), .ZN(n5677) );
  NAND2_X2 U4827 ( .A1(n5679), .A2(n5680), .ZN(w_d[199]) );
  NAND2_X2 U4828 ( .A1(w_q[167]), .A2(n7190), .ZN(n5680) );
  NAND2_X2 U4829 ( .A1(w_q[199]), .A2(n7248), .ZN(n5679) );
  NAND2_X2 U4830 ( .A1(n5681), .A2(n5682), .ZN(w_d[198]) );
  NAND2_X2 U4831 ( .A1(w_q[166]), .A2(n7189), .ZN(n5682) );
  NAND2_X2 U4832 ( .A1(w_q[198]), .A2(n7248), .ZN(n5681) );
  NAND2_X2 U4833 ( .A1(n5683), .A2(n5684), .ZN(w_d[197]) );
  NAND2_X2 U4834 ( .A1(w_q[165]), .A2(n7189), .ZN(n5684) );
  NAND2_X2 U4835 ( .A1(w_q[197]), .A2(n7248), .ZN(n5683) );
  NAND2_X2 U4836 ( .A1(n5685), .A2(n5686), .ZN(w_d[196]) );
  NAND2_X2 U4837 ( .A1(w_q[164]), .A2(n7189), .ZN(n5686) );
  NAND2_X2 U4838 ( .A1(w_q[196]), .A2(n7248), .ZN(n5685) );
  NAND2_X2 U4839 ( .A1(n5687), .A2(n5688), .ZN(w_d[195]) );
  NAND2_X2 U4840 ( .A1(w_q[163]), .A2(n7189), .ZN(n5688) );
  NAND2_X2 U4841 ( .A1(w_q[195]), .A2(n7248), .ZN(n5687) );
  NAND2_X2 U4842 ( .A1(n5689), .A2(n5690), .ZN(w_d[194]) );
  NAND2_X2 U4843 ( .A1(w_q[162]), .A2(n7189), .ZN(n5690) );
  NAND2_X2 U4844 ( .A1(w_q[194]), .A2(n7248), .ZN(n5689) );
  NAND2_X2 U4845 ( .A1(n5691), .A2(n5692), .ZN(w_d[193]) );
  NAND2_X2 U4846 ( .A1(w_q[161]), .A2(n7189), .ZN(n5692) );
  NAND2_X2 U4847 ( .A1(w_q[193]), .A2(n7248), .ZN(n5691) );
  NAND2_X2 U4848 ( .A1(n5693), .A2(n5694), .ZN(w_d[192]) );
  NAND2_X2 U4849 ( .A1(w_q[160]), .A2(n7189), .ZN(n5694) );
  NAND2_X2 U4850 ( .A1(w_q[192]), .A2(n7248), .ZN(n5693) );
  NAND2_X2 U4851 ( .A1(n5695), .A2(n5696), .ZN(w_d[191]) );
  NAND2_X2 U4852 ( .A1(w_q[159]), .A2(n7189), .ZN(n5696) );
  NAND2_X2 U4853 ( .A1(w_q[191]), .A2(n7248), .ZN(n5695) );
  NAND2_X2 U4854 ( .A1(n5697), .A2(n5698), .ZN(w_d[190]) );
  NAND2_X2 U4855 ( .A1(w_q[158]), .A2(n7189), .ZN(n5698) );
  NAND2_X2 U4856 ( .A1(w_q[190]), .A2(n7248), .ZN(n5697) );
  NAND2_X2 U4858 ( .A1(w[18]), .A2(n7160), .ZN(n5701) );
  NAND2_X2 U4859 ( .A1(w_q[18]), .A2(n7248), .ZN(n5700) );
  NAND2_X2 U4861 ( .A1(n5702), .A2(n5703), .ZN(w_d[189]) );
  NAND2_X2 U4862 ( .A1(w_q[157]), .A2(n7189), .ZN(n5703) );
  NAND2_X2 U4863 ( .A1(w_q[189]), .A2(n7247), .ZN(n5702) );
  NAND2_X2 U4864 ( .A1(n5704), .A2(n5705), .ZN(w_d[188]) );
  NAND2_X2 U4865 ( .A1(w_q[156]), .A2(n7189), .ZN(n5705) );
  NAND2_X2 U4866 ( .A1(w_q[188]), .A2(n7247), .ZN(n5704) );
  NAND2_X2 U4867 ( .A1(n5706), .A2(n5707), .ZN(w_d[187]) );
  NAND2_X2 U4868 ( .A1(w_q[155]), .A2(n7188), .ZN(n5707) );
  NAND2_X2 U4869 ( .A1(w_q[187]), .A2(n7247), .ZN(n5706) );
  NAND2_X2 U4870 ( .A1(n5708), .A2(n5709), .ZN(w_d[186]) );
  NAND2_X2 U4871 ( .A1(w_q[154]), .A2(n7188), .ZN(n5709) );
  NAND2_X2 U4872 ( .A1(w_q[186]), .A2(n7247), .ZN(n5708) );
  NAND2_X2 U4873 ( .A1(n5710), .A2(n5711), .ZN(w_d[185]) );
  NAND2_X2 U4874 ( .A1(w_q[153]), .A2(n7188), .ZN(n5711) );
  NAND2_X2 U4875 ( .A1(w_q[185]), .A2(n7247), .ZN(n5710) );
  NAND2_X2 U4876 ( .A1(n5712), .A2(n5713), .ZN(w_d[184]) );
  NAND2_X2 U4877 ( .A1(w_q[152]), .A2(n7188), .ZN(n5713) );
  NAND2_X2 U4878 ( .A1(w_q[184]), .A2(n7247), .ZN(n5712) );
  NAND2_X2 U4879 ( .A1(n5714), .A2(n5715), .ZN(w_d[183]) );
  NAND2_X2 U4880 ( .A1(w_q[151]), .A2(n7188), .ZN(n5715) );
  NAND2_X2 U4881 ( .A1(w_q[183]), .A2(n7247), .ZN(n5714) );
  NAND2_X2 U4882 ( .A1(n5716), .A2(n5717), .ZN(w_d[182]) );
  NAND2_X2 U4883 ( .A1(w_q[150]), .A2(n7188), .ZN(n5717) );
  NAND2_X2 U4884 ( .A1(w_q[182]), .A2(n7247), .ZN(n5716) );
  NAND2_X2 U4885 ( .A1(n5718), .A2(n5719), .ZN(w_d[181]) );
  NAND2_X2 U4886 ( .A1(w_q[149]), .A2(n7188), .ZN(n5719) );
  NAND2_X2 U4887 ( .A1(w_q[181]), .A2(n7247), .ZN(n5718) );
  NAND2_X2 U4888 ( .A1(n5720), .A2(n5721), .ZN(w_d[180]) );
  NAND2_X2 U4889 ( .A1(w_q[148]), .A2(n7188), .ZN(n5721) );
  NAND2_X2 U4890 ( .A1(w_q[180]), .A2(n7247), .ZN(n5720) );
  NAND2_X2 U4892 ( .A1(w[17]), .A2(n7160), .ZN(n5724) );
  NAND2_X2 U4893 ( .A1(w_q[17]), .A2(n7247), .ZN(n5723) );
  NAND2_X2 U4895 ( .A1(n5725), .A2(n5726), .ZN(w_d[179]) );
  NAND2_X2 U4896 ( .A1(w_q[147]), .A2(n7188), .ZN(n5726) );
  NAND2_X2 U4897 ( .A1(w_q[179]), .A2(n7246), .ZN(n5725) );
  NAND2_X2 U4898 ( .A1(n5727), .A2(n5728), .ZN(w_d[178]) );
  NAND2_X2 U4899 ( .A1(w_q[146]), .A2(n7188), .ZN(n5728) );
  NAND2_X2 U4900 ( .A1(w_q[178]), .A2(n7246), .ZN(n5727) );
  NAND2_X2 U4901 ( .A1(n5729), .A2(n5730), .ZN(w_d[177]) );
  NAND2_X2 U4902 ( .A1(w_q[145]), .A2(n7188), .ZN(n5730) );
  NAND2_X2 U4903 ( .A1(w_q[177]), .A2(n7246), .ZN(n5729) );
  NAND2_X2 U4904 ( .A1(n5731), .A2(n5732), .ZN(w_d[176]) );
  NAND2_X2 U4905 ( .A1(w_q[144]), .A2(n7187), .ZN(n5732) );
  NAND2_X2 U4906 ( .A1(w_q[176]), .A2(n7246), .ZN(n5731) );
  NAND2_X2 U4907 ( .A1(n5733), .A2(n5734), .ZN(w_d[175]) );
  NAND2_X2 U4908 ( .A1(w_q[143]), .A2(n7187), .ZN(n5734) );
  NAND2_X2 U4909 ( .A1(w_q[175]), .A2(n7246), .ZN(n5733) );
  NAND2_X2 U4910 ( .A1(n5735), .A2(n5736), .ZN(w_d[174]) );
  NAND2_X2 U4911 ( .A1(w_q[142]), .A2(n7187), .ZN(n5736) );
  NAND2_X2 U4912 ( .A1(w_q[174]), .A2(n7246), .ZN(n5735) );
  NAND2_X2 U4913 ( .A1(n5737), .A2(n5738), .ZN(w_d[173]) );
  NAND2_X2 U4914 ( .A1(w_q[141]), .A2(n7187), .ZN(n5738) );
  NAND2_X2 U4915 ( .A1(w_q[173]), .A2(n7246), .ZN(n5737) );
  NAND2_X2 U4916 ( .A1(n5739), .A2(n5740), .ZN(w_d[172]) );
  NAND2_X2 U4917 ( .A1(w_q[140]), .A2(n7187), .ZN(n5740) );
  NAND2_X2 U4918 ( .A1(w_q[172]), .A2(n7246), .ZN(n5739) );
  NAND2_X2 U4919 ( .A1(n5741), .A2(n5742), .ZN(w_d[171]) );
  NAND2_X2 U4920 ( .A1(w_q[139]), .A2(n7187), .ZN(n5742) );
  NAND2_X2 U4921 ( .A1(w_q[171]), .A2(n7246), .ZN(n5741) );
  NAND2_X2 U4922 ( .A1(n5743), .A2(n5744), .ZN(w_d[170]) );
  NAND2_X2 U4923 ( .A1(w_q[138]), .A2(n7187), .ZN(n5744) );
  NAND2_X2 U4924 ( .A1(w_q[170]), .A2(n7246), .ZN(n5743) );
  NAND2_X2 U4926 ( .A1(w[16]), .A2(n7160), .ZN(n5747) );
  NAND2_X2 U4927 ( .A1(w_q[16]), .A2(n7246), .ZN(n5746) );
  NAND2_X2 U4929 ( .A1(n5748), .A2(n5749), .ZN(w_d[169]) );
  NAND2_X2 U4930 ( .A1(w_q[137]), .A2(n7187), .ZN(n5749) );
  NAND2_X2 U4931 ( .A1(w_q[169]), .A2(n7245), .ZN(n5748) );
  NAND2_X2 U4932 ( .A1(n5750), .A2(n5751), .ZN(w_d[168]) );
  NAND2_X2 U4933 ( .A1(w_q[136]), .A2(n7187), .ZN(n5751) );
  NAND2_X2 U4934 ( .A1(w_q[168]), .A2(n7245), .ZN(n5750) );
  NAND2_X2 U4935 ( .A1(n5752), .A2(n5753), .ZN(w_d[167]) );
  NAND2_X2 U4936 ( .A1(w_q[135]), .A2(n7187), .ZN(n5753) );
  NAND2_X2 U4937 ( .A1(w_q[167]), .A2(n7245), .ZN(n5752) );
  NAND2_X2 U4938 ( .A1(n5754), .A2(n5755), .ZN(w_d[166]) );
  NAND2_X2 U4939 ( .A1(w_q[134]), .A2(n7187), .ZN(n5755) );
  NAND2_X2 U4940 ( .A1(w_q[166]), .A2(n7245), .ZN(n5754) );
  NAND2_X2 U4941 ( .A1(n5756), .A2(n5757), .ZN(w_d[165]) );
  NAND2_X2 U4942 ( .A1(w_q[133]), .A2(n7186), .ZN(n5757) );
  NAND2_X2 U4943 ( .A1(w_q[165]), .A2(n7245), .ZN(n5756) );
  NAND2_X2 U4944 ( .A1(n5758), .A2(n5759), .ZN(w_d[164]) );
  NAND2_X2 U4945 ( .A1(w_q[132]), .A2(n7186), .ZN(n5759) );
  NAND2_X2 U4946 ( .A1(w_q[164]), .A2(n7245), .ZN(n5758) );
  NAND2_X2 U4947 ( .A1(n5760), .A2(n5761), .ZN(w_d[163]) );
  NAND2_X2 U4948 ( .A1(w_q[131]), .A2(n7186), .ZN(n5761) );
  NAND2_X2 U4949 ( .A1(w_q[163]), .A2(n7245), .ZN(n5760) );
  NAND2_X2 U4950 ( .A1(n5762), .A2(n5763), .ZN(w_d[162]) );
  NAND2_X2 U4951 ( .A1(w_q[130]), .A2(n7186), .ZN(n5763) );
  NAND2_X2 U4952 ( .A1(w_q[162]), .A2(n7245), .ZN(n5762) );
  NAND2_X2 U4953 ( .A1(n5764), .A2(n5765), .ZN(w_d[161]) );
  NAND2_X2 U4954 ( .A1(w_q[129]), .A2(n7186), .ZN(n5765) );
  NAND2_X2 U4955 ( .A1(w_q[161]), .A2(n7245), .ZN(n5764) );
  NAND2_X2 U4956 ( .A1(n5766), .A2(n5767), .ZN(w_d[160]) );
  NAND2_X2 U4957 ( .A1(w_q[128]), .A2(n7186), .ZN(n5767) );
  NAND2_X2 U4958 ( .A1(w_q[160]), .A2(n7245), .ZN(n5766) );
  NAND2_X2 U4960 ( .A1(w[15]), .A2(n7160), .ZN(n5770) );
  NAND2_X2 U4961 ( .A1(w_q[15]), .A2(n7245), .ZN(n5769) );
  NAND2_X2 U4963 ( .A1(n5771), .A2(n5772), .ZN(w_d[159]) );
  NAND2_X2 U4964 ( .A1(w_q[127]), .A2(n7186), .ZN(n5772) );
  NAND2_X2 U4965 ( .A1(w_q[159]), .A2(n7244), .ZN(n5771) );
  NAND2_X2 U4966 ( .A1(n5773), .A2(n5774), .ZN(w_d[158]) );
  NAND2_X2 U4967 ( .A1(w_q[126]), .A2(n7186), .ZN(n5774) );
  NAND2_X2 U4968 ( .A1(w_q[158]), .A2(n7244), .ZN(n5773) );
  NAND2_X2 U4969 ( .A1(n5775), .A2(n5776), .ZN(w_d[157]) );
  NAND2_X2 U4970 ( .A1(w_q[125]), .A2(n7186), .ZN(n5776) );
  NAND2_X2 U4971 ( .A1(w_q[157]), .A2(n7244), .ZN(n5775) );
  NAND2_X2 U4972 ( .A1(n5777), .A2(n5778), .ZN(w_d[156]) );
  NAND2_X2 U4973 ( .A1(w_q[124]), .A2(n7186), .ZN(n5778) );
  NAND2_X2 U4974 ( .A1(w_q[156]), .A2(n7244), .ZN(n5777) );
  NAND2_X2 U4975 ( .A1(n5779), .A2(n5780), .ZN(w_d[155]) );
  NAND2_X2 U4976 ( .A1(w_q[123]), .A2(n7186), .ZN(n5780) );
  NAND2_X2 U4977 ( .A1(w_q[155]), .A2(n7244), .ZN(n5779) );
  NAND2_X2 U4978 ( .A1(n5781), .A2(n5782), .ZN(w_d[154]) );
  NAND2_X2 U4979 ( .A1(w_q[122]), .A2(n7185), .ZN(n5782) );
  NAND2_X2 U4980 ( .A1(w_q[154]), .A2(n7244), .ZN(n5781) );
  NAND2_X2 U4981 ( .A1(n5783), .A2(n5784), .ZN(w_d[153]) );
  NAND2_X2 U4982 ( .A1(w_q[121]), .A2(n7185), .ZN(n5784) );
  NAND2_X2 U4983 ( .A1(w_q[153]), .A2(n7244), .ZN(n5783) );
  NAND2_X2 U4984 ( .A1(n5785), .A2(n5786), .ZN(w_d[152]) );
  NAND2_X2 U4985 ( .A1(w_q[120]), .A2(n7185), .ZN(n5786) );
  NAND2_X2 U4986 ( .A1(w_q[152]), .A2(n7244), .ZN(n5785) );
  NAND2_X2 U4987 ( .A1(n5787), .A2(n5788), .ZN(w_d[151]) );
  NAND2_X2 U4988 ( .A1(w_q[119]), .A2(n7185), .ZN(n5788) );
  NAND2_X2 U4989 ( .A1(w_q[151]), .A2(n7244), .ZN(n5787) );
  NAND2_X2 U4990 ( .A1(n5789), .A2(n5790), .ZN(w_d[150]) );
  NAND2_X2 U4991 ( .A1(w_q[118]), .A2(n7185), .ZN(n5790) );
  NAND2_X2 U4992 ( .A1(w_q[150]), .A2(n7244), .ZN(n5789) );
  NAND2_X2 U4994 ( .A1(w[14]), .A2(n7160), .ZN(n5793) );
  NAND2_X2 U4995 ( .A1(w_q[14]), .A2(n7244), .ZN(n5792) );
  NAND2_X2 U4997 ( .A1(n5794), .A2(n5795), .ZN(w_d[149]) );
  NAND2_X2 U4998 ( .A1(w_q[117]), .A2(n7185), .ZN(n5795) );
  NAND2_X2 U4999 ( .A1(w_q[149]), .A2(n7243), .ZN(n5794) );
  NAND2_X2 U5000 ( .A1(n5796), .A2(n5797), .ZN(w_d[148]) );
  NAND2_X2 U5001 ( .A1(w_q[116]), .A2(n7185), .ZN(n5797) );
  NAND2_X2 U5002 ( .A1(w_q[148]), .A2(n7243), .ZN(n5796) );
  NAND2_X2 U5003 ( .A1(n5798), .A2(n5799), .ZN(w_d[147]) );
  NAND2_X2 U5004 ( .A1(w_q[115]), .A2(n7185), .ZN(n5799) );
  NAND2_X2 U5005 ( .A1(w_q[147]), .A2(n7243), .ZN(n5798) );
  NAND2_X2 U5006 ( .A1(n5800), .A2(n5801), .ZN(w_d[146]) );
  NAND2_X2 U5007 ( .A1(w_q[114]), .A2(n7185), .ZN(n5801) );
  NAND2_X2 U5008 ( .A1(w_q[146]), .A2(n7243), .ZN(n5800) );
  NAND2_X2 U5009 ( .A1(n5802), .A2(n5803), .ZN(w_d[145]) );
  NAND2_X2 U5010 ( .A1(w_q[113]), .A2(n7185), .ZN(n5803) );
  NAND2_X2 U5011 ( .A1(w_q[145]), .A2(n7243), .ZN(n5802) );
  NAND2_X2 U5012 ( .A1(n5804), .A2(n5805), .ZN(w_d[144]) );
  NAND2_X2 U5013 ( .A1(w_q[112]), .A2(n7185), .ZN(n5805) );
  NAND2_X2 U5014 ( .A1(w_q[144]), .A2(n7243), .ZN(n5804) );
  NAND2_X2 U5015 ( .A1(n5806), .A2(n5807), .ZN(w_d[143]) );
  NAND2_X2 U5016 ( .A1(w_q[111]), .A2(n7184), .ZN(n5807) );
  NAND2_X2 U5017 ( .A1(w_q[143]), .A2(n7243), .ZN(n5806) );
  NAND2_X2 U5018 ( .A1(n5808), .A2(n5809), .ZN(w_d[142]) );
  NAND2_X2 U5019 ( .A1(w_q[110]), .A2(n7184), .ZN(n5809) );
  NAND2_X2 U5020 ( .A1(w_q[142]), .A2(n7243), .ZN(n5808) );
  NAND2_X2 U5021 ( .A1(n5810), .A2(n5811), .ZN(w_d[141]) );
  NAND2_X2 U5022 ( .A1(w_q[109]), .A2(n7184), .ZN(n5811) );
  NAND2_X2 U5023 ( .A1(w_q[141]), .A2(n7243), .ZN(n5810) );
  NAND2_X2 U5024 ( .A1(n5812), .A2(n5813), .ZN(w_d[140]) );
  NAND2_X2 U5025 ( .A1(w_q[108]), .A2(n7184), .ZN(n5813) );
  NAND2_X2 U5026 ( .A1(w_q[140]), .A2(n7243), .ZN(n5812) );
  NAND2_X2 U5028 ( .A1(w[13]), .A2(n7160), .ZN(n5816) );
  NAND2_X2 U5029 ( .A1(w_q[13]), .A2(n7243), .ZN(n5815) );
  NAND2_X2 U5031 ( .A1(n5817), .A2(n5818), .ZN(w_d[139]) );
  NAND2_X2 U5032 ( .A1(w_q[107]), .A2(n7184), .ZN(n5818) );
  NAND2_X2 U5033 ( .A1(w_q[139]), .A2(n7242), .ZN(n5817) );
  NAND2_X2 U5034 ( .A1(n5819), .A2(n5820), .ZN(w_d[138]) );
  NAND2_X2 U5035 ( .A1(w_q[106]), .A2(n7184), .ZN(n5820) );
  NAND2_X2 U5036 ( .A1(w_q[138]), .A2(n7242), .ZN(n5819) );
  NAND2_X2 U5037 ( .A1(n5821), .A2(n5822), .ZN(w_d[137]) );
  NAND2_X2 U5038 ( .A1(w_q[105]), .A2(n7184), .ZN(n5822) );
  NAND2_X2 U5039 ( .A1(w_q[137]), .A2(n7242), .ZN(n5821) );
  NAND2_X2 U5040 ( .A1(n5823), .A2(n5824), .ZN(w_d[136]) );
  NAND2_X2 U5041 ( .A1(w_q[104]), .A2(n7184), .ZN(n5824) );
  NAND2_X2 U5042 ( .A1(w_q[136]), .A2(n7242), .ZN(n5823) );
  NAND2_X2 U5043 ( .A1(n5825), .A2(n5826), .ZN(w_d[135]) );
  NAND2_X2 U5044 ( .A1(w_q[103]), .A2(n7184), .ZN(n5826) );
  NAND2_X2 U5045 ( .A1(w_q[135]), .A2(n7242), .ZN(n5825) );
  NAND2_X2 U5046 ( .A1(n5827), .A2(n5828), .ZN(w_d[134]) );
  NAND2_X2 U5047 ( .A1(w_q[102]), .A2(n7184), .ZN(n5828) );
  NAND2_X2 U5048 ( .A1(w_q[134]), .A2(n7242), .ZN(n5827) );
  NAND2_X2 U5049 ( .A1(n5829), .A2(n5830), .ZN(w_d[133]) );
  NAND2_X2 U5050 ( .A1(w_q[101]), .A2(n7184), .ZN(n5830) );
  NAND2_X2 U5051 ( .A1(w_q[133]), .A2(n7242), .ZN(n5829) );
  NAND2_X2 U5052 ( .A1(n5831), .A2(n5832), .ZN(w_d[132]) );
  NAND2_X2 U5053 ( .A1(w_q[100]), .A2(n7183), .ZN(n5832) );
  NAND2_X2 U5054 ( .A1(w_q[132]), .A2(n7242), .ZN(n5831) );
  NAND2_X2 U5055 ( .A1(n5833), .A2(n5834), .ZN(w_d[131]) );
  NAND2_X2 U5056 ( .A1(w_q[99]), .A2(n7183), .ZN(n5834) );
  NAND2_X2 U5057 ( .A1(w_q[131]), .A2(n7242), .ZN(n5833) );
  NAND2_X2 U5058 ( .A1(n5835), .A2(n5836), .ZN(w_d[130]) );
  NAND2_X2 U5059 ( .A1(w_q[98]), .A2(n7183), .ZN(n5836) );
  NAND2_X2 U5060 ( .A1(w_q[130]), .A2(n7242), .ZN(n5835) );
  NAND2_X2 U5062 ( .A1(w[12]), .A2(n7160), .ZN(n5839) );
  NAND2_X2 U5063 ( .A1(w_q[12]), .A2(n7242), .ZN(n5838) );
  NAND2_X2 U5065 ( .A1(n5840), .A2(n5841), .ZN(w_d[129]) );
  NAND2_X2 U5066 ( .A1(w_q[97]), .A2(n7183), .ZN(n5841) );
  NAND2_X2 U5067 ( .A1(w_q[129]), .A2(n7241), .ZN(n5840) );
  NAND2_X2 U5068 ( .A1(n5842), .A2(n5843), .ZN(w_d[128]) );
  NAND2_X2 U5069 ( .A1(w_q[96]), .A2(n7183), .ZN(n5843) );
  NAND2_X2 U5070 ( .A1(w_q[128]), .A2(n7241), .ZN(n5842) );
  NAND2_X2 U5071 ( .A1(n5844), .A2(n5845), .ZN(w_d[127]) );
  NAND2_X2 U5072 ( .A1(w_q[95]), .A2(n7183), .ZN(n5845) );
  NAND2_X2 U5073 ( .A1(w_q[127]), .A2(n7241), .ZN(n5844) );
  NAND2_X2 U5074 ( .A1(n5846), .A2(n5847), .ZN(w_d[126]) );
  NAND2_X2 U5075 ( .A1(w_q[94]), .A2(n7183), .ZN(n5847) );
  NAND2_X2 U5076 ( .A1(w_q[126]), .A2(n7241), .ZN(n5846) );
  NAND2_X2 U5077 ( .A1(n5848), .A2(n5849), .ZN(w_d[125]) );
  NAND2_X2 U5078 ( .A1(w_q[93]), .A2(n7183), .ZN(n5849) );
  NAND2_X2 U5079 ( .A1(w_q[125]), .A2(n7241), .ZN(n5848) );
  NAND2_X2 U5080 ( .A1(n5850), .A2(n5851), .ZN(w_d[124]) );
  NAND2_X2 U5081 ( .A1(w_q[92]), .A2(n7183), .ZN(n5851) );
  NAND2_X2 U5082 ( .A1(w_q[124]), .A2(n7241), .ZN(n5850) );
  NAND2_X2 U5083 ( .A1(n5852), .A2(n5853), .ZN(w_d[123]) );
  NAND2_X2 U5084 ( .A1(w_q[91]), .A2(n7183), .ZN(n5853) );
  NAND2_X2 U5085 ( .A1(w_q[123]), .A2(n7241), .ZN(n5852) );
  NAND2_X2 U5086 ( .A1(n5854), .A2(n5855), .ZN(w_d[122]) );
  NAND2_X2 U5087 ( .A1(w_q[90]), .A2(n7183), .ZN(n5855) );
  NAND2_X2 U5088 ( .A1(w_q[122]), .A2(n7241), .ZN(n5854) );
  NAND2_X2 U5089 ( .A1(n5856), .A2(n5857), .ZN(w_d[121]) );
  NAND2_X2 U5090 ( .A1(w_q[89]), .A2(n7216), .ZN(n5857) );
  NAND2_X2 U5091 ( .A1(w_q[121]), .A2(n7241), .ZN(n5856) );
  NAND2_X2 U5092 ( .A1(n5858), .A2(n5859), .ZN(w_d[120]) );
  NAND2_X2 U5093 ( .A1(w_q[88]), .A2(n7216), .ZN(n5859) );
  NAND2_X2 U5094 ( .A1(w_q[120]), .A2(n7241), .ZN(n5858) );
  NAND2_X2 U5096 ( .A1(w[11]), .A2(n7160), .ZN(n5862) );
  NAND2_X2 U5097 ( .A1(w_q[11]), .A2(n7241), .ZN(n5861) );
  NAND2_X2 U5099 ( .A1(n5863), .A2(n5864), .ZN(w_d[119]) );
  NAND2_X2 U5100 ( .A1(w_q[87]), .A2(n7216), .ZN(n5864) );
  NAND2_X2 U5101 ( .A1(w_q[119]), .A2(n7240), .ZN(n5863) );
  NAND2_X2 U5102 ( .A1(n5865), .A2(n5866), .ZN(w_d[118]) );
  NAND2_X2 U5103 ( .A1(w_q[86]), .A2(n7182), .ZN(n5866) );
  NAND2_X2 U5104 ( .A1(w_q[118]), .A2(n7240), .ZN(n5865) );
  NAND2_X2 U5105 ( .A1(n5867), .A2(n5868), .ZN(w_d[117]) );
  NAND2_X2 U5106 ( .A1(w_q[85]), .A2(n7226), .ZN(n5868) );
  NAND2_X2 U5107 ( .A1(w_q[117]), .A2(n7240), .ZN(n5867) );
  NAND2_X2 U5108 ( .A1(n5869), .A2(n5870), .ZN(w_d[116]) );
  NAND2_X2 U5109 ( .A1(w_q[84]), .A2(n7216), .ZN(n5870) );
  NAND2_X2 U5110 ( .A1(w_q[116]), .A2(n7240), .ZN(n5869) );
  NAND2_X2 U5111 ( .A1(n5871), .A2(n5872), .ZN(w_d[115]) );
  NAND2_X2 U5112 ( .A1(w_q[83]), .A2(n7216), .ZN(n5872) );
  NAND2_X2 U5113 ( .A1(w_q[115]), .A2(n7240), .ZN(n5871) );
  NAND2_X2 U5114 ( .A1(n5873), .A2(n5874), .ZN(w_d[114]) );
  NAND2_X2 U5115 ( .A1(w_q[82]), .A2(n7226), .ZN(n5874) );
  NAND2_X2 U5116 ( .A1(w_q[114]), .A2(n7240), .ZN(n5873) );
  NAND2_X2 U5117 ( .A1(n5875), .A2(n5876), .ZN(w_d[113]) );
  NAND2_X2 U5118 ( .A1(w_q[81]), .A2(n7214), .ZN(n5876) );
  NAND2_X2 U5119 ( .A1(w_q[113]), .A2(n7240), .ZN(n5875) );
  NAND2_X2 U5120 ( .A1(n5877), .A2(n5878), .ZN(w_d[112]) );
  NAND2_X2 U5121 ( .A1(w_q[80]), .A2(n7183), .ZN(n5878) );
  NAND2_X2 U5122 ( .A1(w_q[112]), .A2(n7240), .ZN(n5877) );
  NAND2_X2 U5123 ( .A1(n5879), .A2(n5880), .ZN(w_d[111]) );
  NAND2_X2 U5124 ( .A1(w_q[79]), .A2(n7184), .ZN(n5880) );
  NAND2_X2 U5125 ( .A1(w_q[111]), .A2(n7240), .ZN(n5879) );
  NAND2_X2 U5126 ( .A1(n5881), .A2(n5882), .ZN(w_d[110]) );
  NAND2_X2 U5127 ( .A1(w_q[78]), .A2(n7182), .ZN(n5882) );
  NAND2_X2 U5128 ( .A1(w_q[110]), .A2(n7240), .ZN(n5881) );
  NAND2_X2 U5130 ( .A1(w[10]), .A2(n7160), .ZN(n5885) );
  NAND2_X2 U5131 ( .A1(w_q[10]), .A2(n7240), .ZN(n5884) );
  NAND2_X2 U5133 ( .A1(n5886), .A2(n5887), .ZN(w_d[109]) );
  NAND2_X2 U5134 ( .A1(w_q[77]), .A2(n7182), .ZN(n5887) );
  NAND2_X2 U5135 ( .A1(w_q[109]), .A2(n7239), .ZN(n5886) );
  NAND2_X2 U5136 ( .A1(n5888), .A2(n5889), .ZN(w_d[108]) );
  NAND2_X2 U5137 ( .A1(w_q[76]), .A2(n7182), .ZN(n5889) );
  NAND2_X2 U5138 ( .A1(w_q[108]), .A2(n7239), .ZN(n5888) );
  NAND2_X2 U5139 ( .A1(n5890), .A2(n5891), .ZN(w_d[107]) );
  NAND2_X2 U5140 ( .A1(w_q[75]), .A2(n7182), .ZN(n5891) );
  NAND2_X2 U5141 ( .A1(w_q[107]), .A2(n7239), .ZN(n5890) );
  NAND2_X2 U5142 ( .A1(n5892), .A2(n5893), .ZN(w_d[106]) );
  NAND2_X2 U5143 ( .A1(w_q[74]), .A2(n7182), .ZN(n5893) );
  NAND2_X2 U5144 ( .A1(w_q[106]), .A2(n7239), .ZN(n5892) );
  NAND2_X2 U5145 ( .A1(n5894), .A2(n5895), .ZN(w_d[105]) );
  NAND2_X2 U5146 ( .A1(w_q[73]), .A2(n7182), .ZN(n5895) );
  NAND2_X2 U5147 ( .A1(w_q[105]), .A2(n7239), .ZN(n5894) );
  NAND2_X2 U5148 ( .A1(n5896), .A2(n5897), .ZN(w_d[104]) );
  NAND2_X2 U5149 ( .A1(w_q[72]), .A2(n7182), .ZN(n5897) );
  NAND2_X2 U5150 ( .A1(w_q[104]), .A2(n7239), .ZN(n5896) );
  NAND2_X2 U5151 ( .A1(n5898), .A2(n5899), .ZN(w_d[103]) );
  NAND2_X2 U5152 ( .A1(w_q[71]), .A2(n7182), .ZN(n5899) );
  NAND2_X2 U5153 ( .A1(w_q[103]), .A2(n7239), .ZN(n5898) );
  NAND2_X2 U5154 ( .A1(n5900), .A2(n5901), .ZN(w_d[102]) );
  NAND2_X2 U5155 ( .A1(w_q[70]), .A2(n7182), .ZN(n5901) );
  NAND2_X2 U5156 ( .A1(w_q[102]), .A2(n7239), .ZN(n5900) );
  NAND2_X2 U5157 ( .A1(n5902), .A2(n5903), .ZN(w_d[101]) );
  NAND2_X2 U5158 ( .A1(w_q[69]), .A2(n7182), .ZN(n5903) );
  NAND2_X2 U5159 ( .A1(w_q[101]), .A2(n7239), .ZN(n5902) );
  NAND2_X2 U5160 ( .A1(n5904), .A2(n5905), .ZN(w_d[100]) );
  NAND2_X2 U5161 ( .A1(w_q[68]), .A2(n7182), .ZN(n5905) );
  NAND2_X2 U5163 ( .A1(w_q[100]), .A2(n7239), .ZN(n5904) );
  NAND2_X2 U5165 ( .A1(w[0]), .A2(n7160), .ZN(n5908) );
  NAND2_X2 U5166 ( .A1(w_q[0]), .A2(n7239), .ZN(n5907) );
  NAND2_X2 U5170 ( .A1(n5909), .A2(n5910), .ZN(rnd_d[9]) );
  NAND2_X2 U5171 ( .A1(sha1_round_wire[9]), .A2(n7160), .ZN(n5910) );
  NAND2_X2 U5172 ( .A1(n5911), .A2(n5912), .ZN(rnd_d[99]) );
  NAND2_X2 U5173 ( .A1(sha1_round_wire[99]), .A2(n7160), .ZN(n5912) );
  NAND2_X2 U5174 ( .A1(n5913), .A2(n5914), .ZN(rnd_d[98]) );
  NAND2_X2 U5175 ( .A1(sha1_round_wire[98]), .A2(n7160), .ZN(n5914) );
  NAND2_X2 U5176 ( .A1(n5915), .A2(n5916), .ZN(rnd_d[97]) );
  NAND2_X2 U5177 ( .A1(sha1_round_wire[97]), .A2(n7160), .ZN(n5916) );
  NAND2_X2 U5178 ( .A1(n5917), .A2(n5918), .ZN(rnd_d[96]) );
  NAND2_X2 U5179 ( .A1(sha1_round_wire[96]), .A2(n7160), .ZN(n5918) );
  NAND2_X2 U5180 ( .A1(n5919), .A2(n5920), .ZN(rnd_d[95]) );
  NAND2_X2 U5181 ( .A1(sha1_round_wire[95]), .A2(n7160), .ZN(n5920) );
  NAND2_X2 U5182 ( .A1(n5921), .A2(n5922), .ZN(rnd_d[94]) );
  NAND2_X2 U5183 ( .A1(sha1_round_wire[94]), .A2(n7160), .ZN(n5922) );
  NAND2_X2 U5184 ( .A1(n5923), .A2(n5924), .ZN(rnd_d[93]) );
  NAND2_X2 U5185 ( .A1(sha1_round_wire[93]), .A2(n7160), .ZN(n5924) );
  NAND2_X2 U5186 ( .A1(n5925), .A2(n5926), .ZN(rnd_d[92]) );
  NAND2_X2 U5187 ( .A1(sha1_round_wire[92]), .A2(n7161), .ZN(n5926) );
  NAND2_X2 U5188 ( .A1(n5927), .A2(n5928), .ZN(rnd_d[91]) );
  NAND2_X2 U5189 ( .A1(sha1_round_wire[91]), .A2(n7161), .ZN(n5928) );
  NAND2_X2 U5190 ( .A1(n5929), .A2(n5930), .ZN(rnd_d[90]) );
  NAND2_X2 U5191 ( .A1(sha1_round_wire[90]), .A2(n7161), .ZN(n5930) );
  NAND2_X2 U5192 ( .A1(n5931), .A2(n5932), .ZN(rnd_d[8]) );
  NAND2_X2 U5193 ( .A1(sha1_round_wire[8]), .A2(n7161), .ZN(n5932) );
  NAND2_X2 U5194 ( .A1(n5933), .A2(n5934), .ZN(rnd_d[89]) );
  NAND2_X2 U5195 ( .A1(sha1_round_wire[89]), .A2(n7161), .ZN(n5934) );
  NAND2_X2 U5196 ( .A1(n5935), .A2(n5936), .ZN(rnd_d[88]) );
  NAND2_X2 U5197 ( .A1(sha1_round_wire[88]), .A2(n7161), .ZN(n5936) );
  NAND2_X2 U5198 ( .A1(n5937), .A2(n5938), .ZN(rnd_d[87]) );
  NAND2_X2 U5199 ( .A1(sha1_round_wire[87]), .A2(n7161), .ZN(n5938) );
  NAND2_X2 U5200 ( .A1(n5939), .A2(n5940), .ZN(rnd_d[86]) );
  NAND2_X2 U5201 ( .A1(sha1_round_wire[86]), .A2(n7161), .ZN(n5940) );
  NAND2_X2 U5202 ( .A1(n5941), .A2(n5942), .ZN(rnd_d[85]) );
  NAND2_X2 U5203 ( .A1(sha1_round_wire[85]), .A2(n7161), .ZN(n5942) );
  NAND2_X2 U5204 ( .A1(n5943), .A2(n5944), .ZN(rnd_d[84]) );
  NAND2_X2 U5205 ( .A1(sha1_round_wire[84]), .A2(n7161), .ZN(n5944) );
  NAND2_X2 U5206 ( .A1(n5945), .A2(n5946), .ZN(rnd_d[83]) );
  NAND2_X2 U5207 ( .A1(sha1_round_wire[83]), .A2(n7161), .ZN(n5946) );
  NAND2_X2 U5208 ( .A1(n5947), .A2(n5948), .ZN(rnd_d[82]) );
  NAND2_X2 U5209 ( .A1(sha1_round_wire[82]), .A2(n7161), .ZN(n5948) );
  NAND2_X2 U5210 ( .A1(n5949), .A2(n5950), .ZN(rnd_d[81]) );
  NAND2_X2 U5211 ( .A1(sha1_round_wire[81]), .A2(n7161), .ZN(n5950) );
  NAND2_X2 U5212 ( .A1(n5951), .A2(n5952), .ZN(rnd_d[80]) );
  NAND2_X2 U5213 ( .A1(sha1_round_wire[80]), .A2(n7161), .ZN(n5952) );
  NAND2_X2 U5214 ( .A1(n5953), .A2(n5954), .ZN(rnd_d[7]) );
  NAND2_X2 U5215 ( .A1(sha1_round_wire[7]), .A2(n7161), .ZN(n5954) );
  NAND2_X2 U5216 ( .A1(n5955), .A2(n5956), .ZN(rnd_d[79]) );
  NAND2_X2 U5217 ( .A1(sha1_round_wire[79]), .A2(n7161), .ZN(n5956) );
  NAND2_X2 U5218 ( .A1(n5957), .A2(n5958), .ZN(rnd_d[78]) );
  NAND2_X2 U5219 ( .A1(sha1_round_wire[78]), .A2(n7161), .ZN(n5958) );
  NAND2_X2 U5220 ( .A1(n5959), .A2(n5960), .ZN(rnd_d[77]) );
  NAND2_X2 U5221 ( .A1(sha1_round_wire[77]), .A2(n7161), .ZN(n5960) );
  NAND2_X2 U5222 ( .A1(n5961), .A2(n5962), .ZN(rnd_d[76]) );
  NAND2_X2 U5223 ( .A1(sha1_round_wire[76]), .A2(n7161), .ZN(n5962) );
  NAND2_X2 U5224 ( .A1(n5963), .A2(n5964), .ZN(rnd_d[75]) );
  NAND2_X2 U5225 ( .A1(sha1_round_wire[75]), .A2(n7161), .ZN(n5964) );
  NAND2_X2 U5226 ( .A1(n5965), .A2(n5966), .ZN(rnd_d[74]) );
  NAND2_X2 U5227 ( .A1(sha1_round_wire[74]), .A2(n7161), .ZN(n5966) );
  NAND2_X2 U5228 ( .A1(n5967), .A2(n5968), .ZN(rnd_d[73]) );
  NAND2_X2 U5229 ( .A1(sha1_round_wire[73]), .A2(n7161), .ZN(n5968) );
  NAND2_X2 U5230 ( .A1(n5969), .A2(n5970), .ZN(rnd_d[72]) );
  NAND2_X2 U5231 ( .A1(sha1_round_wire[72]), .A2(n7161), .ZN(n5970) );
  NAND2_X2 U5232 ( .A1(n5971), .A2(n5972), .ZN(rnd_d[71]) );
  NAND2_X2 U5233 ( .A1(sha1_round_wire[71]), .A2(n7161), .ZN(n5972) );
  NAND2_X2 U5234 ( .A1(n5973), .A2(n5974), .ZN(rnd_d[70]) );
  NAND2_X2 U5235 ( .A1(sha1_round_wire[70]), .A2(n7161), .ZN(n5974) );
  NAND2_X2 U5236 ( .A1(n5975), .A2(n5976), .ZN(rnd_d[6]) );
  NAND2_X2 U5237 ( .A1(sha1_round_wire[6]), .A2(n7161), .ZN(n5976) );
  NAND2_X2 U5238 ( .A1(n5977), .A2(n5978), .ZN(rnd_d[69]) );
  NAND2_X2 U5239 ( .A1(sha1_round_wire[69]), .A2(n7161), .ZN(n5978) );
  NAND2_X2 U5240 ( .A1(n5979), .A2(n5980), .ZN(rnd_d[68]) );
  NAND2_X2 U5241 ( .A1(sha1_round_wire[68]), .A2(n7162), .ZN(n5980) );
  NAND2_X2 U5242 ( .A1(n5981), .A2(n5982), .ZN(rnd_d[67]) );
  NAND2_X2 U5243 ( .A1(sha1_round_wire[67]), .A2(n7162), .ZN(n5982) );
  NAND2_X2 U5244 ( .A1(n5983), .A2(n5984), .ZN(rnd_d[66]) );
  NAND2_X2 U5245 ( .A1(sha1_round_wire[66]), .A2(n7162), .ZN(n5984) );
  NAND2_X2 U5246 ( .A1(n5985), .A2(n5986), .ZN(rnd_d[65]) );
  NAND2_X2 U5247 ( .A1(sha1_round_wire[65]), .A2(n7162), .ZN(n5986) );
  NAND2_X2 U5248 ( .A1(n5987), .A2(n5988), .ZN(rnd_d[64]) );
  NAND2_X2 U5249 ( .A1(sha1_round_wire[64]), .A2(n7162), .ZN(n5988) );
  NAND2_X2 U5250 ( .A1(n5989), .A2(n5990), .ZN(rnd_d[63]) );
  NAND2_X2 U5251 ( .A1(sha1_round_wire[63]), .A2(n7162), .ZN(n5990) );
  NAND2_X2 U5252 ( .A1(n5991), .A2(n5992), .ZN(rnd_d[62]) );
  NAND2_X2 U5253 ( .A1(sha1_round_wire[62]), .A2(n7162), .ZN(n5992) );
  NAND2_X2 U5254 ( .A1(n5993), .A2(n5994), .ZN(rnd_d[61]) );
  NAND2_X2 U5255 ( .A1(sha1_round_wire[61]), .A2(n7162), .ZN(n5994) );
  NAND2_X2 U5256 ( .A1(n5995), .A2(n5996), .ZN(rnd_d[60]) );
  NAND2_X2 U5257 ( .A1(sha1_round_wire[60]), .A2(n7162), .ZN(n5996) );
  NAND2_X2 U5258 ( .A1(n5997), .A2(n5998), .ZN(rnd_d[5]) );
  NAND2_X2 U5259 ( .A1(sha1_round_wire[5]), .A2(n7162), .ZN(n5998) );
  NAND2_X2 U5260 ( .A1(n5999), .A2(n6000), .ZN(rnd_d[59]) );
  NAND2_X2 U5261 ( .A1(sha1_round_wire[59]), .A2(n7162), .ZN(n6000) );
  NAND2_X2 U5262 ( .A1(n6001), .A2(n6002), .ZN(rnd_d[58]) );
  NAND2_X2 U5263 ( .A1(sha1_round_wire[58]), .A2(n7162), .ZN(n6002) );
  NAND2_X2 U5264 ( .A1(n6003), .A2(n6004), .ZN(rnd_d[57]) );
  NAND2_X2 U5265 ( .A1(sha1_round_wire[57]), .A2(n7162), .ZN(n6004) );
  NAND2_X2 U5266 ( .A1(n6005), .A2(n6006), .ZN(rnd_d[56]) );
  NAND2_X2 U5267 ( .A1(sha1_round_wire[56]), .A2(n7162), .ZN(n6006) );
  NAND2_X2 U5268 ( .A1(n6007), .A2(n6008), .ZN(rnd_d[55]) );
  NAND2_X2 U5269 ( .A1(sha1_round_wire[55]), .A2(n7162), .ZN(n6008) );
  NAND2_X2 U5270 ( .A1(n6009), .A2(n6010), .ZN(rnd_d[54]) );
  NAND2_X2 U5271 ( .A1(sha1_round_wire[54]), .A2(n7162), .ZN(n6010) );
  NAND2_X2 U5272 ( .A1(n6011), .A2(n6012), .ZN(rnd_d[53]) );
  NAND2_X2 U5273 ( .A1(sha1_round_wire[53]), .A2(n7162), .ZN(n6012) );
  NAND2_X2 U5274 ( .A1(n6013), .A2(n6014), .ZN(rnd_d[52]) );
  NAND2_X2 U5275 ( .A1(sha1_round_wire[52]), .A2(n7162), .ZN(n6014) );
  NAND2_X2 U5276 ( .A1(n6015), .A2(n6016), .ZN(rnd_d[51]) );
  NAND2_X2 U5277 ( .A1(sha1_round_wire[51]), .A2(n7162), .ZN(n6016) );
  NAND2_X2 U5278 ( .A1(n6017), .A2(n6018), .ZN(rnd_d[50]) );
  NAND2_X2 U5279 ( .A1(sha1_round_wire[50]), .A2(n7162), .ZN(n6018) );
  NAND2_X2 U5280 ( .A1(n6019), .A2(n6020), .ZN(rnd_d[4]) );
  NAND2_X2 U5281 ( .A1(sha1_round_wire[4]), .A2(n7162), .ZN(n6020) );
  NAND2_X2 U5282 ( .A1(n6021), .A2(n6022), .ZN(rnd_d[49]) );
  NAND2_X2 U5283 ( .A1(sha1_round_wire[49]), .A2(n7162), .ZN(n6022) );
  NAND2_X2 U5284 ( .A1(n6023), .A2(n6024), .ZN(rnd_d[48]) );
  NAND2_X2 U5285 ( .A1(sha1_round_wire[48]), .A2(n7162), .ZN(n6024) );
  NAND2_X2 U5286 ( .A1(n6025), .A2(n6026), .ZN(rnd_d[47]) );
  NAND2_X2 U5287 ( .A1(sha1_round_wire[47]), .A2(n7162), .ZN(n6026) );
  NAND2_X2 U5288 ( .A1(n6027), .A2(n6028), .ZN(rnd_d[46]) );
  NAND2_X2 U5289 ( .A1(sha1_round_wire[46]), .A2(n7162), .ZN(n6028) );
  NAND2_X2 U5290 ( .A1(n6029), .A2(n6030), .ZN(rnd_d[45]) );
  NAND2_X2 U5291 ( .A1(sha1_round_wire[45]), .A2(n7162), .ZN(n6030) );
  NAND2_X2 U5292 ( .A1(n6031), .A2(n6032), .ZN(rnd_d[44]) );
  NAND2_X2 U5293 ( .A1(sha1_round_wire[44]), .A2(n7163), .ZN(n6032) );
  NAND2_X2 U5294 ( .A1(n6033), .A2(n6034), .ZN(rnd_d[43]) );
  NAND2_X2 U5295 ( .A1(sha1_round_wire[43]), .A2(n7163), .ZN(n6034) );
  NAND2_X2 U5296 ( .A1(n6035), .A2(n6036), .ZN(rnd_d[42]) );
  NAND2_X2 U5297 ( .A1(sha1_round_wire[42]), .A2(n7163), .ZN(n6036) );
  NAND2_X2 U5298 ( .A1(n6037), .A2(n6038), .ZN(rnd_d[41]) );
  NAND2_X2 U5299 ( .A1(sha1_round_wire[41]), .A2(n7163), .ZN(n6038) );
  NAND2_X2 U5300 ( .A1(n6039), .A2(n6040), .ZN(rnd_d[40]) );
  NAND2_X2 U5301 ( .A1(sha1_round_wire[40]), .A2(n7163), .ZN(n6040) );
  NAND2_X2 U5302 ( .A1(n6041), .A2(n6042), .ZN(rnd_d[3]) );
  NAND2_X2 U5303 ( .A1(sha1_round_wire[3]), .A2(n7163), .ZN(n6042) );
  NAND2_X2 U5304 ( .A1(n6043), .A2(n6044), .ZN(rnd_d[39]) );
  NAND2_X2 U5305 ( .A1(sha1_round_wire[39]), .A2(n7163), .ZN(n6044) );
  NAND2_X2 U5306 ( .A1(n6045), .A2(n6046), .ZN(rnd_d[38]) );
  NAND2_X2 U5307 ( .A1(sha1_round_wire[38]), .A2(n7163), .ZN(n6046) );
  NAND2_X2 U5308 ( .A1(n6047), .A2(n6048), .ZN(rnd_d[37]) );
  NAND2_X2 U5309 ( .A1(sha1_round_wire[37]), .A2(n7163), .ZN(n6048) );
  NAND2_X2 U5310 ( .A1(n6049), .A2(n6050), .ZN(rnd_d[36]) );
  NAND2_X2 U5311 ( .A1(sha1_round_wire[36]), .A2(n7163), .ZN(n6050) );
  NAND2_X2 U5312 ( .A1(n6051), .A2(n6052), .ZN(rnd_d[35]) );
  NAND2_X2 U5313 ( .A1(sha1_round_wire[35]), .A2(n7163), .ZN(n6052) );
  NAND2_X2 U5314 ( .A1(n6053), .A2(n6054), .ZN(rnd_d[34]) );
  NAND2_X2 U5315 ( .A1(sha1_round_wire[34]), .A2(n7163), .ZN(n6054) );
  NAND2_X2 U5316 ( .A1(n6055), .A2(n6056), .ZN(rnd_d[33]) );
  NAND2_X2 U5317 ( .A1(sha1_round_wire[33]), .A2(n7163), .ZN(n6056) );
  NAND2_X2 U5318 ( .A1(n6057), .A2(n6058), .ZN(rnd_d[32]) );
  NAND2_X2 U5319 ( .A1(sha1_round_wire[32]), .A2(n7163), .ZN(n6058) );
  NAND2_X2 U5320 ( .A1(n6059), .A2(n6060), .ZN(rnd_d[31]) );
  NAND2_X2 U5321 ( .A1(sha1_round_wire[31]), .A2(n7163), .ZN(n6060) );
  NAND2_X2 U5322 ( .A1(n6061), .A2(n6062), .ZN(rnd_d[30]) );
  NAND2_X2 U5323 ( .A1(sha1_round_wire[30]), .A2(n7163), .ZN(n6062) );
  NAND2_X2 U5324 ( .A1(n6063), .A2(n6064), .ZN(rnd_d[2]) );
  NAND2_X2 U5325 ( .A1(sha1_round_wire[2]), .A2(n7163), .ZN(n6064) );
  NAND2_X2 U5326 ( .A1(n6065), .A2(n6066), .ZN(rnd_d[29]) );
  NAND2_X2 U5327 ( .A1(sha1_round_wire[29]), .A2(n7163), .ZN(n6066) );
  NAND2_X2 U5328 ( .A1(n6067), .A2(n6068), .ZN(rnd_d[28]) );
  NAND2_X2 U5329 ( .A1(sha1_round_wire[28]), .A2(n7163), .ZN(n6068) );
  NAND2_X2 U5330 ( .A1(n6069), .A2(n6070), .ZN(rnd_d[27]) );
  NAND2_X2 U5331 ( .A1(sha1_round_wire[27]), .A2(n7163), .ZN(n6070) );
  NAND2_X2 U5332 ( .A1(n6071), .A2(n6072), .ZN(rnd_d[26]) );
  NAND2_X2 U5333 ( .A1(sha1_round_wire[26]), .A2(n7163), .ZN(n6072) );
  NAND2_X2 U5334 ( .A1(n6073), .A2(n6074), .ZN(rnd_d[25]) );
  NAND2_X2 U5335 ( .A1(sha1_round_wire[25]), .A2(n7163), .ZN(n6074) );
  NAND2_X2 U5336 ( .A1(n6075), .A2(n6076), .ZN(rnd_d[24]) );
  NAND2_X2 U5337 ( .A1(sha1_round_wire[24]), .A2(n7163), .ZN(n6076) );
  NAND2_X2 U5338 ( .A1(n6077), .A2(n6078), .ZN(rnd_d[23]) );
  NAND2_X2 U5339 ( .A1(sha1_round_wire[23]), .A2(n7163), .ZN(n6078) );
  NAND2_X2 U5340 ( .A1(n6079), .A2(n6080), .ZN(rnd_d[22]) );
  NAND2_X2 U5341 ( .A1(sha1_round_wire[22]), .A2(n7163), .ZN(n6080) );
  NAND2_X2 U5342 ( .A1(n6081), .A2(n6082), .ZN(rnd_d[21]) );
  NAND2_X2 U5343 ( .A1(sha1_round_wire[21]), .A2(n7163), .ZN(n6082) );
  NAND2_X2 U5344 ( .A1(n6083), .A2(n6084), .ZN(rnd_d[20]) );
  NAND2_X2 U5345 ( .A1(sha1_round_wire[20]), .A2(n7163), .ZN(n6084) );
  NAND2_X2 U5346 ( .A1(n6085), .A2(n6086), .ZN(rnd_d[1]) );
  NAND2_X2 U5347 ( .A1(sha1_round_wire[1]), .A2(n7164), .ZN(n6086) );
  NAND2_X2 U5348 ( .A1(n6087), .A2(n6088), .ZN(rnd_d[19]) );
  NAND2_X2 U5349 ( .A1(sha1_round_wire[19]), .A2(n7164), .ZN(n6088) );
  NAND2_X2 U5350 ( .A1(n6089), .A2(n6090), .ZN(rnd_d[18]) );
  NAND2_X2 U5351 ( .A1(sha1_round_wire[18]), .A2(n7164), .ZN(n6090) );
  NAND2_X2 U5352 ( .A1(n6091), .A2(n6092), .ZN(rnd_d[17]) );
  NAND2_X2 U5353 ( .A1(sha1_round_wire[17]), .A2(n7164), .ZN(n6092) );
  NAND2_X2 U5354 ( .A1(n6093), .A2(n6094), .ZN(rnd_d[16]) );
  NAND2_X2 U5355 ( .A1(sha1_round_wire[16]), .A2(n7164), .ZN(n6094) );
  NAND2_X2 U5356 ( .A1(n6095), .A2(n6096), .ZN(rnd_d[15]) );
  NAND2_X2 U5357 ( .A1(sha1_round_wire[15]), .A2(n7164), .ZN(n6096) );
  NAND2_X2 U5378 ( .A1(n6117), .A2(n6118), .ZN(rnd_d[14]) );
  NAND2_X2 U5379 ( .A1(sha1_round_wire[14]), .A2(n7164), .ZN(n6118) );
  NAND2_X2 U5400 ( .A1(n6139), .A2(n6140), .ZN(rnd_d[13]) );
  NAND2_X2 U5401 ( .A1(sha1_round_wire[13]), .A2(n7164), .ZN(n6140) );
  NAND2_X2 U5406 ( .A1(n6145), .A2(n6146), .ZN(rnd_d[137]) );
  NAND2_X2 U5407 ( .A1(sha1_round_wire[137]), .A2(n7164), .ZN(n6146) );
  NAND2_X2 U5408 ( .A1(n6147), .A2(n6148), .ZN(rnd_d[136]) );
  NAND2_X2 U5409 ( .A1(sha1_round_wire[136]), .A2(n7164), .ZN(n6148) );
  NAND2_X2 U5410 ( .A1(n6149), .A2(n6150), .ZN(rnd_d[135]) );
  NAND2_X2 U5411 ( .A1(sha1_round_wire[135]), .A2(n7164), .ZN(n6150) );
  NAND2_X2 U5412 ( .A1(n6151), .A2(n6152), .ZN(rnd_d[134]) );
  NAND2_X2 U5413 ( .A1(sha1_round_wire[134]), .A2(n7164), .ZN(n6152) );
  NAND2_X2 U5414 ( .A1(n6153), .A2(n6154), .ZN(rnd_d[133]) );
  NAND2_X2 U5415 ( .A1(sha1_round_wire[133]), .A2(n7164), .ZN(n6154) );
  NAND2_X2 U5416 ( .A1(n6155), .A2(n6156), .ZN(rnd_d[132]) );
  NAND2_X2 U5417 ( .A1(sha1_round_wire[132]), .A2(n7164), .ZN(n6156) );
  NAND2_X2 U5418 ( .A1(n6157), .A2(n6158), .ZN(rnd_d[131]) );
  NAND2_X2 U5419 ( .A1(sha1_round_wire[131]), .A2(n7164), .ZN(n6158) );
  NAND2_X2 U5420 ( .A1(n6159), .A2(n6160), .ZN(rnd_d[130]) );
  NAND2_X2 U5421 ( .A1(sha1_round_wire[130]), .A2(n7164), .ZN(n6160) );
  NAND2_X2 U5422 ( .A1(n6161), .A2(n6162), .ZN(rnd_d[12]) );
  NAND2_X2 U5423 ( .A1(sha1_round_wire[12]), .A2(n7164), .ZN(n6162) );
  NAND2_X2 U5424 ( .A1(n6163), .A2(n6164), .ZN(rnd_d[129]) );
  NAND2_X2 U5425 ( .A1(sha1_round_wire[129]), .A2(n7164), .ZN(n6164) );
  NAND2_X2 U5426 ( .A1(n6165), .A2(n6166), .ZN(rnd_d[128]) );
  NAND2_X2 U5427 ( .A1(sha1_round_wire[128]), .A2(n7164), .ZN(n6166) );
  NAND2_X2 U5428 ( .A1(n6167), .A2(n6168), .ZN(rnd_d[127]) );
  NAND2_X2 U5429 ( .A1(sha1_round_wire[127]), .A2(n7164), .ZN(n6168) );
  NAND2_X2 U5430 ( .A1(n6169), .A2(n6170), .ZN(rnd_d[126]) );
  NAND2_X2 U5431 ( .A1(sha1_round_wire[126]), .A2(n7164), .ZN(n6170) );
  NAND2_X2 U5432 ( .A1(n6171), .A2(n6172), .ZN(rnd_d[125]) );
  NAND2_X2 U5433 ( .A1(sha1_round_wire[125]), .A2(n7164), .ZN(n6172) );
  NAND2_X2 U5434 ( .A1(n6173), .A2(n6174), .ZN(rnd_d[124]) );
  NAND2_X2 U5435 ( .A1(sha1_round_wire[124]), .A2(n7164), .ZN(n6174) );
  NAND2_X2 U5436 ( .A1(n6175), .A2(n6176), .ZN(rnd_d[123]) );
  NAND2_X2 U5437 ( .A1(sha1_round_wire[123]), .A2(n7164), .ZN(n6176) );
  NAND2_X2 U5438 ( .A1(n6177), .A2(n6178), .ZN(rnd_d[122]) );
  NAND2_X2 U5439 ( .A1(sha1_round_wire[122]), .A2(n7164), .ZN(n6178) );
  NAND2_X2 U5440 ( .A1(n6179), .A2(n6180), .ZN(rnd_d[121]) );
  NAND2_X2 U5441 ( .A1(sha1_round_wire[121]), .A2(n7164), .ZN(n6180) );
  NAND2_X2 U5442 ( .A1(n6181), .A2(n6182), .ZN(rnd_d[120]) );
  NAND2_X2 U5443 ( .A1(sha1_round_wire[120]), .A2(n7164), .ZN(n6182) );
  NAND2_X2 U5444 ( .A1(n6183), .A2(n6184), .ZN(rnd_d[11]) );
  NAND2_X2 U5445 ( .A1(sha1_round_wire[11]), .A2(n7165), .ZN(n6184) );
  NAND2_X2 U5446 ( .A1(n6185), .A2(n6186), .ZN(rnd_d[119]) );
  NAND2_X2 U5447 ( .A1(sha1_round_wire[119]), .A2(n7165), .ZN(n6186) );
  NAND2_X2 U5448 ( .A1(n6187), .A2(n6188), .ZN(rnd_d[118]) );
  NAND2_X2 U5449 ( .A1(sha1_round_wire[118]), .A2(n7165), .ZN(n6188) );
  NAND2_X2 U5450 ( .A1(n6189), .A2(n6190), .ZN(rnd_d[117]) );
  NAND2_X2 U5451 ( .A1(sha1_round_wire[117]), .A2(n7165), .ZN(n6190) );
  NAND2_X2 U5452 ( .A1(n6191), .A2(n6192), .ZN(rnd_d[116]) );
  NAND2_X2 U5453 ( .A1(sha1_round_wire[116]), .A2(n7165), .ZN(n6192) );
  NAND2_X2 U5454 ( .A1(n6193), .A2(n6194), .ZN(rnd_d[115]) );
  NAND2_X2 U5455 ( .A1(sha1_round_wire[115]), .A2(n7165), .ZN(n6194) );
  NAND2_X2 U5456 ( .A1(n6195), .A2(n6196), .ZN(rnd_d[114]) );
  NAND2_X2 U5457 ( .A1(sha1_round_wire[114]), .A2(n7165), .ZN(n6196) );
  NAND2_X2 U5458 ( .A1(n6197), .A2(n6198), .ZN(rnd_d[113]) );
  NAND2_X2 U5459 ( .A1(sha1_round_wire[113]), .A2(n7155), .ZN(n6198) );
  NAND2_X2 U5460 ( .A1(n6199), .A2(n6200), .ZN(rnd_d[112]) );
  NAND2_X2 U5461 ( .A1(sha1_round_wire[112]), .A2(n7152), .ZN(n6200) );
  NAND2_X2 U5462 ( .A1(n6201), .A2(n6202), .ZN(rnd_d[111]) );
  NAND2_X2 U5463 ( .A1(sha1_round_wire[111]), .A2(n7152), .ZN(n6202) );
  NAND2_X2 U5464 ( .A1(n6203), .A2(n6204), .ZN(rnd_d[110]) );
  NAND2_X2 U5465 ( .A1(sha1_round_wire[110]), .A2(n7152), .ZN(n6204) );
  NAND2_X2 U5466 ( .A1(n6205), .A2(n6206), .ZN(rnd_d[10]) );
  NAND2_X2 U5467 ( .A1(sha1_round_wire[10]), .A2(n7152), .ZN(n6206) );
  NAND2_X2 U5468 ( .A1(n6207), .A2(n6208), .ZN(rnd_d[109]) );
  NAND2_X2 U5469 ( .A1(sha1_round_wire[109]), .A2(n7152), .ZN(n6208) );
  NAND2_X2 U5470 ( .A1(n6209), .A2(n6210), .ZN(rnd_d[108]) );
  NAND2_X2 U5471 ( .A1(sha1_round_wire[108]), .A2(n7152), .ZN(n6210) );
  NAND2_X2 U5472 ( .A1(n6211), .A2(n6212), .ZN(rnd_d[107]) );
  NAND2_X2 U5473 ( .A1(sha1_round_wire[107]), .A2(n7152), .ZN(n6212) );
  NAND2_X2 U5474 ( .A1(n6213), .A2(n6214), .ZN(rnd_d[106]) );
  NAND2_X2 U5475 ( .A1(sha1_round_wire[106]), .A2(n7152), .ZN(n6214) );
  NAND2_X2 U5476 ( .A1(n6215), .A2(n6216), .ZN(rnd_d[105]) );
  NAND2_X2 U5477 ( .A1(sha1_round_wire[105]), .A2(n7152), .ZN(n6216) );
  NAND2_X2 U5478 ( .A1(n6217), .A2(n6218), .ZN(rnd_d[104]) );
  NAND2_X2 U5479 ( .A1(sha1_round_wire[104]), .A2(n7152), .ZN(n6218) );
  NAND2_X2 U5480 ( .A1(n6219), .A2(n6220), .ZN(rnd_d[103]) );
  NAND2_X2 U5481 ( .A1(sha1_round_wire[103]), .A2(n7152), .ZN(n6220) );
  NAND2_X2 U5482 ( .A1(n6221), .A2(n6222), .ZN(rnd_d[102]) );
  NAND2_X2 U5483 ( .A1(sha1_round_wire[102]), .A2(n7152), .ZN(n6222) );
  NAND2_X2 U5484 ( .A1(n6223), .A2(n6224), .ZN(rnd_d[101]) );
  NAND2_X2 U5485 ( .A1(sha1_round_wire[101]), .A2(n7152), .ZN(n6224) );
  NAND2_X2 U5486 ( .A1(n6225), .A2(n6226), .ZN(rnd_d[100]) );
  NAND2_X2 U5487 ( .A1(sha1_round_wire[100]), .A2(n7152), .ZN(n6226) );
  NAND2_X2 U5488 ( .A1(n6227), .A2(n6228), .ZN(rnd_d[0]) );
  NAND2_X2 U5489 ( .A1(sha1_round_wire[0]), .A2(n7152), .ZN(n6228) );
  XNOR2_X2 U5494 ( .A(n6232), .B(n7398), .ZN(n6233) );
  NAND2_X2 U5500 ( .A1(n6237), .A2(n6238), .ZN(rnd_cnt_d[2]) );
  NAND4_X2 U5501 ( .A1(n7396), .A2(rnd_cnt_q[1]), .A3(rnd_cnt_q[0]), .A4(n7400), .ZN(n6238) );
  NAND2_X2 U5503 ( .A1(n7397), .A2(n6240), .ZN(n6239) );
  NAND2_X2 U5504 ( .A1(n7396), .A2(n7401), .ZN(n6240) );
  NAND2_X2 U5505 ( .A1(n6241), .A2(n6242), .ZN(rnd_cnt_d[1]) );
  NAND2_X2 U5507 ( .A1(rnd_cnt_d[0]), .A2(rnd_cnt_q[1]), .ZN(n6241) );
  AND2_X2 U5509 ( .A1(state[0]), .A2(state[1]), .ZN(out_valid) );
  NAND2_X2 U5514 ( .A1(n7176), .A2(n7402), .ZN(n6247) );
  AND2_X2 U5517 ( .A1(rnd_cnt_q[3]), .A2(n6236), .ZN(n5038) );
  NAND2_X2 U6001 ( .A1(n5909), .A2(n6569), .ZN(cv_d[9]) );
  NAND2_X2 U6002 ( .A1(cv_q[9]), .A2(n7152), .ZN(n6569) );
  NAND2_X2 U6004 ( .A1(cv[9]), .A2(n7124), .ZN(n6571) );
  NAND2_X2 U6005 ( .A1(cv_next[9]), .A2(n7139), .ZN(n6570) );
  NAND2_X2 U6006 ( .A1(n5911), .A2(n6574), .ZN(cv_d[99]) );
  NAND2_X2 U6007 ( .A1(cv_q[99]), .A2(n7152), .ZN(n6574) );
  NAND2_X2 U6009 ( .A1(cv[99]), .A2(n7124), .ZN(n6576) );
  NAND2_X2 U6010 ( .A1(cv_next[99]), .A2(n7139), .ZN(n6575) );
  NAND2_X2 U6011 ( .A1(n5913), .A2(n6577), .ZN(cv_d[98]) );
  NAND2_X2 U6012 ( .A1(cv_q[98]), .A2(n7152), .ZN(n6577) );
  NAND2_X2 U6014 ( .A1(cv[98]), .A2(n7124), .ZN(n6579) );
  NAND2_X2 U6015 ( .A1(cv_next[98]), .A2(n7139), .ZN(n6578) );
  NAND2_X2 U6016 ( .A1(n5915), .A2(n6580), .ZN(cv_d[97]) );
  NAND2_X2 U6017 ( .A1(cv_q[97]), .A2(n7153), .ZN(n6580) );
  NAND2_X2 U6019 ( .A1(cv[97]), .A2(n7124), .ZN(n6582) );
  NAND2_X2 U6020 ( .A1(cv_next[97]), .A2(n7139), .ZN(n6581) );
  NAND2_X2 U6021 ( .A1(n5917), .A2(n6583), .ZN(cv_d[96]) );
  NAND2_X2 U6022 ( .A1(cv_q[96]), .A2(n7152), .ZN(n6583) );
  NAND2_X2 U6024 ( .A1(cv[96]), .A2(n7124), .ZN(n6585) );
  NAND2_X2 U6025 ( .A1(cv_next[96]), .A2(n7139), .ZN(n6584) );
  NAND2_X2 U6026 ( .A1(n5919), .A2(n6586), .ZN(cv_d[95]) );
  NAND2_X2 U6027 ( .A1(cv_q[95]), .A2(n7152), .ZN(n6586) );
  NAND2_X2 U6029 ( .A1(cv[95]), .A2(n7124), .ZN(n6588) );
  NAND2_X2 U6030 ( .A1(cv_next[95]), .A2(n7139), .ZN(n6587) );
  NAND2_X2 U6031 ( .A1(n5921), .A2(n6589), .ZN(cv_d[94]) );
  NAND2_X2 U6032 ( .A1(cv_q[94]), .A2(n7153), .ZN(n6589) );
  NAND2_X2 U6034 ( .A1(cv[94]), .A2(n7124), .ZN(n6591) );
  NAND2_X2 U6035 ( .A1(cv_next[94]), .A2(n7139), .ZN(n6590) );
  NAND2_X2 U6036 ( .A1(n5923), .A2(n6592), .ZN(cv_d[93]) );
  NAND2_X2 U6037 ( .A1(cv_q[93]), .A2(n7153), .ZN(n6592) );
  NAND2_X2 U6039 ( .A1(cv[93]), .A2(n7124), .ZN(n6594) );
  NAND2_X2 U6040 ( .A1(cv_next[93]), .A2(n7139), .ZN(n6593) );
  NAND2_X2 U6041 ( .A1(n5925), .A2(n6595), .ZN(cv_d[92]) );
  NAND2_X2 U6042 ( .A1(cv_q[92]), .A2(n7153), .ZN(n6595) );
  NAND2_X2 U6044 ( .A1(cv[92]), .A2(n7124), .ZN(n6597) );
  NAND2_X2 U6045 ( .A1(cv_next[92]), .A2(n7139), .ZN(n6596) );
  NAND2_X2 U6046 ( .A1(n5927), .A2(n6598), .ZN(cv_d[91]) );
  NAND2_X2 U6047 ( .A1(cv_q[91]), .A2(n7153), .ZN(n6598) );
  NAND2_X2 U6049 ( .A1(cv[91]), .A2(n7124), .ZN(n6600) );
  NAND2_X2 U6050 ( .A1(cv_next[91]), .A2(n7139), .ZN(n6599) );
  NAND2_X2 U6051 ( .A1(n5929), .A2(n6601), .ZN(cv_d[90]) );
  NAND2_X2 U6052 ( .A1(cv_q[90]), .A2(n7153), .ZN(n6601) );
  NAND2_X2 U6054 ( .A1(cv[90]), .A2(n7124), .ZN(n6603) );
  NAND2_X2 U6055 ( .A1(cv_next[90]), .A2(n7139), .ZN(n6602) );
  NAND2_X2 U6056 ( .A1(n5931), .A2(n6604), .ZN(cv_d[8]) );
  NAND2_X2 U6057 ( .A1(cv_q[8]), .A2(n7153), .ZN(n6604) );
  NAND2_X2 U6059 ( .A1(cv[8]), .A2(n7125), .ZN(n6606) );
  NAND2_X2 U6060 ( .A1(cv_next[8]), .A2(n7140), .ZN(n6605) );
  NAND2_X2 U6061 ( .A1(n5933), .A2(n6607), .ZN(cv_d[89]) );
  NAND2_X2 U6062 ( .A1(cv_q[89]), .A2(n7153), .ZN(n6607) );
  NAND2_X2 U6064 ( .A1(cv[89]), .A2(n7125), .ZN(n6609) );
  NAND2_X2 U6065 ( .A1(cv_next[89]), .A2(n7140), .ZN(n6608) );
  NAND2_X2 U6066 ( .A1(n5935), .A2(n6610), .ZN(cv_d[88]) );
  NAND2_X2 U6067 ( .A1(cv_q[88]), .A2(n7153), .ZN(n6610) );
  NAND2_X2 U6069 ( .A1(cv[88]), .A2(n7125), .ZN(n6612) );
  NAND2_X2 U6070 ( .A1(cv_next[88]), .A2(n7140), .ZN(n6611) );
  NAND2_X2 U6071 ( .A1(n5937), .A2(n6613), .ZN(cv_d[87]) );
  NAND2_X2 U6072 ( .A1(cv_q[87]), .A2(n7153), .ZN(n6613) );
  NAND2_X2 U6074 ( .A1(cv[87]), .A2(n7125), .ZN(n6615) );
  NAND2_X2 U6075 ( .A1(cv_next[87]), .A2(n7140), .ZN(n6614) );
  NAND2_X2 U6076 ( .A1(n5939), .A2(n6616), .ZN(cv_d[86]) );
  NAND2_X2 U6077 ( .A1(cv_q[86]), .A2(n7153), .ZN(n6616) );
  NAND2_X2 U6079 ( .A1(cv[86]), .A2(n7125), .ZN(n6618) );
  NAND2_X2 U6080 ( .A1(cv_next[86]), .A2(n7140), .ZN(n6617) );
  NAND2_X2 U6081 ( .A1(n5941), .A2(n6619), .ZN(cv_d[85]) );
  NAND2_X2 U6082 ( .A1(cv_q[85]), .A2(n7153), .ZN(n6619) );
  NAND2_X2 U6084 ( .A1(cv[85]), .A2(n7125), .ZN(n6621) );
  NAND2_X2 U6085 ( .A1(cv_next[85]), .A2(n7140), .ZN(n6620) );
  NAND2_X2 U6086 ( .A1(n5943), .A2(n6622), .ZN(cv_d[84]) );
  NAND2_X2 U6087 ( .A1(cv_q[84]), .A2(n7153), .ZN(n6622) );
  NAND2_X2 U6089 ( .A1(cv[84]), .A2(n7125), .ZN(n6624) );
  NAND2_X2 U6090 ( .A1(cv_next[84]), .A2(n7140), .ZN(n6623) );
  NAND2_X2 U6091 ( .A1(n5945), .A2(n6625), .ZN(cv_d[83]) );
  NAND2_X2 U6092 ( .A1(cv_q[83]), .A2(n7153), .ZN(n6625) );
  NAND2_X2 U6094 ( .A1(cv[83]), .A2(n7125), .ZN(n6627) );
  NAND2_X2 U6095 ( .A1(cv_next[83]), .A2(n7140), .ZN(n6626) );
  NAND2_X2 U6096 ( .A1(n5947), .A2(n6628), .ZN(cv_d[82]) );
  NAND2_X2 U6097 ( .A1(cv_q[82]), .A2(n7153), .ZN(n6628) );
  NAND2_X2 U6099 ( .A1(cv[82]), .A2(n7125), .ZN(n6630) );
  NAND2_X2 U6100 ( .A1(cv_next[82]), .A2(n7140), .ZN(n6629) );
  NAND2_X2 U6101 ( .A1(n5949), .A2(n6631), .ZN(cv_d[81]) );
  NAND2_X2 U6102 ( .A1(cv_q[81]), .A2(n7153), .ZN(n6631) );
  NAND2_X2 U6104 ( .A1(cv[81]), .A2(n7125), .ZN(n6633) );
  NAND2_X2 U6105 ( .A1(cv_next[81]), .A2(n7140), .ZN(n6632) );
  NAND2_X2 U6106 ( .A1(n5951), .A2(n6634), .ZN(cv_d[80]) );
  NAND2_X2 U6107 ( .A1(cv_q[80]), .A2(n7153), .ZN(n6634) );
  NAND2_X2 U6109 ( .A1(cv[80]), .A2(n7125), .ZN(n6636) );
  NAND2_X2 U6110 ( .A1(cv_next[80]), .A2(n7140), .ZN(n6635) );
  NAND2_X2 U6111 ( .A1(n5953), .A2(n6637), .ZN(cv_d[7]) );
  NAND2_X2 U6112 ( .A1(cv_q[7]), .A2(n7153), .ZN(n6637) );
  NAND2_X2 U6114 ( .A1(cv[7]), .A2(n7126), .ZN(n6639) );
  NAND2_X2 U6115 ( .A1(cv_next[7]), .A2(n7141), .ZN(n6638) );
  NAND2_X2 U6116 ( .A1(n5955), .A2(n6640), .ZN(cv_d[79]) );
  NAND2_X2 U6117 ( .A1(cv_q[79]), .A2(n7153), .ZN(n6640) );
  NAND2_X2 U6119 ( .A1(cv[79]), .A2(n7126), .ZN(n6642) );
  NAND2_X2 U6120 ( .A1(cv_next[79]), .A2(n7141), .ZN(n6641) );
  NAND2_X2 U6121 ( .A1(n5957), .A2(n6643), .ZN(cv_d[78]) );
  NAND2_X2 U6122 ( .A1(cv_q[78]), .A2(n7153), .ZN(n6643) );
  NAND2_X2 U6124 ( .A1(cv[78]), .A2(n7126), .ZN(n6645) );
  NAND2_X2 U6125 ( .A1(cv_next[78]), .A2(n7141), .ZN(n6644) );
  NAND2_X2 U6126 ( .A1(n5959), .A2(n6646), .ZN(cv_d[77]) );
  NAND2_X2 U6127 ( .A1(cv_q[77]), .A2(n7153), .ZN(n6646) );
  NAND2_X2 U6129 ( .A1(cv[77]), .A2(n7126), .ZN(n6648) );
  NAND2_X2 U6130 ( .A1(cv_next[77]), .A2(n7141), .ZN(n6647) );
  NAND2_X2 U6131 ( .A1(n5961), .A2(n6649), .ZN(cv_d[76]) );
  NAND2_X2 U6132 ( .A1(cv_q[76]), .A2(n7153), .ZN(n6649) );
  NAND2_X2 U6134 ( .A1(cv[76]), .A2(n7126), .ZN(n6651) );
  NAND2_X2 U6135 ( .A1(cv_next[76]), .A2(n7141), .ZN(n6650) );
  NAND2_X2 U6136 ( .A1(n5963), .A2(n6652), .ZN(cv_d[75]) );
  NAND2_X2 U6137 ( .A1(cv_q[75]), .A2(n7153), .ZN(n6652) );
  NAND2_X2 U6139 ( .A1(cv[75]), .A2(n7126), .ZN(n6654) );
  NAND2_X2 U6140 ( .A1(cv_next[75]), .A2(n7141), .ZN(n6653) );
  NAND2_X2 U6141 ( .A1(n5965), .A2(n6655), .ZN(cv_d[74]) );
  NAND2_X2 U6142 ( .A1(cv_q[74]), .A2(n7153), .ZN(n6655) );
  NAND2_X2 U6144 ( .A1(cv[74]), .A2(n7126), .ZN(n6657) );
  NAND2_X2 U6145 ( .A1(cv_next[74]), .A2(n7141), .ZN(n6656) );
  NAND2_X2 U6146 ( .A1(n5967), .A2(n6658), .ZN(cv_d[73]) );
  NAND2_X2 U6147 ( .A1(cv_q[73]), .A2(n7153), .ZN(n6658) );
  NAND2_X2 U6149 ( .A1(cv[73]), .A2(n7126), .ZN(n6660) );
  NAND2_X2 U6150 ( .A1(cv_next[73]), .A2(n7141), .ZN(n6659) );
  NAND2_X2 U6151 ( .A1(n5969), .A2(n6661), .ZN(cv_d[72]) );
  NAND2_X2 U6152 ( .A1(cv_q[72]), .A2(n7154), .ZN(n6661) );
  NAND2_X2 U6154 ( .A1(cv[72]), .A2(n7126), .ZN(n6663) );
  NAND2_X2 U6155 ( .A1(cv_next[72]), .A2(n7141), .ZN(n6662) );
  NAND2_X2 U6156 ( .A1(n5971), .A2(n6664), .ZN(cv_d[71]) );
  NAND2_X2 U6157 ( .A1(cv_q[71]), .A2(n7153), .ZN(n6664) );
  NAND2_X2 U6159 ( .A1(cv[71]), .A2(n7126), .ZN(n6666) );
  NAND2_X2 U6160 ( .A1(cv_next[71]), .A2(n7141), .ZN(n6665) );
  NAND2_X2 U6161 ( .A1(n5973), .A2(n6667), .ZN(cv_d[70]) );
  NAND2_X2 U6162 ( .A1(cv_q[70]), .A2(n7153), .ZN(n6667) );
  NAND2_X2 U6164 ( .A1(cv[70]), .A2(n7126), .ZN(n6669) );
  NAND2_X2 U6165 ( .A1(cv_next[70]), .A2(n7141), .ZN(n6668) );
  NAND2_X2 U6166 ( .A1(n5975), .A2(n6670), .ZN(cv_d[6]) );
  NAND2_X2 U6167 ( .A1(cv_q[6]), .A2(n7154), .ZN(n6670) );
  NAND2_X2 U6169 ( .A1(cv[6]), .A2(n7127), .ZN(n6672) );
  NAND2_X2 U6170 ( .A1(cv_next[6]), .A2(n7142), .ZN(n6671) );
  NAND2_X2 U6171 ( .A1(n5977), .A2(n6673), .ZN(cv_d[69]) );
  NAND2_X2 U6172 ( .A1(cv_q[69]), .A2(n7154), .ZN(n6673) );
  NAND2_X2 U6174 ( .A1(cv[69]), .A2(n7127), .ZN(n6675) );
  NAND2_X2 U6175 ( .A1(cv_next[69]), .A2(n7142), .ZN(n6674) );
  NAND2_X2 U6176 ( .A1(n5979), .A2(n6676), .ZN(cv_d[68]) );
  NAND2_X2 U6177 ( .A1(cv_q[68]), .A2(n7154), .ZN(n6676) );
  NAND2_X2 U6179 ( .A1(cv[68]), .A2(n7127), .ZN(n6678) );
  NAND2_X2 U6180 ( .A1(cv_next[68]), .A2(n7142), .ZN(n6677) );
  NAND2_X2 U6181 ( .A1(n5981), .A2(n6679), .ZN(cv_d[67]) );
  NAND2_X2 U6182 ( .A1(cv_q[67]), .A2(n7154), .ZN(n6679) );
  NAND2_X2 U6184 ( .A1(cv[67]), .A2(n7127), .ZN(n6681) );
  NAND2_X2 U6185 ( .A1(cv_next[67]), .A2(n7142), .ZN(n6680) );
  NAND2_X2 U6186 ( .A1(n5983), .A2(n6682), .ZN(cv_d[66]) );
  NAND2_X2 U6187 ( .A1(cv_q[66]), .A2(n7154), .ZN(n6682) );
  NAND2_X2 U6189 ( .A1(cv[66]), .A2(n7127), .ZN(n6684) );
  NAND2_X2 U6190 ( .A1(cv_next[66]), .A2(n7142), .ZN(n6683) );
  NAND2_X2 U6191 ( .A1(n5985), .A2(n6685), .ZN(cv_d[65]) );
  NAND2_X2 U6192 ( .A1(cv_q[65]), .A2(n7154), .ZN(n6685) );
  NAND2_X2 U6194 ( .A1(cv[65]), .A2(n7127), .ZN(n6687) );
  NAND2_X2 U6195 ( .A1(cv_next[65]), .A2(n7142), .ZN(n6686) );
  NAND2_X2 U6196 ( .A1(n5987), .A2(n6688), .ZN(cv_d[64]) );
  NAND2_X2 U6197 ( .A1(cv_q[64]), .A2(n7154), .ZN(n6688) );
  NAND2_X2 U6199 ( .A1(cv[64]), .A2(n7127), .ZN(n6690) );
  NAND2_X2 U6200 ( .A1(cv_next[64]), .A2(n7142), .ZN(n6689) );
  NAND2_X2 U6201 ( .A1(n5989), .A2(n6691), .ZN(cv_d[63]) );
  NAND2_X2 U6202 ( .A1(cv_q[63]), .A2(n7154), .ZN(n6691) );
  NAND2_X2 U6204 ( .A1(cv[63]), .A2(n7127), .ZN(n6693) );
  NAND2_X2 U6205 ( .A1(cv_next[63]), .A2(n7142), .ZN(n6692) );
  NAND2_X2 U6206 ( .A1(n5991), .A2(n6694), .ZN(cv_d[62]) );
  NAND2_X2 U6207 ( .A1(cv_q[62]), .A2(n7154), .ZN(n6694) );
  NAND2_X2 U6209 ( .A1(cv[62]), .A2(n7127), .ZN(n6696) );
  NAND2_X2 U6210 ( .A1(cv_next[62]), .A2(n7142), .ZN(n6695) );
  NAND2_X2 U6211 ( .A1(n5993), .A2(n6697), .ZN(cv_d[61]) );
  NAND2_X2 U6212 ( .A1(cv_q[61]), .A2(n7154), .ZN(n6697) );
  NAND2_X2 U6214 ( .A1(cv[61]), .A2(n7127), .ZN(n6699) );
  NAND2_X2 U6215 ( .A1(cv_next[61]), .A2(n7142), .ZN(n6698) );
  NAND2_X2 U6216 ( .A1(n5995), .A2(n6700), .ZN(cv_d[60]) );
  NAND2_X2 U6217 ( .A1(cv_q[60]), .A2(n7154), .ZN(n6700) );
  NAND2_X2 U6219 ( .A1(cv[60]), .A2(n7127), .ZN(n6702) );
  NAND2_X2 U6220 ( .A1(cv_next[60]), .A2(n7142), .ZN(n6701) );
  NAND2_X2 U6221 ( .A1(n5997), .A2(n6703), .ZN(cv_d[5]) );
  NAND2_X2 U6222 ( .A1(cv_q[5]), .A2(n7154), .ZN(n6703) );
  NAND2_X2 U6224 ( .A1(cv[5]), .A2(n7128), .ZN(n6705) );
  NAND2_X2 U6225 ( .A1(cv_next[5]), .A2(n7143), .ZN(n6704) );
  NAND2_X2 U6226 ( .A1(n5999), .A2(n6706), .ZN(cv_d[59]) );
  NAND2_X2 U6227 ( .A1(cv_q[59]), .A2(n7154), .ZN(n6706) );
  NAND2_X2 U6229 ( .A1(cv[59]), .A2(n7128), .ZN(n6708) );
  NAND2_X2 U6230 ( .A1(cv_next[59]), .A2(n7143), .ZN(n6707) );
  NAND2_X2 U6231 ( .A1(n6001), .A2(n6709), .ZN(cv_d[58]) );
  NAND2_X2 U6232 ( .A1(cv_q[58]), .A2(n7154), .ZN(n6709) );
  NAND2_X2 U6234 ( .A1(cv[58]), .A2(n7128), .ZN(n6711) );
  NAND2_X2 U6235 ( .A1(cv_next[58]), .A2(n7143), .ZN(n6710) );
  NAND2_X2 U6236 ( .A1(n6003), .A2(n6712), .ZN(cv_d[57]) );
  NAND2_X2 U6237 ( .A1(cv_q[57]), .A2(n7154), .ZN(n6712) );
  NAND2_X2 U6239 ( .A1(cv[57]), .A2(n7128), .ZN(n6714) );
  NAND2_X2 U6240 ( .A1(cv_next[57]), .A2(n7143), .ZN(n6713) );
  NAND2_X2 U6241 ( .A1(n6005), .A2(n6715), .ZN(cv_d[56]) );
  NAND2_X2 U6242 ( .A1(cv_q[56]), .A2(n7154), .ZN(n6715) );
  NAND2_X2 U6244 ( .A1(cv[56]), .A2(n7128), .ZN(n6717) );
  NAND2_X2 U6245 ( .A1(cv_next[56]), .A2(n7143), .ZN(n6716) );
  NAND2_X2 U6246 ( .A1(n6007), .A2(n6718), .ZN(cv_d[55]) );
  NAND2_X2 U6247 ( .A1(cv_q[55]), .A2(n7154), .ZN(n6718) );
  NAND2_X2 U6249 ( .A1(cv[55]), .A2(n7128), .ZN(n6720) );
  NAND2_X2 U6250 ( .A1(cv_next[55]), .A2(n7143), .ZN(n6719) );
  NAND2_X2 U6251 ( .A1(n6009), .A2(n6721), .ZN(cv_d[54]) );
  NAND2_X2 U6252 ( .A1(cv_q[54]), .A2(n7154), .ZN(n6721) );
  NAND2_X2 U6254 ( .A1(cv[54]), .A2(n7128), .ZN(n6723) );
  NAND2_X2 U6255 ( .A1(cv_next[54]), .A2(n7143), .ZN(n6722) );
  NAND2_X2 U6256 ( .A1(n6011), .A2(n6724), .ZN(cv_d[53]) );
  NAND2_X2 U6257 ( .A1(cv_q[53]), .A2(n7154), .ZN(n6724) );
  NAND2_X2 U6259 ( .A1(cv[53]), .A2(n7128), .ZN(n6726) );
  NAND2_X2 U6260 ( .A1(cv_next[53]), .A2(n7143), .ZN(n6725) );
  NAND2_X2 U6261 ( .A1(n6013), .A2(n6727), .ZN(cv_d[52]) );
  NAND2_X2 U6262 ( .A1(cv_q[52]), .A2(n7154), .ZN(n6727) );
  NAND2_X2 U6264 ( .A1(cv[52]), .A2(n7128), .ZN(n6729) );
  NAND2_X2 U6265 ( .A1(cv_next[52]), .A2(n7143), .ZN(n6728) );
  NAND2_X2 U6266 ( .A1(n6015), .A2(n6730), .ZN(cv_d[51]) );
  NAND2_X2 U6267 ( .A1(cv_q[51]), .A2(n7154), .ZN(n6730) );
  NAND2_X2 U6269 ( .A1(cv[51]), .A2(n7128), .ZN(n6732) );
  NAND2_X2 U6270 ( .A1(cv_next[51]), .A2(n7143), .ZN(n6731) );
  NAND2_X2 U6271 ( .A1(n6017), .A2(n6733), .ZN(cv_d[50]) );
  NAND2_X2 U6272 ( .A1(cv_q[50]), .A2(n7154), .ZN(n6733) );
  NAND2_X2 U6274 ( .A1(cv[50]), .A2(n7128), .ZN(n6735) );
  NAND2_X2 U6275 ( .A1(cv_next[50]), .A2(n7143), .ZN(n6734) );
  NAND2_X2 U6276 ( .A1(n6019), .A2(n6736), .ZN(cv_d[4]) );
  NAND2_X2 U6277 ( .A1(cv_q[4]), .A2(n7154), .ZN(n6736) );
  NAND2_X2 U6279 ( .A1(cv[4]), .A2(n7129), .ZN(n6738) );
  NAND2_X2 U6280 ( .A1(cv_next[4]), .A2(n7144), .ZN(n6737) );
  NAND2_X2 U6281 ( .A1(n6021), .A2(n6739), .ZN(cv_d[49]) );
  NAND2_X2 U6282 ( .A1(cv_q[49]), .A2(n7154), .ZN(n6739) );
  NAND2_X2 U6284 ( .A1(cv[49]), .A2(n7129), .ZN(n6741) );
  NAND2_X2 U6285 ( .A1(cv_next[49]), .A2(n7144), .ZN(n6740) );
  NAND2_X2 U6286 ( .A1(n6023), .A2(n6742), .ZN(cv_d[48]) );
  NAND2_X2 U6287 ( .A1(cv_q[48]), .A2(n7154), .ZN(n6742) );
  NAND2_X2 U6289 ( .A1(cv[48]), .A2(n7129), .ZN(n6744) );
  NAND2_X2 U6290 ( .A1(cv_next[48]), .A2(n7144), .ZN(n6743) );
  NAND2_X2 U6291 ( .A1(n6025), .A2(n6745), .ZN(cv_d[47]) );
  NAND2_X2 U6292 ( .A1(cv_q[47]), .A2(n7154), .ZN(n6745) );
  NAND2_X2 U6294 ( .A1(cv[47]), .A2(n7129), .ZN(n6747) );
  NAND2_X2 U6295 ( .A1(cv_next[47]), .A2(n7144), .ZN(n6746) );
  NAND2_X2 U6296 ( .A1(n6027), .A2(n6748), .ZN(cv_d[46]) );
  NAND2_X2 U6297 ( .A1(cv_q[46]), .A2(n7155), .ZN(n6748) );
  NAND2_X2 U6299 ( .A1(cv[46]), .A2(n7129), .ZN(n6750) );
  NAND2_X2 U6300 ( .A1(cv_next[46]), .A2(n7144), .ZN(n6749) );
  NAND2_X2 U6301 ( .A1(n6029), .A2(n6751), .ZN(cv_d[45]) );
  NAND2_X2 U6302 ( .A1(cv_q[45]), .A2(n7155), .ZN(n6751) );
  NAND2_X2 U6304 ( .A1(cv[45]), .A2(n7129), .ZN(n6753) );
  NAND2_X2 U6305 ( .A1(cv_next[45]), .A2(n7144), .ZN(n6752) );
  NAND2_X2 U6306 ( .A1(n6031), .A2(n6754), .ZN(cv_d[44]) );
  NAND2_X2 U6307 ( .A1(cv_q[44]), .A2(n7155), .ZN(n6754) );
  NAND2_X2 U6309 ( .A1(cv[44]), .A2(n7129), .ZN(n6756) );
  NAND2_X2 U6310 ( .A1(cv_next[44]), .A2(n7144), .ZN(n6755) );
  NAND2_X2 U6311 ( .A1(n6033), .A2(n6757), .ZN(cv_d[43]) );
  NAND2_X2 U6312 ( .A1(cv_q[43]), .A2(n7155), .ZN(n6757) );
  NAND2_X2 U6314 ( .A1(cv[43]), .A2(n7129), .ZN(n6759) );
  NAND2_X2 U6315 ( .A1(cv_next[43]), .A2(n7144), .ZN(n6758) );
  NAND2_X2 U6316 ( .A1(n6035), .A2(n6760), .ZN(cv_d[42]) );
  NAND2_X2 U6317 ( .A1(cv_q[42]), .A2(n7155), .ZN(n6760) );
  NAND2_X2 U6319 ( .A1(cv[42]), .A2(n7129), .ZN(n6762) );
  NAND2_X2 U6320 ( .A1(cv_next[42]), .A2(n7144), .ZN(n6761) );
  NAND2_X2 U6321 ( .A1(n6037), .A2(n6763), .ZN(cv_d[41]) );
  NAND2_X2 U6322 ( .A1(cv_q[41]), .A2(n7155), .ZN(n6763) );
  NAND2_X2 U6324 ( .A1(cv[41]), .A2(n7129), .ZN(n6765) );
  NAND2_X2 U6325 ( .A1(cv_next[41]), .A2(n7144), .ZN(n6764) );
  NAND2_X2 U6326 ( .A1(n6039), .A2(n6766), .ZN(cv_d[40]) );
  NAND2_X2 U6327 ( .A1(cv_q[40]), .A2(n7155), .ZN(n6766) );
  NAND2_X2 U6329 ( .A1(cv[40]), .A2(n7129), .ZN(n6768) );
  NAND2_X2 U6330 ( .A1(cv_next[40]), .A2(n7144), .ZN(n6767) );
  NAND2_X2 U6331 ( .A1(n6041), .A2(n6769), .ZN(cv_d[3]) );
  NAND2_X2 U6332 ( .A1(cv_q[3]), .A2(n7155), .ZN(n6769) );
  NAND2_X2 U6334 ( .A1(cv[3]), .A2(n7130), .ZN(n6771) );
  NAND2_X2 U6335 ( .A1(cv_next[3]), .A2(n7145), .ZN(n6770) );
  NAND2_X2 U6336 ( .A1(n6043), .A2(n6772), .ZN(cv_d[39]) );
  NAND2_X2 U6337 ( .A1(cv_q[39]), .A2(n7155), .ZN(n6772) );
  NAND2_X2 U6339 ( .A1(cv[39]), .A2(n7130), .ZN(n6774) );
  NAND2_X2 U6340 ( .A1(cv_next[39]), .A2(n7145), .ZN(n6773) );
  NAND2_X2 U6341 ( .A1(n6045), .A2(n6775), .ZN(cv_d[38]) );
  NAND2_X2 U6342 ( .A1(cv_q[38]), .A2(n7155), .ZN(n6775) );
  NAND2_X2 U6344 ( .A1(cv[38]), .A2(n7130), .ZN(n6777) );
  NAND2_X2 U6345 ( .A1(cv_next[38]), .A2(n7145), .ZN(n6776) );
  NAND2_X2 U6346 ( .A1(n6047), .A2(n6778), .ZN(cv_d[37]) );
  NAND2_X2 U6347 ( .A1(cv_q[37]), .A2(n7155), .ZN(n6778) );
  NAND2_X2 U6349 ( .A1(cv[37]), .A2(n7130), .ZN(n6780) );
  NAND2_X2 U6350 ( .A1(cv_next[37]), .A2(n7145), .ZN(n6779) );
  NAND2_X2 U6351 ( .A1(n6049), .A2(n6781), .ZN(cv_d[36]) );
  NAND2_X2 U6352 ( .A1(cv_q[36]), .A2(n7155), .ZN(n6781) );
  NAND2_X2 U6354 ( .A1(cv[36]), .A2(n7130), .ZN(n6783) );
  NAND2_X2 U6355 ( .A1(cv_next[36]), .A2(n7145), .ZN(n6782) );
  NAND2_X2 U6356 ( .A1(n6051), .A2(n6784), .ZN(cv_d[35]) );
  NAND2_X2 U6357 ( .A1(cv_q[35]), .A2(n7155), .ZN(n6784) );
  NAND2_X2 U6359 ( .A1(cv[35]), .A2(n7130), .ZN(n6786) );
  NAND2_X2 U6360 ( .A1(cv_next[35]), .A2(n7145), .ZN(n6785) );
  NAND2_X2 U6361 ( .A1(n6053), .A2(n6787), .ZN(cv_d[34]) );
  NAND2_X2 U6362 ( .A1(cv_q[34]), .A2(n7155), .ZN(n6787) );
  NAND2_X2 U6364 ( .A1(cv[34]), .A2(n7130), .ZN(n6789) );
  NAND2_X2 U6365 ( .A1(cv_next[34]), .A2(n7145), .ZN(n6788) );
  NAND2_X2 U6366 ( .A1(n6055), .A2(n6790), .ZN(cv_d[33]) );
  NAND2_X2 U6367 ( .A1(cv_q[33]), .A2(n7155), .ZN(n6790) );
  NAND2_X2 U6369 ( .A1(cv[33]), .A2(n7130), .ZN(n6792) );
  NAND2_X2 U6370 ( .A1(cv_next[33]), .A2(n7145), .ZN(n6791) );
  NAND2_X2 U6371 ( .A1(n6057), .A2(n6793), .ZN(cv_d[32]) );
  NAND2_X2 U6372 ( .A1(cv_q[32]), .A2(n7155), .ZN(n6793) );
  NAND2_X2 U6374 ( .A1(cv[32]), .A2(n7130), .ZN(n6795) );
  NAND2_X2 U6375 ( .A1(cv_next[32]), .A2(n7145), .ZN(n6794) );
  NAND2_X2 U6376 ( .A1(n6059), .A2(n6796), .ZN(cv_d[31]) );
  NAND2_X2 U6377 ( .A1(cv_q[31]), .A2(n7155), .ZN(n6796) );
  NAND2_X2 U6379 ( .A1(cv[31]), .A2(n7130), .ZN(n6798) );
  NAND2_X2 U6380 ( .A1(cv_next[31]), .A2(n7145), .ZN(n6797) );
  NAND2_X2 U6381 ( .A1(n6061), .A2(n6799), .ZN(cv_d[30]) );
  NAND2_X2 U6382 ( .A1(cv_q[30]), .A2(n7155), .ZN(n6799) );
  NAND2_X2 U6384 ( .A1(cv[30]), .A2(n7130), .ZN(n6801) );
  NAND2_X2 U6385 ( .A1(cv_next[30]), .A2(n7145), .ZN(n6800) );
  NAND2_X2 U6386 ( .A1(n6063), .A2(n6802), .ZN(cv_d[2]) );
  NAND2_X2 U6387 ( .A1(cv_q[2]), .A2(n7155), .ZN(n6802) );
  NAND2_X2 U6389 ( .A1(cv[2]), .A2(n7131), .ZN(n6804) );
  NAND2_X2 U6390 ( .A1(cv_next[2]), .A2(n7146), .ZN(n6803) );
  NAND2_X2 U6391 ( .A1(n6065), .A2(n6805), .ZN(cv_d[29]) );
  NAND2_X2 U6392 ( .A1(cv_q[29]), .A2(n7155), .ZN(n6805) );
  NAND2_X2 U6394 ( .A1(cv[29]), .A2(n7131), .ZN(n6807) );
  NAND2_X2 U6395 ( .A1(cv_next[29]), .A2(n7146), .ZN(n6806) );
  NAND2_X2 U6396 ( .A1(n6067), .A2(n6808), .ZN(cv_d[28]) );
  NAND2_X2 U6397 ( .A1(cv_q[28]), .A2(n7155), .ZN(n6808) );
  NAND2_X2 U6399 ( .A1(cv[28]), .A2(n7131), .ZN(n6810) );
  NAND2_X2 U6400 ( .A1(cv_next[28]), .A2(n7146), .ZN(n6809) );
  NAND2_X2 U6401 ( .A1(n6069), .A2(n6811), .ZN(cv_d[27]) );
  NAND2_X2 U6402 ( .A1(cv_q[27]), .A2(n7155), .ZN(n6811) );
  NAND2_X2 U6404 ( .A1(cv[27]), .A2(n7131), .ZN(n6813) );
  NAND2_X2 U6405 ( .A1(cv_next[27]), .A2(n7146), .ZN(n6812) );
  NAND2_X2 U6406 ( .A1(n6071), .A2(n6814), .ZN(cv_d[26]) );
  NAND2_X2 U6407 ( .A1(cv_q[26]), .A2(n7155), .ZN(n6814) );
  NAND2_X2 U6409 ( .A1(cv[26]), .A2(n7131), .ZN(n6816) );
  NAND2_X2 U6410 ( .A1(cv_next[26]), .A2(n7146), .ZN(n6815) );
  NAND2_X2 U6411 ( .A1(n6073), .A2(n6817), .ZN(cv_d[25]) );
  NAND2_X2 U6412 ( .A1(cv_q[25]), .A2(n7155), .ZN(n6817) );
  NAND2_X2 U6414 ( .A1(cv[25]), .A2(n7131), .ZN(n6819) );
  NAND2_X2 U6415 ( .A1(cv_next[25]), .A2(n7146), .ZN(n6818) );
  NAND2_X2 U6416 ( .A1(n6075), .A2(n6820), .ZN(cv_d[24]) );
  NAND2_X2 U6417 ( .A1(cv_q[24]), .A2(n7155), .ZN(n6820) );
  NAND2_X2 U6419 ( .A1(cv[24]), .A2(n7131), .ZN(n6822) );
  NAND2_X2 U6420 ( .A1(cv_next[24]), .A2(n7146), .ZN(n6821) );
  NAND2_X2 U6421 ( .A1(n6077), .A2(n6823), .ZN(cv_d[23]) );
  NAND2_X2 U6422 ( .A1(cv_q[23]), .A2(n7155), .ZN(n6823) );
  NAND2_X2 U6424 ( .A1(cv[23]), .A2(n7131), .ZN(n6825) );
  NAND2_X2 U6425 ( .A1(cv_next[23]), .A2(n7146), .ZN(n6824) );
  NAND2_X2 U6426 ( .A1(n6079), .A2(n6826), .ZN(cv_d[22]) );
  NAND2_X2 U6427 ( .A1(cv_q[22]), .A2(n7156), .ZN(n6826) );
  NAND2_X2 U6429 ( .A1(cv[22]), .A2(n7131), .ZN(n6828) );
  NAND2_X2 U6430 ( .A1(cv_next[22]), .A2(n7146), .ZN(n6827) );
  NAND2_X2 U6431 ( .A1(n6081), .A2(n6829), .ZN(cv_d[21]) );
  NAND2_X2 U6432 ( .A1(cv_q[21]), .A2(n7156), .ZN(n6829) );
  NAND2_X2 U6434 ( .A1(cv[21]), .A2(n7131), .ZN(n6831) );
  NAND2_X2 U6435 ( .A1(cv_next[21]), .A2(n7146), .ZN(n6830) );
  NAND2_X2 U6436 ( .A1(n6083), .A2(n6832), .ZN(cv_d[20]) );
  NAND2_X2 U6437 ( .A1(cv_q[20]), .A2(n7156), .ZN(n6832) );
  NAND2_X2 U6439 ( .A1(cv[20]), .A2(n7131), .ZN(n6834) );
  NAND2_X2 U6440 ( .A1(cv_next[20]), .A2(n7146), .ZN(n6833) );
  NAND2_X2 U6441 ( .A1(n6085), .A2(n6835), .ZN(cv_d[1]) );
  NAND2_X2 U6442 ( .A1(cv_q[1]), .A2(n7156), .ZN(n6835) );
  NAND2_X2 U6444 ( .A1(cv[1]), .A2(n7132), .ZN(n6837) );
  NAND2_X2 U6445 ( .A1(cv_next[1]), .A2(n7147), .ZN(n6836) );
  NAND2_X2 U6446 ( .A1(n6087), .A2(n6838), .ZN(cv_d[19]) );
  NAND2_X2 U6447 ( .A1(cv_q[19]), .A2(n7156), .ZN(n6838) );
  NAND2_X2 U6449 ( .A1(cv[19]), .A2(n7132), .ZN(n6840) );
  NAND2_X2 U6450 ( .A1(cv_next[19]), .A2(n7147), .ZN(n6839) );
  NAND2_X2 U6451 ( .A1(n6089), .A2(n6841), .ZN(cv_d[18]) );
  NAND2_X2 U6452 ( .A1(cv_q[18]), .A2(n7156), .ZN(n6841) );
  NAND2_X2 U6454 ( .A1(cv[18]), .A2(n7132), .ZN(n6843) );
  NAND2_X2 U6455 ( .A1(cv_next[18]), .A2(n7147), .ZN(n6842) );
  NAND2_X2 U6456 ( .A1(n6091), .A2(n6844), .ZN(cv_d[17]) );
  NAND2_X2 U6457 ( .A1(cv_q[17]), .A2(n7156), .ZN(n6844) );
  NAND2_X2 U6459 ( .A1(cv[17]), .A2(n7132), .ZN(n6846) );
  NAND2_X2 U6460 ( .A1(cv_next[17]), .A2(n7147), .ZN(n6845) );
  NAND2_X2 U6461 ( .A1(n6093), .A2(n6847), .ZN(cv_d[16]) );
  NAND2_X2 U6462 ( .A1(cv_q[16]), .A2(n7156), .ZN(n6847) );
  NAND2_X2 U6464 ( .A1(cv[16]), .A2(n7132), .ZN(n6849) );
  NAND2_X2 U6465 ( .A1(cv_next[16]), .A2(n7147), .ZN(n6848) );
  NAND2_X2 U6466 ( .A1(n6095), .A2(n6850), .ZN(cv_d[15]) );
  NAND2_X2 U6467 ( .A1(cv_q[15]), .A2(n7156), .ZN(n6850) );
  NAND2_X2 U6469 ( .A1(cv[15]), .A2(n7132), .ZN(n6852) );
  NAND2_X2 U6470 ( .A1(cv_next[15]), .A2(n7147), .ZN(n6851) );
  NAND2_X2 U6471 ( .A1(n7373), .A2(n6853), .ZN(cv_d[159]) );
  NAND2_X2 U6472 ( .A1(cv_q[159]), .A2(n7156), .ZN(n6853) );
  NAND2_X2 U6477 ( .A1(cv_q[158]), .A2(n7156), .ZN(n6856) );
  NAND2_X2 U6481 ( .A1(n7375), .A2(n6859), .ZN(cv_d[157]) );
  NAND2_X2 U6482 ( .A1(cv_q[157]), .A2(n7156), .ZN(n6859) );
  NAND2_X2 U6486 ( .A1(n7376), .A2(n6862), .ZN(cv_d[156]) );
  NAND2_X2 U6487 ( .A1(cv_q[156]), .A2(n7156), .ZN(n6862) );
  NAND2_X2 U6492 ( .A1(cv_q[155]), .A2(n7156), .ZN(n6865) );
  NAND2_X2 U6497 ( .A1(cv_q[154]), .A2(n7156), .ZN(n6868) );
  NAND2_X2 U6502 ( .A1(cv_q[153]), .A2(n7156), .ZN(n6871) );
  NAND2_X2 U6506 ( .A1(n7380), .A2(n6874), .ZN(cv_d[152]) );
  NAND2_X2 U6507 ( .A1(cv_q[152]), .A2(n7156), .ZN(n6874) );
  NAND2_X2 U6511 ( .A1(n7381), .A2(n6877), .ZN(cv_d[151]) );
  NAND2_X2 U6512 ( .A1(cv_q[151]), .A2(n7156), .ZN(n6877) );
  NAND2_X2 U6516 ( .A1(n7382), .A2(n6880), .ZN(cv_d[150]) );
  NAND2_X2 U6517 ( .A1(cv_q[150]), .A2(n7156), .ZN(n6880) );
  NAND2_X2 U6521 ( .A1(n6117), .A2(n6883), .ZN(cv_d[14]) );
  NAND2_X2 U6522 ( .A1(cv_q[14]), .A2(n7156), .ZN(n6883) );
  NAND2_X2 U6524 ( .A1(cv[14]), .A2(n7132), .ZN(n6885) );
  NAND2_X2 U6525 ( .A1(cv_next[14]), .A2(n7147), .ZN(n6884) );
  NAND2_X2 U6527 ( .A1(cv_q[149]), .A2(n7156), .ZN(n6886) );
  NAND2_X2 U6531 ( .A1(n7384), .A2(n6889), .ZN(cv_d[148]) );
  NAND2_X2 U6532 ( .A1(cv_q[148]), .A2(n7156), .ZN(n6889) );
  NAND2_X2 U6536 ( .A1(n7385), .A2(n6892), .ZN(cv_d[147]) );
  NAND2_X2 U6537 ( .A1(cv_q[147]), .A2(n7156), .ZN(n6892) );
  NAND2_X2 U6541 ( .A1(n7386), .A2(n6895), .ZN(cv_d[146]) );
  NAND2_X2 U6542 ( .A1(cv_q[146]), .A2(n7156), .ZN(n6895) );
  NAND2_X2 U6546 ( .A1(n7387), .A2(n6898), .ZN(cv_d[145]) );
  NAND2_X2 U6547 ( .A1(cv_q[145]), .A2(n7156), .ZN(n6898) );
  NAND2_X2 U6551 ( .A1(n7388), .A2(n6901), .ZN(cv_d[144]) );
  NAND2_X2 U6552 ( .A1(cv_q[144]), .A2(n7156), .ZN(n6901) );
  NAND2_X2 U6556 ( .A1(n7389), .A2(n6904), .ZN(cv_d[143]) );
  NAND2_X2 U6557 ( .A1(cv_q[143]), .A2(n7156), .ZN(n6904) );
  NAND2_X2 U6561 ( .A1(n7390), .A2(n6907), .ZN(cv_d[142]) );
  NAND2_X2 U6562 ( .A1(cv_q[142]), .A2(n7157), .ZN(n6907) );
  NAND2_X2 U6566 ( .A1(n7391), .A2(n6910), .ZN(cv_d[141]) );
  NAND2_X2 U6567 ( .A1(cv_q[141]), .A2(n7157), .ZN(n6910) );
  NAND2_X2 U6571 ( .A1(n7392), .A2(n6913), .ZN(cv_d[140]) );
  NAND2_X2 U6572 ( .A1(cv_q[140]), .A2(n7157), .ZN(n6913) );
  NAND2_X2 U6576 ( .A1(n6139), .A2(n6916), .ZN(cv_d[13]) );
  NAND2_X2 U6577 ( .A1(cv_q[13]), .A2(n7157), .ZN(n6916) );
  NAND2_X2 U6579 ( .A1(cv[13]), .A2(n7132), .ZN(n6918) );
  NAND2_X2 U6580 ( .A1(cv_next[13]), .A2(n7147), .ZN(n6917) );
  NAND2_X2 U6581 ( .A1(n7393), .A2(n6919), .ZN(cv_d[139]) );
  NAND2_X2 U6582 ( .A1(cv_q[139]), .A2(n7157), .ZN(n6919) );
  NAND2_X2 U6586 ( .A1(n7394), .A2(n6922), .ZN(cv_d[138]) );
  NAND2_X2 U6587 ( .A1(cv_q[138]), .A2(n7157), .ZN(n6922) );
  NAND2_X2 U6591 ( .A1(n6145), .A2(n6925), .ZN(cv_d[137]) );
  NAND2_X2 U6592 ( .A1(cv_q[137]), .A2(n7157), .ZN(n6925) );
  NAND2_X2 U6594 ( .A1(cv[137]), .A2(n7132), .ZN(n6927) );
  NAND2_X2 U6595 ( .A1(cv_next[137]), .A2(n7147), .ZN(n6926) );
  NAND2_X2 U6596 ( .A1(n6147), .A2(n6928), .ZN(cv_d[136]) );
  NAND2_X2 U6597 ( .A1(cv_q[136]), .A2(n7157), .ZN(n6928) );
  NAND2_X2 U6599 ( .A1(cv[136]), .A2(n7132), .ZN(n6930) );
  NAND2_X2 U6600 ( .A1(cv_next[136]), .A2(n7147), .ZN(n6929) );
  NAND2_X2 U6601 ( .A1(n6149), .A2(n6931), .ZN(cv_d[135]) );
  NAND2_X2 U6602 ( .A1(cv_q[135]), .A2(n7157), .ZN(n6931) );
  NAND2_X2 U6604 ( .A1(cv[135]), .A2(n7132), .ZN(n6933) );
  NAND2_X2 U6605 ( .A1(cv_next[135]), .A2(n7147), .ZN(n6932) );
  NAND2_X2 U6606 ( .A1(n6151), .A2(n6934), .ZN(cv_d[134]) );
  NAND2_X2 U6607 ( .A1(cv_q[134]), .A2(n7157), .ZN(n6934) );
  NAND2_X2 U6609 ( .A1(cv[134]), .A2(n7133), .ZN(n6936) );
  NAND2_X2 U6610 ( .A1(cv_next[134]), .A2(n7148), .ZN(n6935) );
  NAND2_X2 U6611 ( .A1(n6153), .A2(n6937), .ZN(cv_d[133]) );
  NAND2_X2 U6612 ( .A1(cv_q[133]), .A2(n7157), .ZN(n6937) );
  NAND2_X2 U6614 ( .A1(cv[133]), .A2(n7133), .ZN(n6939) );
  NAND2_X2 U6615 ( .A1(cv_next[133]), .A2(n7148), .ZN(n6938) );
  NAND2_X2 U6616 ( .A1(n6155), .A2(n6940), .ZN(cv_d[132]) );
  NAND2_X2 U6617 ( .A1(cv_q[132]), .A2(n7157), .ZN(n6940) );
  NAND2_X2 U6619 ( .A1(cv[132]), .A2(n7133), .ZN(n6942) );
  NAND2_X2 U6620 ( .A1(cv_next[132]), .A2(n7148), .ZN(n6941) );
  NAND2_X2 U6621 ( .A1(n6157), .A2(n6943), .ZN(cv_d[131]) );
  NAND2_X2 U6622 ( .A1(cv_q[131]), .A2(n7157), .ZN(n6943) );
  NAND2_X2 U6624 ( .A1(cv[131]), .A2(n7133), .ZN(n6945) );
  NAND2_X2 U6625 ( .A1(cv_next[131]), .A2(n7148), .ZN(n6944) );
  NAND2_X2 U6626 ( .A1(n6159), .A2(n6946), .ZN(cv_d[130]) );
  NAND2_X2 U6627 ( .A1(cv_q[130]), .A2(n7157), .ZN(n6946) );
  NAND2_X2 U6629 ( .A1(cv[130]), .A2(n7133), .ZN(n6948) );
  NAND2_X2 U6630 ( .A1(cv_next[130]), .A2(n7148), .ZN(n6947) );
  NAND2_X2 U6631 ( .A1(n6161), .A2(n6949), .ZN(cv_d[12]) );
  NAND2_X2 U6632 ( .A1(cv_q[12]), .A2(n7157), .ZN(n6949) );
  NAND2_X2 U6634 ( .A1(cv[12]), .A2(n7133), .ZN(n6951) );
  NAND2_X2 U6635 ( .A1(cv_next[12]), .A2(n7148), .ZN(n6950) );
  NAND2_X2 U6636 ( .A1(n6163), .A2(n6952), .ZN(cv_d[129]) );
  NAND2_X2 U6637 ( .A1(cv_q[129]), .A2(n7157), .ZN(n6952) );
  NAND2_X2 U6639 ( .A1(cv[129]), .A2(n7133), .ZN(n6954) );
  NAND2_X2 U6640 ( .A1(cv_next[129]), .A2(n7148), .ZN(n6953) );
  NAND2_X2 U6641 ( .A1(n6165), .A2(n6955), .ZN(cv_d[128]) );
  NAND2_X2 U6642 ( .A1(cv_q[128]), .A2(n7157), .ZN(n6955) );
  NAND2_X2 U6644 ( .A1(cv[128]), .A2(n7133), .ZN(n6957) );
  NAND2_X2 U6645 ( .A1(cv_next[128]), .A2(n7148), .ZN(n6956) );
  NAND2_X2 U6646 ( .A1(n6167), .A2(n6958), .ZN(cv_d[127]) );
  NAND2_X2 U6647 ( .A1(cv_q[127]), .A2(n7157), .ZN(n6958) );
  NAND2_X2 U6649 ( .A1(cv[127]), .A2(n7133), .ZN(n6960) );
  NAND2_X2 U6650 ( .A1(cv_next[127]), .A2(n7148), .ZN(n6959) );
  NAND2_X2 U6651 ( .A1(n6169), .A2(n6961), .ZN(cv_d[126]) );
  NAND2_X2 U6652 ( .A1(cv_q[126]), .A2(n7157), .ZN(n6961) );
  NAND2_X2 U6654 ( .A1(cv[126]), .A2(n7133), .ZN(n6963) );
  NAND2_X2 U6655 ( .A1(cv_next[126]), .A2(n7148), .ZN(n6962) );
  NAND2_X2 U6656 ( .A1(n6171), .A2(n6964), .ZN(cv_d[125]) );
  NAND2_X2 U6657 ( .A1(cv_q[125]), .A2(n7157), .ZN(n6964) );
  NAND2_X2 U6659 ( .A1(cv[125]), .A2(n7133), .ZN(n6966) );
  NAND2_X2 U6660 ( .A1(cv_next[125]), .A2(n7148), .ZN(n6965) );
  NAND2_X2 U6661 ( .A1(n6173), .A2(n6967), .ZN(cv_d[124]) );
  NAND2_X2 U6662 ( .A1(cv_q[124]), .A2(n7157), .ZN(n6967) );
  NAND2_X2 U6664 ( .A1(cv[124]), .A2(n7134), .ZN(n6969) );
  NAND2_X2 U6665 ( .A1(cv_next[124]), .A2(n7149), .ZN(n6968) );
  NAND2_X2 U6666 ( .A1(n6175), .A2(n6970), .ZN(cv_d[123]) );
  NAND2_X2 U6667 ( .A1(cv_q[123]), .A2(n7157), .ZN(n6970) );
  NAND2_X2 U6669 ( .A1(cv[123]), .A2(n7134), .ZN(n6972) );
  NAND2_X2 U6670 ( .A1(cv_next[123]), .A2(n7149), .ZN(n6971) );
  NAND2_X2 U6671 ( .A1(n6177), .A2(n6973), .ZN(cv_d[122]) );
  NAND2_X2 U6672 ( .A1(cv_q[122]), .A2(n7157), .ZN(n6973) );
  NAND2_X2 U6674 ( .A1(cv[122]), .A2(n7134), .ZN(n6975) );
  NAND2_X2 U6675 ( .A1(cv_next[122]), .A2(n7149), .ZN(n6974) );
  NAND2_X2 U6676 ( .A1(n6179), .A2(n6976), .ZN(cv_d[121]) );
  NAND2_X2 U6677 ( .A1(cv_q[121]), .A2(n7157), .ZN(n6976) );
  NAND2_X2 U6679 ( .A1(cv[121]), .A2(n7134), .ZN(n6978) );
  NAND2_X2 U6680 ( .A1(cv_next[121]), .A2(n7149), .ZN(n6977) );
  NAND2_X2 U6681 ( .A1(n6181), .A2(n6979), .ZN(cv_d[120]) );
  NAND2_X2 U6682 ( .A1(cv_q[120]), .A2(n7157), .ZN(n6979) );
  NAND2_X2 U6684 ( .A1(cv[120]), .A2(n7134), .ZN(n6981) );
  NAND2_X2 U6685 ( .A1(cv_next[120]), .A2(n7149), .ZN(n6980) );
  NAND2_X2 U6686 ( .A1(n6183), .A2(n6982), .ZN(cv_d[11]) );
  NAND2_X2 U6687 ( .A1(cv_q[11]), .A2(n7157), .ZN(n6982) );
  NAND2_X2 U6689 ( .A1(cv[11]), .A2(n7134), .ZN(n6984) );
  NAND2_X2 U6690 ( .A1(cv_next[11]), .A2(n7149), .ZN(n6983) );
  NAND2_X2 U6691 ( .A1(n6185), .A2(n6985), .ZN(cv_d[119]) );
  NAND2_X2 U6692 ( .A1(cv_q[119]), .A2(n7157), .ZN(n6985) );
  NAND2_X2 U6694 ( .A1(cv[119]), .A2(n7134), .ZN(n6987) );
  NAND2_X2 U6695 ( .A1(cv_next[119]), .A2(n7149), .ZN(n6986) );
  NAND2_X2 U6696 ( .A1(n6187), .A2(n6988), .ZN(cv_d[118]) );
  NAND2_X2 U6697 ( .A1(cv_q[118]), .A2(n7158), .ZN(n6988) );
  NAND2_X2 U6699 ( .A1(cv[118]), .A2(n7134), .ZN(n6990) );
  NAND2_X2 U6700 ( .A1(cv_next[118]), .A2(n7149), .ZN(n6989) );
  NAND2_X2 U6701 ( .A1(n6189), .A2(n6991), .ZN(cv_d[117]) );
  NAND2_X2 U6702 ( .A1(cv_q[117]), .A2(n7158), .ZN(n6991) );
  NAND2_X2 U6704 ( .A1(cv[117]), .A2(n7134), .ZN(n6993) );
  NAND2_X2 U6705 ( .A1(cv_next[117]), .A2(n7149), .ZN(n6992) );
  NAND2_X2 U6706 ( .A1(n6191), .A2(n6994), .ZN(cv_d[116]) );
  NAND2_X2 U6707 ( .A1(cv_q[116]), .A2(n7158), .ZN(n6994) );
  NAND2_X2 U6709 ( .A1(cv[116]), .A2(n7134), .ZN(n6996) );
  NAND2_X2 U6710 ( .A1(cv_next[116]), .A2(n7149), .ZN(n6995) );
  NAND2_X2 U6711 ( .A1(n6193), .A2(n6997), .ZN(cv_d[115]) );
  NAND2_X2 U6712 ( .A1(cv_q[115]), .A2(n7158), .ZN(n6997) );
  NAND2_X2 U6714 ( .A1(cv[115]), .A2(n7134), .ZN(n6999) );
  NAND2_X2 U6715 ( .A1(cv_next[115]), .A2(n7149), .ZN(n6998) );
  NAND2_X2 U6716 ( .A1(n6195), .A2(n7000), .ZN(cv_d[114]) );
  NAND2_X2 U6717 ( .A1(cv_q[114]), .A2(n7158), .ZN(n7000) );
  NAND2_X2 U6719 ( .A1(cv[114]), .A2(n7135), .ZN(n7002) );
  NAND2_X2 U6720 ( .A1(cv_next[114]), .A2(n7150), .ZN(n7001) );
  NAND2_X2 U6721 ( .A1(n6197), .A2(n7003), .ZN(cv_d[113]) );
  NAND2_X2 U6722 ( .A1(cv_q[113]), .A2(n7158), .ZN(n7003) );
  NAND2_X2 U6724 ( .A1(cv[113]), .A2(n7135), .ZN(n7005) );
  NAND2_X2 U6725 ( .A1(cv_next[113]), .A2(n7150), .ZN(n7004) );
  NAND2_X2 U6726 ( .A1(n6199), .A2(n7006), .ZN(cv_d[112]) );
  NAND2_X2 U6727 ( .A1(cv_q[112]), .A2(n7158), .ZN(n7006) );
  NAND2_X2 U6729 ( .A1(cv[112]), .A2(n7135), .ZN(n7008) );
  NAND2_X2 U6730 ( .A1(cv_next[112]), .A2(n7150), .ZN(n7007) );
  NAND2_X2 U6731 ( .A1(n6201), .A2(n7009), .ZN(cv_d[111]) );
  NAND2_X2 U6732 ( .A1(cv_q[111]), .A2(n7158), .ZN(n7009) );
  NAND2_X2 U6734 ( .A1(cv[111]), .A2(n7135), .ZN(n7011) );
  NAND2_X2 U6735 ( .A1(cv_next[111]), .A2(n7150), .ZN(n7010) );
  NAND2_X2 U6736 ( .A1(n6203), .A2(n7012), .ZN(cv_d[110]) );
  NAND2_X2 U6737 ( .A1(cv_q[110]), .A2(n7158), .ZN(n7012) );
  NAND2_X2 U6739 ( .A1(cv[110]), .A2(n7135), .ZN(n7014) );
  NAND2_X2 U6740 ( .A1(cv_next[110]), .A2(n7150), .ZN(n7013) );
  NAND2_X2 U6741 ( .A1(n6205), .A2(n7015), .ZN(cv_d[10]) );
  NAND2_X2 U6742 ( .A1(cv_q[10]), .A2(n7158), .ZN(n7015) );
  NAND2_X2 U6744 ( .A1(cv[10]), .A2(n7135), .ZN(n7017) );
  NAND2_X2 U6745 ( .A1(cv_next[10]), .A2(n7150), .ZN(n7016) );
  NAND2_X2 U6746 ( .A1(n6207), .A2(n7018), .ZN(cv_d[109]) );
  NAND2_X2 U6747 ( .A1(cv_q[109]), .A2(n7158), .ZN(n7018) );
  NAND2_X2 U6749 ( .A1(cv[109]), .A2(n7135), .ZN(n7020) );
  NAND2_X2 U6750 ( .A1(cv_next[109]), .A2(n7150), .ZN(n7019) );
  NAND2_X2 U6751 ( .A1(n6209), .A2(n7021), .ZN(cv_d[108]) );
  NAND2_X2 U6752 ( .A1(cv_q[108]), .A2(n7158), .ZN(n7021) );
  NAND2_X2 U6754 ( .A1(cv[108]), .A2(n7135), .ZN(n7023) );
  NAND2_X2 U6755 ( .A1(cv_next[108]), .A2(n7150), .ZN(n7022) );
  NAND2_X2 U6756 ( .A1(n6211), .A2(n7024), .ZN(cv_d[107]) );
  NAND2_X2 U6757 ( .A1(cv_q[107]), .A2(n7158), .ZN(n7024) );
  NAND2_X2 U6759 ( .A1(cv[107]), .A2(n7135), .ZN(n7026) );
  NAND2_X2 U6760 ( .A1(cv_next[107]), .A2(n7150), .ZN(n7025) );
  NAND2_X2 U6761 ( .A1(n6213), .A2(n7027), .ZN(cv_d[106]) );
  NAND2_X2 U6762 ( .A1(cv_q[106]), .A2(n7158), .ZN(n7027) );
  NAND2_X2 U6764 ( .A1(cv[106]), .A2(n7135), .ZN(n7029) );
  NAND2_X2 U6765 ( .A1(cv_next[106]), .A2(n7150), .ZN(n7028) );
  NAND2_X2 U6766 ( .A1(n6215), .A2(n7030), .ZN(cv_d[105]) );
  NAND2_X2 U6767 ( .A1(cv_q[105]), .A2(n7158), .ZN(n7030) );
  NAND2_X2 U6769 ( .A1(cv[105]), .A2(n7135), .ZN(n7032) );
  NAND2_X2 U6770 ( .A1(cv_next[105]), .A2(n7150), .ZN(n7031) );
  NAND2_X2 U6771 ( .A1(n6217), .A2(n7033), .ZN(cv_d[104]) );
  NAND2_X2 U6772 ( .A1(cv_q[104]), .A2(n7158), .ZN(n7033) );
  NAND2_X2 U6774 ( .A1(cv[104]), .A2(n7136), .ZN(n7035) );
  NAND2_X2 U6775 ( .A1(cv_next[104]), .A2(n7151), .ZN(n7034) );
  NAND2_X2 U6776 ( .A1(n6219), .A2(n7036), .ZN(cv_d[103]) );
  NAND2_X2 U6777 ( .A1(cv_q[103]), .A2(n7158), .ZN(n7036) );
  NAND2_X2 U6779 ( .A1(cv[103]), .A2(n7136), .ZN(n7038) );
  NAND2_X2 U6780 ( .A1(cv_next[103]), .A2(n7151), .ZN(n7037) );
  NAND2_X2 U6781 ( .A1(n6221), .A2(n7039), .ZN(cv_d[102]) );
  NAND2_X2 U6782 ( .A1(cv_q[102]), .A2(n7158), .ZN(n7039) );
  NAND2_X2 U6784 ( .A1(cv[102]), .A2(n7136), .ZN(n7041) );
  NAND2_X2 U6785 ( .A1(cv_next[102]), .A2(n7151), .ZN(n7040) );
  NAND2_X2 U6786 ( .A1(n6223), .A2(n7042), .ZN(cv_d[101]) );
  NAND2_X2 U6787 ( .A1(cv_q[101]), .A2(n7158), .ZN(n7042) );
  NAND2_X2 U6789 ( .A1(cv[101]), .A2(n7136), .ZN(n7044) );
  NAND2_X2 U6790 ( .A1(cv_next[101]), .A2(n7151), .ZN(n7043) );
  NAND2_X2 U6791 ( .A1(n6225), .A2(n7045), .ZN(cv_d[100]) );
  NAND2_X2 U6792 ( .A1(cv_q[100]), .A2(n7158), .ZN(n7045) );
  NAND2_X2 U6794 ( .A1(cv[100]), .A2(n7136), .ZN(n7047) );
  NAND2_X2 U6795 ( .A1(cv_next[100]), .A2(n7151), .ZN(n7046) );
  NAND2_X2 U6796 ( .A1(n6227), .A2(n7048), .ZN(cv_d[0]) );
  NAND2_X2 U6797 ( .A1(cv_q[0]), .A2(n7158), .ZN(n7048) );
  NAND2_X2 U6799 ( .A1(cv[0]), .A2(n7136), .ZN(n7050) );
  NAND2_X2 U6801 ( .A1(cv_next[0]), .A2(n7151), .ZN(n7049) );
  NAND2_X2 U6803 ( .A1(state[0]), .A2(n7395), .ZN(busy) );
  NAND2_X1 U6818 ( .A1(n7377), .A2(n6865), .ZN(cv_d[155]) );
  NAND2_X4 U6819 ( .A1(n7372), .A2(n7373), .ZN(rnd_d[159]) );
  INV_X8 U6820 ( .A(n7118), .ZN(n7119) );
  NAND2_X4 U6821 ( .A1(sha1_round_wire[151]), .A2(n7159), .ZN(n7340) );
  NAND2_X4 U6822 ( .A1(sha1_round_wire[159]), .A2(n7159), .ZN(n7372) );
  NAND2_X2 U6823 ( .A1(n7381), .A2(n7340), .ZN(rnd_d[151]) );
  NAND2_X2 U6824 ( .A1(sha1_round_wire[157]), .A2(n7159), .ZN(n7364) );
  INV_X8 U6825 ( .A(rnd_cnt_q[2]), .ZN(n7118) );
  NAND2_X2 U6826 ( .A1(n7356), .A2(n7377), .ZN(rnd_d[155]) );
  INV_X1 U6827 ( .A(n7331), .ZN(n7383) );
  INV_X1 U6828 ( .A(n7351), .ZN(n7378) );
  INV_X1 U6829 ( .A(n7367), .ZN(n7374) );
  INV_X1 U6830 ( .A(n7347), .ZN(n7379) );
  AND2_X1 U6831 ( .A1(n7049), .A2(n7050), .ZN(n6227) );
  AND2_X1 U6832 ( .A1(n6836), .A2(n6837), .ZN(n6085) );
  AND2_X1 U6833 ( .A1(n6803), .A2(n6804), .ZN(n6063) );
  AND2_X1 U6834 ( .A1(n6770), .A2(n6771), .ZN(n6041) );
  AND2_X1 U6835 ( .A1(n6737), .A2(n6738), .ZN(n6019) );
  AND2_X1 U6836 ( .A1(n6704), .A2(n6705), .ZN(n5997) );
  AND2_X1 U6837 ( .A1(n6671), .A2(n6672), .ZN(n5975) );
  AND2_X1 U6838 ( .A1(n6638), .A2(n6639), .ZN(n5953) );
  AND2_X1 U6839 ( .A1(n6605), .A2(n6606), .ZN(n5931) );
  AND2_X1 U6840 ( .A1(n6570), .A2(n6571), .ZN(n5909) );
  AND2_X1 U6841 ( .A1(n7016), .A2(n7017), .ZN(n6205) );
  AND2_X1 U6842 ( .A1(n6983), .A2(n6984), .ZN(n6183) );
  AND2_X1 U6843 ( .A1(n6950), .A2(n6951), .ZN(n6161) );
  AND2_X1 U6844 ( .A1(n6917), .A2(n6918), .ZN(n6139) );
  AND2_X1 U6845 ( .A1(n6884), .A2(n6885), .ZN(n6117) );
  AND2_X1 U6846 ( .A1(n6851), .A2(n6852), .ZN(n6095) );
  AND2_X1 U6847 ( .A1(n6848), .A2(n6849), .ZN(n6093) );
  AND2_X1 U6848 ( .A1(n6845), .A2(n6846), .ZN(n6091) );
  AND2_X1 U6849 ( .A1(n6842), .A2(n6843), .ZN(n6089) );
  AND2_X1 U6850 ( .A1(n6839), .A2(n6840), .ZN(n6087) );
  AND2_X1 U6851 ( .A1(n6833), .A2(n6834), .ZN(n6083) );
  AND2_X1 U6852 ( .A1(n6830), .A2(n6831), .ZN(n6081) );
  AND2_X1 U6853 ( .A1(n6827), .A2(n6828), .ZN(n6079) );
  AND2_X1 U6854 ( .A1(n6824), .A2(n6825), .ZN(n6077) );
  AND2_X1 U6855 ( .A1(n6821), .A2(n6822), .ZN(n6075) );
  AND2_X1 U6856 ( .A1(n6818), .A2(n6819), .ZN(n6073) );
  AND2_X1 U6857 ( .A1(n6815), .A2(n6816), .ZN(n6071) );
  AND2_X1 U6858 ( .A1(n6812), .A2(n6813), .ZN(n6069) );
  AND2_X1 U6859 ( .A1(n6809), .A2(n6810), .ZN(n6067) );
  AND2_X1 U6860 ( .A1(n6806), .A2(n6807), .ZN(n6065) );
  AND2_X1 U6861 ( .A1(n6800), .A2(n6801), .ZN(n6061) );
  AND2_X1 U6862 ( .A1(n6797), .A2(n6798), .ZN(n6059) );
  AND2_X1 U6863 ( .A1(n6794), .A2(n6795), .ZN(n6057) );
  AND2_X1 U6864 ( .A1(n6791), .A2(n6792), .ZN(n6055) );
  AND2_X1 U6865 ( .A1(n6788), .A2(n6789), .ZN(n6053) );
  AND2_X1 U6866 ( .A1(n6785), .A2(n6786), .ZN(n6051) );
  AND2_X1 U6867 ( .A1(n6782), .A2(n6783), .ZN(n6049) );
  AND2_X1 U6868 ( .A1(n6779), .A2(n6780), .ZN(n6047) );
  AND2_X1 U6869 ( .A1(n6776), .A2(n6777), .ZN(n6045) );
  AND2_X1 U6870 ( .A1(n6773), .A2(n6774), .ZN(n6043) );
  AND2_X1 U6871 ( .A1(n6767), .A2(n6768), .ZN(n6039) );
  AND2_X1 U6872 ( .A1(n6764), .A2(n6765), .ZN(n6037) );
  AND2_X1 U6873 ( .A1(n6761), .A2(n6762), .ZN(n6035) );
  AND2_X1 U6874 ( .A1(n6758), .A2(n6759), .ZN(n6033) );
  AND2_X1 U6875 ( .A1(n6755), .A2(n6756), .ZN(n6031) );
  AND2_X1 U6876 ( .A1(n6752), .A2(n6753), .ZN(n6029) );
  AND2_X1 U6877 ( .A1(n6749), .A2(n6750), .ZN(n6027) );
  AND2_X1 U6878 ( .A1(n6746), .A2(n6747), .ZN(n6025) );
  AND2_X1 U6879 ( .A1(n6743), .A2(n6744), .ZN(n6023) );
  AND2_X1 U6880 ( .A1(n6740), .A2(n6741), .ZN(n6021) );
  AND2_X1 U6881 ( .A1(n6734), .A2(n6735), .ZN(n6017) );
  AND2_X1 U6882 ( .A1(n6731), .A2(n6732), .ZN(n6015) );
  AND2_X1 U6883 ( .A1(n6728), .A2(n6729), .ZN(n6013) );
  AND2_X1 U6884 ( .A1(n6725), .A2(n6726), .ZN(n6011) );
  AND2_X1 U6885 ( .A1(n6722), .A2(n6723), .ZN(n6009) );
  AND2_X1 U6886 ( .A1(n6719), .A2(n6720), .ZN(n6007) );
  AND2_X1 U6887 ( .A1(n6716), .A2(n6717), .ZN(n6005) );
  AND2_X1 U6888 ( .A1(n6713), .A2(n6714), .ZN(n6003) );
  AND2_X1 U6889 ( .A1(n6710), .A2(n6711), .ZN(n6001) );
  AND2_X1 U6890 ( .A1(n6707), .A2(n6708), .ZN(n5999) );
  AND2_X1 U6891 ( .A1(n6701), .A2(n6702), .ZN(n5995) );
  AND2_X1 U6892 ( .A1(n6698), .A2(n6699), .ZN(n5993) );
  AND2_X1 U6893 ( .A1(n6695), .A2(n6696), .ZN(n5991) );
  AND2_X1 U6894 ( .A1(n6692), .A2(n6693), .ZN(n5989) );
  AND2_X1 U6895 ( .A1(n6689), .A2(n6690), .ZN(n5987) );
  AND2_X1 U6896 ( .A1(n6686), .A2(n6687), .ZN(n5985) );
  AND2_X1 U6897 ( .A1(n6683), .A2(n6684), .ZN(n5983) );
  AND2_X1 U6898 ( .A1(n6680), .A2(n6681), .ZN(n5981) );
  AND2_X1 U6899 ( .A1(n6677), .A2(n6678), .ZN(n5979) );
  AND2_X1 U6900 ( .A1(n6674), .A2(n6675), .ZN(n5977) );
  AND2_X1 U6901 ( .A1(n6668), .A2(n6669), .ZN(n5973) );
  AND2_X1 U6902 ( .A1(n6665), .A2(n6666), .ZN(n5971) );
  AND2_X1 U6903 ( .A1(n6662), .A2(n6663), .ZN(n5969) );
  AND2_X1 U6904 ( .A1(n6659), .A2(n6660), .ZN(n5967) );
  AND2_X1 U6905 ( .A1(n6656), .A2(n6657), .ZN(n5965) );
  AND2_X1 U6906 ( .A1(n6653), .A2(n6654), .ZN(n5963) );
  AND2_X1 U6907 ( .A1(n6650), .A2(n6651), .ZN(n5961) );
  AND2_X1 U6908 ( .A1(n6647), .A2(n6648), .ZN(n5959) );
  AND2_X1 U6909 ( .A1(n6644), .A2(n6645), .ZN(n5957) );
  AND2_X1 U6910 ( .A1(n6641), .A2(n6642), .ZN(n5955) );
  AND2_X1 U6911 ( .A1(n6635), .A2(n6636), .ZN(n5951) );
  AND2_X1 U6912 ( .A1(n6632), .A2(n6633), .ZN(n5949) );
  AND2_X1 U6913 ( .A1(n6629), .A2(n6630), .ZN(n5947) );
  AND2_X1 U6914 ( .A1(n6626), .A2(n6627), .ZN(n5945) );
  AND2_X1 U6915 ( .A1(n6623), .A2(n6624), .ZN(n5943) );
  AND2_X1 U6916 ( .A1(n6620), .A2(n6621), .ZN(n5941) );
  AND2_X1 U6917 ( .A1(n6617), .A2(n6618), .ZN(n5939) );
  AND2_X1 U6918 ( .A1(n6614), .A2(n6615), .ZN(n5937) );
  AND2_X1 U6919 ( .A1(n6611), .A2(n6612), .ZN(n5935) );
  AND2_X1 U6920 ( .A1(n6608), .A2(n6609), .ZN(n5933) );
  AND2_X1 U6921 ( .A1(n6602), .A2(n6603), .ZN(n5929) );
  AND2_X1 U6922 ( .A1(n6599), .A2(n6600), .ZN(n5927) );
  AND2_X1 U6923 ( .A1(n6596), .A2(n6597), .ZN(n5925) );
  AND2_X1 U6924 ( .A1(n6593), .A2(n6594), .ZN(n5923) );
  AND2_X1 U6925 ( .A1(n6590), .A2(n6591), .ZN(n5921) );
  AND2_X1 U6926 ( .A1(n6587), .A2(n6588), .ZN(n5919) );
  AND2_X1 U6927 ( .A1(n6584), .A2(n6585), .ZN(n5917) );
  AND2_X1 U6928 ( .A1(n6581), .A2(n6582), .ZN(n5915) );
  AND2_X1 U6929 ( .A1(n6578), .A2(n6579), .ZN(n5913) );
  AND2_X1 U6930 ( .A1(n6575), .A2(n6576), .ZN(n5911) );
  AND2_X1 U6931 ( .A1(n7046), .A2(n7047), .ZN(n6225) );
  AND2_X1 U6932 ( .A1(n7043), .A2(n7044), .ZN(n6223) );
  AND2_X1 U6933 ( .A1(n7040), .A2(n7041), .ZN(n6221) );
  AND2_X1 U6934 ( .A1(n7037), .A2(n7038), .ZN(n6219) );
  AND2_X1 U6935 ( .A1(n7034), .A2(n7035), .ZN(n6217) );
  AND2_X1 U6936 ( .A1(n7031), .A2(n7032), .ZN(n6215) );
  AND2_X1 U6937 ( .A1(n7028), .A2(n7029), .ZN(n6213) );
  AND2_X1 U6938 ( .A1(n7025), .A2(n7026), .ZN(n6211) );
  AND2_X1 U6939 ( .A1(n7022), .A2(n7023), .ZN(n6209) );
  AND2_X1 U6940 ( .A1(n7019), .A2(n7020), .ZN(n6207) );
  AND2_X1 U6941 ( .A1(n7013), .A2(n7014), .ZN(n6203) );
  AND2_X1 U6942 ( .A1(n7010), .A2(n7011), .ZN(n6201) );
  AND2_X1 U6943 ( .A1(n7007), .A2(n7008), .ZN(n6199) );
  AND2_X1 U6944 ( .A1(n7004), .A2(n7005), .ZN(n6197) );
  AND2_X1 U6945 ( .A1(n7001), .A2(n7002), .ZN(n6195) );
  AND2_X1 U6946 ( .A1(n6998), .A2(n6999), .ZN(n6193) );
  AND2_X1 U6947 ( .A1(n6995), .A2(n6996), .ZN(n6191) );
  AND2_X1 U6948 ( .A1(n6992), .A2(n6993), .ZN(n6189) );
  AND2_X1 U6949 ( .A1(n6989), .A2(n6990), .ZN(n6187) );
  AND2_X1 U6950 ( .A1(n6986), .A2(n6987), .ZN(n6185) );
  AND2_X1 U6951 ( .A1(n6980), .A2(n6981), .ZN(n6181) );
  AND2_X1 U6952 ( .A1(n6977), .A2(n6978), .ZN(n6179) );
  AND2_X1 U6953 ( .A1(n6974), .A2(n6975), .ZN(n6177) );
  AND2_X1 U6954 ( .A1(n6971), .A2(n6972), .ZN(n6175) );
  AND2_X1 U6955 ( .A1(n6968), .A2(n6969), .ZN(n6173) );
  AND2_X1 U6956 ( .A1(n6965), .A2(n6966), .ZN(n6171) );
  AND2_X1 U6957 ( .A1(n6962), .A2(n6963), .ZN(n6169) );
  AND2_X1 U6958 ( .A1(n6959), .A2(n6960), .ZN(n6167) );
  AND2_X1 U6959 ( .A1(n6956), .A2(n6957), .ZN(n6165) );
  AND2_X1 U6960 ( .A1(n6953), .A2(n6954), .ZN(n6163) );
  AND2_X1 U6961 ( .A1(n6947), .A2(n6948), .ZN(n6159) );
  AND2_X1 U6962 ( .A1(n6944), .A2(n6945), .ZN(n6157) );
  AND2_X1 U6963 ( .A1(n6941), .A2(n6942), .ZN(n6155) );
  AND2_X1 U6964 ( .A1(n6938), .A2(n6939), .ZN(n6153) );
  AND2_X1 U6965 ( .A1(n6935), .A2(n6936), .ZN(n6151) );
  AND2_X1 U6966 ( .A1(n6932), .A2(n6933), .ZN(n6149) );
  AND2_X1 U6967 ( .A1(n6929), .A2(n6930), .ZN(n6147) );
  AND2_X1 U6968 ( .A1(n6926), .A2(n6927), .ZN(n6145) );
  INV_X8 U6969 ( .A(n7287), .ZN(n7394) );
  NAND2_X1 U6970 ( .A1(cv[138]), .A2(n7122), .ZN(n7286) );
  NAND2_X1 U6971 ( .A1(n7286), .A2(n7285), .ZN(n7287) );
  INV_X8 U6972 ( .A(n7291), .ZN(n7393) );
  NAND2_X1 U6973 ( .A1(cv[139]), .A2(n7122), .ZN(n7290) );
  NAND2_X1 U6974 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
  INV_X8 U6975 ( .A(n7295), .ZN(n7392) );
  NAND2_X1 U6976 ( .A1(cv[140]), .A2(n7122), .ZN(n7294) );
  NAND2_X1 U6977 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  INV_X8 U6978 ( .A(n7299), .ZN(n7391) );
  NAND2_X1 U6979 ( .A1(cv[141]), .A2(n7122), .ZN(n7298) );
  NAND2_X1 U6980 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  INV_X8 U6981 ( .A(n7303), .ZN(n7390) );
  NAND2_X1 U6982 ( .A1(cv[142]), .A2(n7122), .ZN(n7302) );
  NAND2_X1 U6983 ( .A1(n7302), .A2(n7301), .ZN(n7303) );
  INV_X8 U6984 ( .A(n7307), .ZN(n7389) );
  NAND2_X1 U6985 ( .A1(cv[143]), .A2(n7122), .ZN(n7306) );
  NAND2_X1 U6986 ( .A1(n7306), .A2(n7305), .ZN(n7307) );
  INV_X8 U6987 ( .A(n7311), .ZN(n7388) );
  NAND2_X1 U6988 ( .A1(cv[144]), .A2(n7122), .ZN(n7310) );
  NAND2_X1 U6989 ( .A1(n7310), .A2(n7309), .ZN(n7311) );
  INV_X8 U6990 ( .A(n7315), .ZN(n7387) );
  NAND2_X1 U6991 ( .A1(cv[145]), .A2(n7122), .ZN(n7314) );
  NAND2_X1 U6992 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  INV_X8 U6993 ( .A(n7319), .ZN(n7386) );
  NAND2_X1 U6994 ( .A1(cv[146]), .A2(n7122), .ZN(n7318) );
  NAND2_X1 U6995 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
  INV_X8 U6996 ( .A(n7323), .ZN(n7385) );
  NAND2_X1 U6997 ( .A1(cv[147]), .A2(n7122), .ZN(n7322) );
  NAND2_X1 U6998 ( .A1(n7322), .A2(n7321), .ZN(n7323) );
  INV_X8 U6999 ( .A(n7327), .ZN(n7384) );
  NAND2_X1 U7000 ( .A1(cv[148]), .A2(n7122), .ZN(n7326) );
  NAND2_X1 U7001 ( .A1(n7326), .A2(n7325), .ZN(n7327) );
  NAND2_X1 U7002 ( .A1(n7383), .A2(n6886), .ZN(cv_d[149]) );
  NAND2_X1 U7003 ( .A1(cv[149]), .A2(n7123), .ZN(n7330) );
  NAND2_X1 U7004 ( .A1(n7330), .A2(n7329), .ZN(n7331) );
  INV_X8 U7005 ( .A(n7339), .ZN(n7381) );
  NAND2_X1 U7006 ( .A1(cv[151]), .A2(n7123), .ZN(n7338) );
  NAND2_X1 U7007 ( .A1(n7338), .A2(n7337), .ZN(n7339) );
  INV_X8 U7008 ( .A(n7343), .ZN(n7380) );
  NAND2_X1 U7009 ( .A1(cv[152]), .A2(n7123), .ZN(n7342) );
  NAND2_X1 U7010 ( .A1(n7342), .A2(n7341), .ZN(n7343) );
  NAND2_X1 U7011 ( .A1(n7379), .A2(n6871), .ZN(cv_d[153]) );
  NAND2_X1 U7012 ( .A1(cv[153]), .A2(n7123), .ZN(n7346) );
  NAND2_X1 U7013 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
  NAND2_X1 U7014 ( .A1(n7378), .A2(n6868), .ZN(cv_d[154]) );
  NAND2_X1 U7015 ( .A1(cv[154]), .A2(n7123), .ZN(n7350) );
  NAND2_X1 U7016 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  INV_X1 U7017 ( .A(n7355), .ZN(n7377) );
  NAND2_X1 U7018 ( .A1(cv[155]), .A2(n7123), .ZN(n7354) );
  NAND2_X1 U7019 ( .A1(n7354), .A2(n7353), .ZN(n7355) );
  INV_X8 U7020 ( .A(n7359), .ZN(n7376) );
  NAND2_X1 U7021 ( .A1(cv[156]), .A2(n7123), .ZN(n7358) );
  NAND2_X1 U7022 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  INV_X8 U7023 ( .A(n7363), .ZN(n7375) );
  NAND2_X1 U7024 ( .A1(cv[157]), .A2(n7123), .ZN(n7362) );
  NAND2_X1 U7025 ( .A1(n7362), .A2(n7361), .ZN(n7363) );
  NAND2_X1 U7026 ( .A1(n7374), .A2(n6856), .ZN(cv_d[158]) );
  NAND2_X1 U7027 ( .A1(cv[158]), .A2(n7123), .ZN(n7366) );
  NAND2_X1 U7028 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  INV_X1 U7029 ( .A(n5906), .ZN(n7052) );
  INV_X4 U7030 ( .A(n7052), .ZN(n7053) );
  NAND2_X1 U7031 ( .A1(data_in[0]), .A2(n7228), .ZN(n5906) );
  NAND3_X1 U7032 ( .A1(n7053), .A2(n5907), .A3(n5908), .ZN(w_d[0]) );
  INV_X1 U7033 ( .A(n5673), .ZN(n7054) );
  INV_X4 U7034 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U7035 ( .A1(data_in[1]), .A2(n7228), .ZN(n5673) );
  NAND3_X1 U7036 ( .A1(n7055), .A2(n5674), .A3(n5675), .ZN(w_d[1]) );
  INV_X1 U7037 ( .A(n5440), .ZN(n7056) );
  INV_X4 U7038 ( .A(n7056), .ZN(n7057) );
  NAND2_X1 U7039 ( .A1(data_in[2]), .A2(n7229), .ZN(n5440) );
  NAND3_X1 U7040 ( .A1(n7057), .A2(n5441), .A3(n5442), .ZN(w_d[2]) );
  INV_X1 U7041 ( .A(n5215), .ZN(n7058) );
  INV_X4 U7042 ( .A(n7058), .ZN(n7059) );
  NAND2_X1 U7043 ( .A1(data_in[3]), .A2(n7229), .ZN(n5215) );
  NAND3_X1 U7044 ( .A1(n7059), .A2(n5216), .A3(n5217), .ZN(w_d[3]) );
  INV_X1 U7045 ( .A(n4829), .ZN(n7060) );
  INV_X4 U7046 ( .A(n7060), .ZN(n7061) );
  NAND2_X1 U7047 ( .A1(data_in[4]), .A2(n7229), .ZN(n4829) );
  NAND3_X1 U7048 ( .A1(n7061), .A2(n4830), .A3(n4831), .ZN(w_d[4]) );
  INV_X1 U7049 ( .A(n4686), .ZN(n7062) );
  INV_X4 U7050 ( .A(n7062), .ZN(n7063) );
  NAND2_X1 U7051 ( .A1(data_in[5]), .A2(n7229), .ZN(n4686) );
  NAND3_X1 U7052 ( .A1(n7063), .A2(n4687), .A3(n4688), .ZN(w_d[5]) );
  INV_X1 U7053 ( .A(n4675), .ZN(n7064) );
  INV_X4 U7054 ( .A(n7064), .ZN(n7065) );
  NAND2_X1 U7055 ( .A1(data_in[6]), .A2(n7229), .ZN(n4675) );
  NAND3_X1 U7056 ( .A1(n7065), .A2(n4676), .A3(n4677), .ZN(w_d[6]) );
  INV_X1 U7057 ( .A(n4672), .ZN(n7066) );
  INV_X4 U7058 ( .A(n7066), .ZN(n7067) );
  NAND2_X1 U7059 ( .A1(data_in[7]), .A2(n7229), .ZN(n4672) );
  NAND3_X1 U7060 ( .A1(n7067), .A2(n4673), .A3(n4674), .ZN(w_d[7]) );
  INV_X1 U7061 ( .A(n4669), .ZN(n7068) );
  INV_X4 U7062 ( .A(n7068), .ZN(n7069) );
  NAND2_X1 U7063 ( .A1(data_in[8]), .A2(n7229), .ZN(n4669) );
  NAND3_X1 U7064 ( .A1(n7069), .A2(n4670), .A3(n4671), .ZN(w_d[8]) );
  INV_X1 U7065 ( .A(n4654), .ZN(n7070) );
  INV_X4 U7066 ( .A(n7070), .ZN(n7071) );
  NAND2_X1 U7067 ( .A1(data_in[9]), .A2(n7227), .ZN(n4654) );
  NAND3_X1 U7068 ( .A1(n7071), .A2(n4655), .A3(n4656), .ZN(w_d[9]) );
  INV_X1 U7069 ( .A(n5883), .ZN(n7072) );
  INV_X4 U7070 ( .A(n7072), .ZN(n7073) );
  NAND2_X1 U7071 ( .A1(data_in[10]), .A2(n7227), .ZN(n5883) );
  NAND3_X1 U7072 ( .A1(n7073), .A2(n5884), .A3(n5885), .ZN(w_d[10]) );
  INV_X1 U7073 ( .A(n5860), .ZN(n7074) );
  INV_X4 U7074 ( .A(n7074), .ZN(n7075) );
  NAND2_X1 U7075 ( .A1(data_in[11]), .A2(n7227), .ZN(n5860) );
  NAND3_X1 U7076 ( .A1(n7075), .A2(n5861), .A3(n5862), .ZN(w_d[11]) );
  INV_X1 U7077 ( .A(n5837), .ZN(n7076) );
  INV_X4 U7078 ( .A(n7076), .ZN(n7077) );
  NAND2_X1 U7079 ( .A1(data_in[12]), .A2(n7227), .ZN(n5837) );
  NAND3_X1 U7080 ( .A1(n7077), .A2(n5838), .A3(n5839), .ZN(w_d[12]) );
  INV_X1 U7081 ( .A(n5814), .ZN(n7078) );
  INV_X4 U7082 ( .A(n7078), .ZN(n7079) );
  NAND2_X1 U7083 ( .A1(data_in[13]), .A2(n7227), .ZN(n5814) );
  NAND3_X1 U7084 ( .A1(n7079), .A2(n5815), .A3(n5816), .ZN(w_d[13]) );
  INV_X1 U7085 ( .A(n5791), .ZN(n7080) );
  INV_X4 U7086 ( .A(n7080), .ZN(n7081) );
  NAND2_X1 U7087 ( .A1(data_in[14]), .A2(n7227), .ZN(n5791) );
  NAND3_X1 U7088 ( .A1(n7081), .A2(n5792), .A3(n5793), .ZN(w_d[14]) );
  INV_X1 U7089 ( .A(n5768), .ZN(n7082) );
  INV_X4 U7090 ( .A(n7082), .ZN(n7083) );
  NAND2_X1 U7091 ( .A1(data_in[15]), .A2(n7227), .ZN(n5768) );
  NAND3_X1 U7092 ( .A1(n7083), .A2(n5769), .A3(n5770), .ZN(w_d[15]) );
  INV_X1 U7093 ( .A(n5745), .ZN(n7084) );
  INV_X4 U7094 ( .A(n7084), .ZN(n7085) );
  NAND2_X1 U7095 ( .A1(data_in[16]), .A2(n7227), .ZN(n5745) );
  NAND3_X1 U7096 ( .A1(n7085), .A2(n5746), .A3(n5747), .ZN(w_d[16]) );
  INV_X1 U7097 ( .A(n5722), .ZN(n7086) );
  INV_X4 U7098 ( .A(n7086), .ZN(n7087) );
  NAND2_X1 U7099 ( .A1(data_in[17]), .A2(n7227), .ZN(n5722) );
  NAND3_X1 U7100 ( .A1(n7087), .A2(n5723), .A3(n5724), .ZN(w_d[17]) );
  INV_X1 U7101 ( .A(n5699), .ZN(n7088) );
  INV_X4 U7102 ( .A(n7088), .ZN(n7089) );
  NAND2_X1 U7103 ( .A1(data_in[18]), .A2(n7227), .ZN(n5699) );
  NAND3_X1 U7104 ( .A1(n7089), .A2(n5700), .A3(n5701), .ZN(w_d[18]) );
  INV_X1 U7105 ( .A(n5676), .ZN(n7090) );
  INV_X4 U7106 ( .A(n7090), .ZN(n7091) );
  NAND2_X1 U7107 ( .A1(data_in[19]), .A2(n7227), .ZN(n5676) );
  NAND3_X1 U7108 ( .A1(n7091), .A2(n5677), .A3(n5678), .ZN(w_d[19]) );
  INV_X1 U7109 ( .A(n5650), .ZN(n7092) );
  INV_X4 U7110 ( .A(n7092), .ZN(n7093) );
  NAND2_X1 U7111 ( .A1(data_in[20]), .A2(n7228), .ZN(n5650) );
  NAND3_X1 U7112 ( .A1(n7093), .A2(n5651), .A3(n5652), .ZN(w_d[20]) );
  INV_X1 U7113 ( .A(n5627), .ZN(n7094) );
  INV_X4 U7114 ( .A(n7094), .ZN(n7095) );
  NAND2_X1 U7115 ( .A1(data_in[21]), .A2(n7228), .ZN(n5627) );
  NAND3_X1 U7116 ( .A1(n7095), .A2(n5628), .A3(n5629), .ZN(w_d[21]) );
  INV_X1 U7117 ( .A(n5604), .ZN(n7096) );
  INV_X4 U7118 ( .A(n7096), .ZN(n7097) );
  NAND2_X1 U7119 ( .A1(data_in[22]), .A2(n7228), .ZN(n5604) );
  NAND3_X1 U7120 ( .A1(n7097), .A2(n5605), .A3(n5606), .ZN(w_d[22]) );
  INV_X1 U7121 ( .A(n5581), .ZN(n7098) );
  INV_X4 U7122 ( .A(n7098), .ZN(n7099) );
  NAND2_X1 U7123 ( .A1(data_in[23]), .A2(n7228), .ZN(n5581) );
  NAND3_X1 U7124 ( .A1(n7099), .A2(n5582), .A3(n5583), .ZN(w_d[23]) );
  INV_X1 U7125 ( .A(n5558), .ZN(n7100) );
  INV_X4 U7126 ( .A(n7100), .ZN(n7101) );
  NAND2_X1 U7127 ( .A1(data_in[24]), .A2(n7228), .ZN(n5558) );
  NAND3_X1 U7128 ( .A1(n7101), .A2(n5559), .A3(n5560), .ZN(w_d[24]) );
  INV_X1 U7129 ( .A(n5535), .ZN(n7102) );
  INV_X4 U7130 ( .A(n7102), .ZN(n7103) );
  NAND2_X1 U7131 ( .A1(data_in[25]), .A2(n7228), .ZN(n5535) );
  NAND3_X1 U7132 ( .A1(n7103), .A2(n5536), .A3(n5537), .ZN(w_d[25]) );
  INV_X1 U7133 ( .A(n5512), .ZN(n7104) );
  INV_X4 U7134 ( .A(n7104), .ZN(n7105) );
  NAND2_X1 U7135 ( .A1(data_in[26]), .A2(n7228), .ZN(n5512) );
  NAND3_X1 U7136 ( .A1(n7105), .A2(n5513), .A3(n5514), .ZN(w_d[26]) );
  INV_X1 U7137 ( .A(n5489), .ZN(n7106) );
  INV_X4 U7138 ( .A(n7106), .ZN(n7107) );
  NAND2_X1 U7139 ( .A1(data_in[27]), .A2(n7228), .ZN(n5489) );
  NAND3_X1 U7140 ( .A1(n7107), .A2(n5490), .A3(n5491), .ZN(w_d[27]) );
  INV_X1 U7141 ( .A(n5466), .ZN(n7108) );
  INV_X4 U7142 ( .A(n7108), .ZN(n7109) );
  NAND2_X1 U7143 ( .A1(data_in[28]), .A2(n7228), .ZN(n5466) );
  NAND3_X1 U7144 ( .A1(n7109), .A2(n5467), .A3(n5468), .ZN(w_d[28]) );
  INV_X1 U7145 ( .A(n5443), .ZN(n7110) );
  INV_X4 U7146 ( .A(n7110), .ZN(n7111) );
  NAND2_X1 U7147 ( .A1(data_in[29]), .A2(n7229), .ZN(n5443) );
  NAND3_X1 U7148 ( .A1(n7111), .A2(n5444), .A3(n5445), .ZN(w_d[29]) );
  INV_X1 U7149 ( .A(n5417), .ZN(n7112) );
  INV_X4 U7150 ( .A(n7112), .ZN(n7113) );
  NAND2_X1 U7151 ( .A1(data_in[30]), .A2(n7229), .ZN(n5417) );
  NAND3_X1 U7152 ( .A1(n7113), .A2(n5418), .A3(n5419), .ZN(w_d[30]) );
  INV_X1 U7153 ( .A(n5394), .ZN(n7114) );
  INV_X4 U7154 ( .A(n7114), .ZN(n7115) );
  NAND2_X1 U7155 ( .A1(data_in[31]), .A2(n7229), .ZN(n5394) );
  NAND3_X1 U7156 ( .A1(n7115), .A2(n5395), .A3(n5396), .ZN(w_d[31]) );
  CLKBUF_X1 U7157 ( .A(start), .Z(n7116) );
  CLKBUF_X1 U7158 ( .A(reset), .Z(n7117) );
  NOR2_X1 U7159 ( .A1(n7116), .A2(n6243), .ZN(next_state[1]) );
  INV_X1 U7160 ( .A(n7371), .ZN(n7373) );
  NAND2_X1 U7161 ( .A1(cv[159]), .A2(n7123), .ZN(n7370) );
  NAND2_X1 U7162 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  INV_X8 U7163 ( .A(n7335), .ZN(n7382) );
  NAND2_X1 U7164 ( .A1(cv[150]), .A2(n7123), .ZN(n7334) );
  NAND2_X1 U7165 ( .A1(n7334), .A2(n7333), .ZN(n7335) );
  INV_X1 U7166 ( .A(rnd_cnt_q[5]), .ZN(n7398) );
  XNOR2_X1 U7167 ( .A(rnd_cnt_q[6]), .B(n6231), .ZN(n6229) );
  NAND4_X1 U7168 ( .A1(rnd_cnt_q[6]), .A2(n5038), .A3(n7399), .A4(n7398), .ZN(
        n6245) );
  NAND2_X1 U7169 ( .A1(w[11]), .A2(n7238), .ZN(n4922) );
  BUF_X4 U7170 ( .A(n4662), .Z(n7193) );
  BUF_X4 U7171 ( .A(n4662), .Z(n7194) );
  BUF_X4 U7172 ( .A(n4662), .Z(n7211) );
  BUF_X4 U7173 ( .A(n4662), .Z(n7215) );
  BUF_X4 U7174 ( .A(n7226), .Z(n7182) );
  BUF_X4 U7175 ( .A(n7225), .Z(n7183) );
  BUF_X4 U7176 ( .A(n7225), .Z(n7184) );
  BUF_X4 U7177 ( .A(n7225), .Z(n7185) );
  BUF_X4 U7178 ( .A(n7224), .Z(n7186) );
  BUF_X4 U7179 ( .A(n7224), .Z(n7187) );
  BUF_X4 U7180 ( .A(n7224), .Z(n7188) );
  BUF_X4 U7181 ( .A(n7223), .Z(n7189) );
  BUF_X4 U7182 ( .A(n7223), .Z(n7190) );
  BUF_X4 U7183 ( .A(n7223), .Z(n7191) );
  BUF_X4 U7184 ( .A(n4662), .Z(n7192) );
  BUF_X4 U7185 ( .A(n4662), .Z(n7195) );
  BUF_X4 U7186 ( .A(n7226), .Z(n7196) );
  BUF_X4 U7187 ( .A(n7188), .Z(n7197) );
  BUF_X4 U7188 ( .A(n7222), .Z(n7198) );
  BUF_X4 U7189 ( .A(n7222), .Z(n7199) );
  BUF_X4 U7190 ( .A(n7222), .Z(n7200) );
  BUF_X4 U7191 ( .A(n7221), .Z(n7201) );
  BUF_X4 U7192 ( .A(n7221), .Z(n7202) );
  BUF_X4 U7193 ( .A(n7221), .Z(n7203) );
  BUF_X4 U7194 ( .A(n7220), .Z(n7204) );
  BUF_X4 U7195 ( .A(n7220), .Z(n7205) );
  BUF_X4 U7196 ( .A(n7220), .Z(n7206) );
  BUF_X4 U7197 ( .A(n7219), .Z(n7207) );
  BUF_X4 U7198 ( .A(n7219), .Z(n7208) );
  BUF_X4 U7199 ( .A(n7219), .Z(n7209) );
  BUF_X4 U7200 ( .A(n4662), .Z(n7210) );
  BUF_X4 U7201 ( .A(n7218), .Z(n7212) );
  BUF_X4 U7202 ( .A(n7218), .Z(n7213) );
  BUF_X4 U7203 ( .A(n7217), .Z(n7214) );
  BUF_X4 U7204 ( .A(n7196), .Z(n7216) );
  BUF_X4 U7205 ( .A(n4662), .Z(n7217) );
  BUF_X4 U7206 ( .A(n4662), .Z(n7225) );
  BUF_X4 U7207 ( .A(n4662), .Z(n7224) );
  BUF_X4 U7208 ( .A(n4662), .Z(n7223) );
  BUF_X4 U7209 ( .A(n4662), .Z(n7222) );
  BUF_X4 U7210 ( .A(n4662), .Z(n7221) );
  BUF_X4 U7211 ( .A(n4662), .Z(n7220) );
  BUF_X4 U7212 ( .A(n4662), .Z(n7219) );
  BUF_X4 U7213 ( .A(n4662), .Z(n7218) );
  BUF_X4 U7214 ( .A(n4662), .Z(n7226) );
  INV_X4 U7215 ( .A(n7395), .ZN(n7152) );
  INV_X4 U7216 ( .A(n7166), .ZN(n7165) );
  INV_X4 U7217 ( .A(n7166), .ZN(n7163) );
  INV_X4 U7218 ( .A(n7166), .ZN(n7161) );
  INV_X4 U7219 ( .A(n7166), .ZN(n7164) );
  INV_X4 U7220 ( .A(n7166), .ZN(n7162) );
  INV_X4 U7221 ( .A(n7166), .ZN(n7158) );
  INV_X4 U7222 ( .A(n7166), .ZN(n7157) );
  INV_X4 U7223 ( .A(n7166), .ZN(n7160) );
  INV_X4 U7224 ( .A(n7166), .ZN(n7159) );
  INV_X4 U7225 ( .A(n7166), .ZN(n7155) );
  INV_X4 U7226 ( .A(n7166), .ZN(n7154) );
  INV_X4 U7227 ( .A(n7166), .ZN(n7156) );
  INV_X4 U7228 ( .A(n7395), .ZN(n7153) );
  INV_X4 U7229 ( .A(n6248), .ZN(n7176) );
  INV_X4 U7230 ( .A(n6248), .ZN(n7175) );
  INV_X4 U7231 ( .A(n6248), .ZN(n7174) );
  INV_X4 U7232 ( .A(n6248), .ZN(n7173) );
  INV_X4 U7233 ( .A(n6248), .ZN(n7171) );
  INV_X4 U7234 ( .A(n6248), .ZN(n7170) );
  INV_X4 U7235 ( .A(n6248), .ZN(n7172) );
  INV_X4 U7236 ( .A(n6248), .ZN(n7169) );
  INV_X4 U7237 ( .A(n7153), .ZN(n7166) );
  INV_X4 U7238 ( .A(n6248), .ZN(n7168) );
  INV_X4 U7239 ( .A(n6248), .ZN(n7167) );
  INV_X4 U7240 ( .A(n7283), .ZN(n7131) );
  INV_X4 U7241 ( .A(n7284), .ZN(n7146) );
  INV_X4 U7242 ( .A(n7283), .ZN(n7130) );
  INV_X4 U7243 ( .A(n7284), .ZN(n7145) );
  INV_X4 U7244 ( .A(n7283), .ZN(n7129) );
  INV_X4 U7245 ( .A(n7284), .ZN(n7144) );
  INV_X4 U7246 ( .A(n7283), .ZN(n7128) );
  INV_X4 U7247 ( .A(n7284), .ZN(n7143) );
  INV_X4 U7248 ( .A(n7283), .ZN(n7135) );
  INV_X4 U7249 ( .A(n7284), .ZN(n7150) );
  INV_X4 U7250 ( .A(n7283), .ZN(n7134) );
  INV_X4 U7251 ( .A(n7284), .ZN(n7149) );
  INV_X4 U7252 ( .A(n7283), .ZN(n7133) );
  INV_X4 U7253 ( .A(n7284), .ZN(n7148) );
  INV_X4 U7254 ( .A(n7283), .ZN(n7132) );
  INV_X4 U7255 ( .A(n7284), .ZN(n7147) );
  INV_X4 U7256 ( .A(n7284), .ZN(n7137) );
  INV_X4 U7257 ( .A(n7283), .ZN(n7122) );
  INV_X4 U7258 ( .A(n7284), .ZN(n7138) );
  INV_X4 U7259 ( .A(n7283), .ZN(n7123) );
  INV_X4 U7260 ( .A(n7283), .ZN(n7127) );
  INV_X4 U7261 ( .A(n7284), .ZN(n7142) );
  INV_X4 U7262 ( .A(n7283), .ZN(n7126) );
  INV_X4 U7263 ( .A(n7284), .ZN(n7141) );
  INV_X4 U7264 ( .A(n7283), .ZN(n7125) );
  INV_X4 U7265 ( .A(n7284), .ZN(n7140) );
  INV_X4 U7266 ( .A(n7283), .ZN(n7124) );
  INV_X4 U7267 ( .A(n7284), .ZN(n7139) );
  INV_X4 U7268 ( .A(n7283), .ZN(n7136) );
  INV_X4 U7269 ( .A(n7284), .ZN(n7151) );
  BUF_X4 U7270 ( .A(n7237), .Z(n7269) );
  BUF_X4 U7271 ( .A(n4658), .Z(n7270) );
  BUF_X4 U7272 ( .A(n7237), .Z(n7271) );
  BUF_X4 U7273 ( .A(n7237), .Z(n7276) );
  BUF_X4 U7274 ( .A(n7237), .Z(n7277) );
  BUF_X4 U7275 ( .A(n7238), .Z(n7278) );
  BUF_X4 U7276 ( .A(n7279), .Z(n7239) );
  BUF_X4 U7277 ( .A(n7279), .Z(n7240) );
  BUF_X4 U7278 ( .A(n7279), .Z(n7241) );
  BUF_X4 U7279 ( .A(n7230), .Z(n7242) );
  BUF_X4 U7280 ( .A(n7230), .Z(n7243) );
  BUF_X4 U7281 ( .A(n7230), .Z(n7244) );
  BUF_X4 U7282 ( .A(n7231), .Z(n7245) );
  BUF_X4 U7283 ( .A(n7231), .Z(n7246) );
  BUF_X4 U7284 ( .A(n7231), .Z(n7247) );
  BUF_X4 U7285 ( .A(n7232), .Z(n7248) );
  BUF_X4 U7286 ( .A(n7232), .Z(n7249) );
  BUF_X4 U7287 ( .A(n7232), .Z(n7250) );
  BUF_X4 U7288 ( .A(n4658), .Z(n7251) );
  BUF_X4 U7289 ( .A(n7237), .Z(n7252) );
  BUF_X4 U7290 ( .A(n7267), .Z(n7253) );
  BUF_X4 U7291 ( .A(n7274), .Z(n7254) );
  BUF_X4 U7292 ( .A(n7233), .Z(n7255) );
  BUF_X4 U7293 ( .A(n7233), .Z(n7256) );
  BUF_X4 U7294 ( .A(n7233), .Z(n7257) );
  BUF_X4 U7295 ( .A(n7234), .Z(n7258) );
  BUF_X4 U7296 ( .A(n7234), .Z(n7259) );
  BUF_X4 U7297 ( .A(n7234), .Z(n7260) );
  BUF_X4 U7298 ( .A(n7235), .Z(n7261) );
  BUF_X4 U7299 ( .A(n7235), .Z(n7262) );
  BUF_X4 U7300 ( .A(n7235), .Z(n7263) );
  BUF_X4 U7301 ( .A(n7236), .Z(n7264) );
  BUF_X4 U7302 ( .A(n7236), .Z(n7265) );
  BUF_X4 U7303 ( .A(n7236), .Z(n7266) );
  BUF_X4 U7304 ( .A(n7236), .Z(n7267) );
  BUF_X4 U7305 ( .A(n4658), .Z(n7268) );
  BUF_X4 U7306 ( .A(n7237), .Z(n7272) );
  BUF_X4 U7307 ( .A(n7237), .Z(n7273) );
  BUF_X4 U7308 ( .A(n7237), .Z(n7274) );
  BUF_X4 U7309 ( .A(n7237), .Z(n7275) );
  BUF_X4 U7310 ( .A(n7238), .Z(n7279) );
  INV_X4 U7311 ( .A(n7120), .ZN(n7229) );
  INV_X4 U7312 ( .A(n7120), .ZN(n7227) );
  INV_X4 U7313 ( .A(n7120), .ZN(n7228) );
  INV_X4 U7314 ( .A(n7181), .ZN(n7177) );
  INV_X4 U7315 ( .A(n7181), .ZN(n7178) );
  INV_X4 U7316 ( .A(n7181), .ZN(n7179) );
  BUF_X4 U7317 ( .A(n4658), .Z(n7230) );
  BUF_X4 U7318 ( .A(n4658), .Z(n7231) );
  BUF_X4 U7319 ( .A(n4658), .Z(n7232) );
  BUF_X4 U7320 ( .A(n4658), .Z(n7233) );
  BUF_X4 U7321 ( .A(n4658), .Z(n7234) );
  BUF_X4 U7322 ( .A(n4658), .Z(n7235) );
  BUF_X4 U7323 ( .A(n4658), .Z(n7236) );
  BUF_X4 U7324 ( .A(n4658), .Z(n7237) );
  BUF_X4 U7325 ( .A(n4658), .Z(n7238) );
  OR2_X2 U7326 ( .A1(n7403), .A2(n7152), .ZN(n7120) );
  NAND3_X2 U7327 ( .A1(n6245), .A2(n7402), .A3(n7152), .ZN(n6230) );
  INV_X4 U7328 ( .A(n7121), .ZN(n7180) );
  NOR2_X2 U7329 ( .A1(n6233), .A2(n6230), .ZN(rnd_cnt_d[5]) );
  NOR2_X2 U7330 ( .A1(n6234), .A2(n6230), .ZN(rnd_cnt_d[4]) );
  INV_X4 U7331 ( .A(n7121), .ZN(n7181) );
  NOR2_X2 U7332 ( .A1(n7152), .A2(load_in), .ZN(n4658) );
  NOR2_X2 U7333 ( .A1(n6230), .A2(rnd_cnt_q[0]), .ZN(rnd_cnt_d[0]) );
  AND2_X2 U7334 ( .A1(n5037), .A2(n7403), .ZN(n7121) );
  NOR2_X2 U7335 ( .A1(n6244), .A2(n7167), .ZN(n6243) );
  NOR2_X2 U7336 ( .A1(n7395), .A2(n6245), .ZN(n6244) );
  NAND3_X2 U7337 ( .A1(n6246), .A2(n6230), .A3(n6247), .ZN(next_state[0]) );
  NAND3_X2 U7338 ( .A1(n6248), .A2(n7395), .A3(n7116), .ZN(n6246) );
  NAND3_X2 U7339 ( .A1(rnd_cnt_q[0]), .A2(n7401), .A3(n7396), .ZN(n6242) );
  NOR2_X2 U7340 ( .A1(n6229), .A2(n6230), .ZN(rnd_cnt_d[6]) );
  NOR2_X2 U7341 ( .A1(n6232), .A2(n7398), .ZN(n6231) );
  NOR2_X2 U7342 ( .A1(n6235), .A2(n6230), .ZN(rnd_cnt_d[3]) );
  XNOR2_X1 U7343 ( .A(n6236), .B(rnd_cnt_q[3]), .ZN(n6235) );
  INV_X1 U7344 ( .A(n7119), .ZN(n7400) );
  INV_X1 U7345 ( .A(rnd_cnt_q[4]), .ZN(n7399) );
  NAND2_X1 U7346 ( .A1(n7119), .A2(n6239), .ZN(n6237) );
  AND3_X4 U7347 ( .A1(rnd_cnt_q[1]), .A2(rnd_cnt_q[0]), .A3(n7119), .ZN(n6236)
         );
  XNOR2_X1 U7348 ( .A(rnd_cnt_q[4]), .B(n5038), .ZN(n6234) );
  NAND2_X1 U7349 ( .A1(rnd_cnt_q[4]), .A2(n5038), .ZN(n6232) );
  OR4_X1 U7350 ( .A1(n5038), .A2(rnd_cnt_q[4]), .A3(rnd_cnt_q[5]), .A4(
        rnd_cnt_q[6]), .ZN(n5037) );
  OR2_X4 U7351 ( .A1(n7165), .A2(n7229), .ZN(n4662) );
  INV_X4 U7352 ( .A(state[0]), .ZN(n7280) );
  NAND2_X2 U7353 ( .A1(state[1]), .A2(n7280), .ZN(n6248) );
  MUX2_X2 U7354 ( .A(cv_next[0]), .B(N157), .S(n7167), .Z(cv_next_d[0]) );
  MUX2_X2 U7355 ( .A(cv_next[1]), .B(N158), .S(n7168), .Z(cv_next_d[1]) );
  MUX2_X2 U7356 ( .A(cv_next[2]), .B(N159), .S(n7167), .Z(cv_next_d[2]) );
  MUX2_X2 U7357 ( .A(cv_next[3]), .B(N160), .S(n7176), .Z(cv_next_d[3]) );
  MUX2_X2 U7358 ( .A(cv_next[4]), .B(N161), .S(n7176), .Z(cv_next_d[4]) );
  MUX2_X2 U7359 ( .A(cv_next[5]), .B(N162), .S(n7176), .Z(cv_next_d[5]) );
  MUX2_X2 U7360 ( .A(cv_next[6]), .B(N163), .S(n7176), .Z(cv_next_d[6]) );
  MUX2_X2 U7361 ( .A(cv_next[7]), .B(N164), .S(n7176), .Z(cv_next_d[7]) );
  MUX2_X2 U7362 ( .A(cv_next[8]), .B(N165), .S(n7176), .Z(cv_next_d[8]) );
  MUX2_X2 U7363 ( .A(cv_next[9]), .B(N166), .S(n7176), .Z(cv_next_d[9]) );
  MUX2_X2 U7364 ( .A(cv_next[10]), .B(N167), .S(n7176), .Z(cv_next_d[10]) );
  MUX2_X2 U7365 ( .A(cv_next[11]), .B(N168), .S(n7176), .Z(cv_next_d[11]) );
  MUX2_X2 U7366 ( .A(cv_next[12]), .B(N169), .S(n7176), .Z(cv_next_d[12]) );
  MUX2_X2 U7367 ( .A(cv_next[13]), .B(N170), .S(n7176), .Z(cv_next_d[13]) );
  MUX2_X2 U7368 ( .A(cv_next[14]), .B(N171), .S(n7176), .Z(cv_next_d[14]) );
  MUX2_X2 U7369 ( .A(cv_next[15]), .B(N172), .S(n7176), .Z(cv_next_d[15]) );
  MUX2_X2 U7370 ( .A(cv_next[16]), .B(N173), .S(n7176), .Z(cv_next_d[16]) );
  MUX2_X2 U7371 ( .A(cv_next[17]), .B(N174), .S(n7176), .Z(cv_next_d[17]) );
  MUX2_X2 U7372 ( .A(cv_next[18]), .B(N175), .S(n7176), .Z(cv_next_d[18]) );
  MUX2_X2 U7373 ( .A(cv_next[19]), .B(N176), .S(n7175), .Z(cv_next_d[19]) );
  MUX2_X2 U7374 ( .A(cv_next[20]), .B(N177), .S(n7175), .Z(cv_next_d[20]) );
  MUX2_X2 U7375 ( .A(cv_next[21]), .B(N178), .S(n7175), .Z(cv_next_d[21]) );
  MUX2_X2 U7376 ( .A(cv_next[22]), .B(N179), .S(n7175), .Z(cv_next_d[22]) );
  MUX2_X2 U7377 ( .A(cv_next[23]), .B(N180), .S(n7175), .Z(cv_next_d[23]) );
  MUX2_X2 U7378 ( .A(cv_next[24]), .B(N181), .S(n7175), .Z(cv_next_d[24]) );
  MUX2_X2 U7379 ( .A(cv_next[25]), .B(N182), .S(n7175), .Z(cv_next_d[25]) );
  MUX2_X2 U7380 ( .A(cv_next[26]), .B(N183), .S(n7175), .Z(cv_next_d[26]) );
  MUX2_X2 U7381 ( .A(cv_next[27]), .B(N184), .S(n7175), .Z(cv_next_d[27]) );
  MUX2_X2 U7382 ( .A(cv_next[28]), .B(N185), .S(n7175), .Z(cv_next_d[28]) );
  MUX2_X2 U7383 ( .A(cv_next[29]), .B(N186), .S(n7175), .Z(cv_next_d[29]) );
  MUX2_X2 U7384 ( .A(cv_next[30]), .B(N187), .S(n7175), .Z(cv_next_d[30]) );
  MUX2_X2 U7385 ( .A(cv_next[31]), .B(N188), .S(n7175), .Z(cv_next_d[31]) );
  MUX2_X2 U7386 ( .A(cv_next[32]), .B(N125), .S(n7175), .Z(cv_next_d[32]) );
  MUX2_X2 U7387 ( .A(cv_next[33]), .B(N126), .S(n7175), .Z(cv_next_d[33]) );
  MUX2_X2 U7388 ( .A(cv_next[34]), .B(N127), .S(n7175), .Z(cv_next_d[34]) );
  MUX2_X2 U7389 ( .A(cv_next[35]), .B(N128), .S(n7174), .Z(cv_next_d[35]) );
  MUX2_X2 U7390 ( .A(cv_next[36]), .B(N129), .S(n7174), .Z(cv_next_d[36]) );
  MUX2_X2 U7391 ( .A(cv_next[37]), .B(N130), .S(n7174), .Z(cv_next_d[37]) );
  MUX2_X2 U7392 ( .A(cv_next[38]), .B(N131), .S(n7174), .Z(cv_next_d[38]) );
  MUX2_X2 U7393 ( .A(cv_next[39]), .B(N132), .S(n7174), .Z(cv_next_d[39]) );
  MUX2_X2 U7394 ( .A(cv_next[40]), .B(N133), .S(n7174), .Z(cv_next_d[40]) );
  MUX2_X2 U7395 ( .A(cv_next[41]), .B(N134), .S(n7174), .Z(cv_next_d[41]) );
  MUX2_X2 U7396 ( .A(cv_next[42]), .B(N135), .S(n7174), .Z(cv_next_d[42]) );
  MUX2_X2 U7397 ( .A(cv_next[43]), .B(N136), .S(n7174), .Z(cv_next_d[43]) );
  MUX2_X2 U7398 ( .A(cv_next[44]), .B(N137), .S(n7174), .Z(cv_next_d[44]) );
  MUX2_X2 U7399 ( .A(cv_next[45]), .B(N138), .S(n7174), .Z(cv_next_d[45]) );
  MUX2_X2 U7400 ( .A(cv_next[46]), .B(N139), .S(n7174), .Z(cv_next_d[46]) );
  MUX2_X2 U7401 ( .A(cv_next[47]), .B(N140), .S(n7174), .Z(cv_next_d[47]) );
  MUX2_X2 U7402 ( .A(cv_next[48]), .B(N141), .S(n7174), .Z(cv_next_d[48]) );
  MUX2_X2 U7403 ( .A(cv_next[49]), .B(N142), .S(n7174), .Z(cv_next_d[49]) );
  MUX2_X2 U7404 ( .A(cv_next[50]), .B(N143), .S(n7174), .Z(cv_next_d[50]) );
  MUX2_X2 U7405 ( .A(cv_next[51]), .B(N144), .S(n7173), .Z(cv_next_d[51]) );
  MUX2_X2 U7406 ( .A(cv_next[52]), .B(N145), .S(n7173), .Z(cv_next_d[52]) );
  MUX2_X2 U7407 ( .A(cv_next[53]), .B(N146), .S(n7173), .Z(cv_next_d[53]) );
  MUX2_X2 U7408 ( .A(cv_next[54]), .B(N147), .S(n7173), .Z(cv_next_d[54]) );
  MUX2_X2 U7409 ( .A(cv_next[55]), .B(N148), .S(n7173), .Z(cv_next_d[55]) );
  MUX2_X2 U7410 ( .A(cv_next[56]), .B(N149), .S(n7173), .Z(cv_next_d[56]) );
  MUX2_X2 U7411 ( .A(cv_next[57]), .B(N150), .S(n7173), .Z(cv_next_d[57]) );
  MUX2_X2 U7412 ( .A(cv_next[58]), .B(N151), .S(n7173), .Z(cv_next_d[58]) );
  MUX2_X2 U7413 ( .A(cv_next[59]), .B(N152), .S(n7173), .Z(cv_next_d[59]) );
  MUX2_X2 U7414 ( .A(cv_next[60]), .B(N153), .S(n7173), .Z(cv_next_d[60]) );
  MUX2_X2 U7415 ( .A(cv_next[61]), .B(N154), .S(n7173), .Z(cv_next_d[61]) );
  MUX2_X2 U7416 ( .A(cv_next[62]), .B(N155), .S(n7173), .Z(cv_next_d[62]) );
  MUX2_X2 U7417 ( .A(cv_next[63]), .B(N156), .S(n7173), .Z(cv_next_d[63]) );
  MUX2_X2 U7418 ( .A(cv_next[64]), .B(N93), .S(n7173), .Z(cv_next_d[64]) );
  MUX2_X2 U7419 ( .A(cv_next[65]), .B(N94), .S(n7173), .Z(cv_next_d[65]) );
  MUX2_X2 U7420 ( .A(cv_next[66]), .B(N95), .S(n7173), .Z(cv_next_d[66]) );
  MUX2_X2 U7421 ( .A(cv_next[67]), .B(N96), .S(n7172), .Z(cv_next_d[67]) );
  MUX2_X2 U7422 ( .A(cv_next[68]), .B(N97), .S(n7172), .Z(cv_next_d[68]) );
  MUX2_X2 U7423 ( .A(cv_next[69]), .B(N98), .S(n7172), .Z(cv_next_d[69]) );
  MUX2_X2 U7424 ( .A(cv_next[70]), .B(N99), .S(n7172), .Z(cv_next_d[70]) );
  MUX2_X2 U7425 ( .A(cv_next[71]), .B(N100), .S(n7172), .Z(cv_next_d[71]) );
  MUX2_X2 U7426 ( .A(cv_next[72]), .B(N101), .S(n7172), .Z(cv_next_d[72]) );
  MUX2_X2 U7427 ( .A(cv_next[73]), .B(N102), .S(n7172), .Z(cv_next_d[73]) );
  MUX2_X2 U7428 ( .A(cv_next[74]), .B(N103), .S(n7172), .Z(cv_next_d[74]) );
  MUX2_X2 U7429 ( .A(cv_next[75]), .B(N104), .S(n7172), .Z(cv_next_d[75]) );
  MUX2_X2 U7430 ( .A(cv_next[76]), .B(N105), .S(n7172), .Z(cv_next_d[76]) );
  MUX2_X2 U7431 ( .A(cv_next[77]), .B(N106), .S(n7172), .Z(cv_next_d[77]) );
  MUX2_X2 U7432 ( .A(cv_next[78]), .B(N107), .S(n7172), .Z(cv_next_d[78]) );
  MUX2_X2 U7433 ( .A(cv_next[79]), .B(N108), .S(n7172), .Z(cv_next_d[79]) );
  MUX2_X2 U7434 ( .A(cv_next[80]), .B(N109), .S(n7172), .Z(cv_next_d[80]) );
  MUX2_X2 U7435 ( .A(cv_next[81]), .B(N110), .S(n7172), .Z(cv_next_d[81]) );
  MUX2_X2 U7436 ( .A(cv_next[82]), .B(N111), .S(n7171), .Z(cv_next_d[82]) );
  MUX2_X2 U7437 ( .A(cv_next[83]), .B(N112), .S(n7171), .Z(cv_next_d[83]) );
  MUX2_X2 U7438 ( .A(cv_next[84]), .B(N113), .S(n7171), .Z(cv_next_d[84]) );
  MUX2_X2 U7439 ( .A(cv_next[85]), .B(N114), .S(n7171), .Z(cv_next_d[85]) );
  MUX2_X2 U7440 ( .A(cv_next[86]), .B(N115), .S(n7171), .Z(cv_next_d[86]) );
  MUX2_X2 U7441 ( .A(cv_next[87]), .B(N116), .S(n7171), .Z(cv_next_d[87]) );
  MUX2_X2 U7442 ( .A(cv_next[88]), .B(N117), .S(n7171), .Z(cv_next_d[88]) );
  MUX2_X2 U7443 ( .A(cv_next[89]), .B(N118), .S(n7171), .Z(cv_next_d[89]) );
  MUX2_X2 U7444 ( .A(cv_next[90]), .B(N119), .S(n7171), .Z(cv_next_d[90]) );
  MUX2_X2 U7445 ( .A(cv_next[91]), .B(N120), .S(n7171), .Z(cv_next_d[91]) );
  MUX2_X2 U7446 ( .A(cv_next[92]), .B(N121), .S(n7171), .Z(cv_next_d[92]) );
  MUX2_X2 U7447 ( .A(cv_next[93]), .B(N122), .S(n7171), .Z(cv_next_d[93]) );
  MUX2_X2 U7448 ( .A(cv_next[94]), .B(N123), .S(n7171), .Z(cv_next_d[94]) );
  MUX2_X2 U7449 ( .A(cv_next[95]), .B(N124), .S(n7171), .Z(cv_next_d[95]) );
  MUX2_X2 U7450 ( .A(cv_next[96]), .B(N61), .S(n7171), .Z(cv_next_d[96]) );
  MUX2_X2 U7451 ( .A(cv_next[97]), .B(N62), .S(n7171), .Z(cv_next_d[97]) );
  MUX2_X2 U7452 ( .A(cv_next[98]), .B(N63), .S(n7170), .Z(cv_next_d[98]) );
  MUX2_X2 U7453 ( .A(cv_next[99]), .B(N64), .S(n7170), .Z(cv_next_d[99]) );
  MUX2_X2 U7454 ( .A(cv_next[100]), .B(N65), .S(n7170), .Z(cv_next_d[100]) );
  MUX2_X2 U7455 ( .A(cv_next[101]), .B(N66), .S(n7170), .Z(cv_next_d[101]) );
  MUX2_X2 U7456 ( .A(cv_next[102]), .B(N67), .S(n7170), .Z(cv_next_d[102]) );
  MUX2_X2 U7457 ( .A(cv_next[103]), .B(N68), .S(n7170), .Z(cv_next_d[103]) );
  MUX2_X2 U7458 ( .A(cv_next[104]), .B(N69), .S(n7170), .Z(cv_next_d[104]) );
  MUX2_X2 U7459 ( .A(cv_next[105]), .B(N70), .S(n7170), .Z(cv_next_d[105]) );
  MUX2_X2 U7460 ( .A(cv_next[106]), .B(N71), .S(n7170), .Z(cv_next_d[106]) );
  MUX2_X2 U7461 ( .A(cv_next[107]), .B(N72), .S(n7170), .Z(cv_next_d[107]) );
  MUX2_X2 U7462 ( .A(cv_next[108]), .B(N73), .S(n7170), .Z(cv_next_d[108]) );
  MUX2_X2 U7463 ( .A(cv_next[109]), .B(N74), .S(n7170), .Z(cv_next_d[109]) );
  MUX2_X2 U7464 ( .A(cv_next[110]), .B(N75), .S(n7170), .Z(cv_next_d[110]) );
  MUX2_X2 U7465 ( .A(cv_next[111]), .B(N76), .S(n7170), .Z(cv_next_d[111]) );
  MUX2_X2 U7466 ( .A(cv_next[112]), .B(N77), .S(n7170), .Z(cv_next_d[112]) );
  MUX2_X2 U7467 ( .A(cv_next[113]), .B(N78), .S(n7170), .Z(cv_next_d[113]) );
  MUX2_X2 U7468 ( .A(cv_next[114]), .B(N79), .S(n7169), .Z(cv_next_d[114]) );
  MUX2_X2 U7469 ( .A(cv_next[115]), .B(N80), .S(n7169), .Z(cv_next_d[115]) );
  MUX2_X2 U7470 ( .A(cv_next[116]), .B(N81), .S(n7169), .Z(cv_next_d[116]) );
  MUX2_X2 U7471 ( .A(cv_next[117]), .B(N82), .S(n7169), .Z(cv_next_d[117]) );
  MUX2_X2 U7472 ( .A(cv_next[118]), .B(N83), .S(n7169), .Z(cv_next_d[118]) );
  MUX2_X2 U7473 ( .A(cv_next[119]), .B(N84), .S(n7169), .Z(cv_next_d[119]) );
  MUX2_X2 U7474 ( .A(cv_next[120]), .B(N85), .S(n7169), .Z(cv_next_d[120]) );
  MUX2_X2 U7475 ( .A(cv_next[121]), .B(N86), .S(n7172), .Z(cv_next_d[121]) );
  MUX2_X2 U7476 ( .A(cv_next[122]), .B(N87), .S(n7169), .Z(cv_next_d[122]) );
  MUX2_X2 U7477 ( .A(cv_next[123]), .B(N88), .S(n7169), .Z(cv_next_d[123]) );
  MUX2_X2 U7478 ( .A(cv_next[124]), .B(N89), .S(n7169), .Z(cv_next_d[124]) );
  MUX2_X2 U7479 ( .A(cv_next[125]), .B(N90), .S(n7169), .Z(cv_next_d[125]) );
  MUX2_X2 U7480 ( .A(cv_next[126]), .B(N91), .S(n7169), .Z(cv_next_d[126]) );
  MUX2_X2 U7481 ( .A(cv_next[127]), .B(N92), .S(n7169), .Z(cv_next_d[127]) );
  MUX2_X2 U7482 ( .A(cv_next[128]), .B(N29), .S(n7169), .Z(cv_next_d[128]) );
  MUX2_X2 U7483 ( .A(cv_next[129]), .B(N30), .S(n7169), .Z(cv_next_d[129]) );
  MUX2_X2 U7484 ( .A(cv_next[130]), .B(N31), .S(n7169), .Z(cv_next_d[130]) );
  MUX2_X2 U7485 ( .A(cv_next[131]), .B(N32), .S(n7168), .Z(cv_next_d[131]) );
  MUX2_X2 U7486 ( .A(cv_next[132]), .B(N33), .S(n7168), .Z(cv_next_d[132]) );
  MUX2_X2 U7487 ( .A(cv_next[133]), .B(N34), .S(n7168), .Z(cv_next_d[133]) );
  MUX2_X2 U7488 ( .A(cv_next[134]), .B(N35), .S(n7168), .Z(cv_next_d[134]) );
  MUX2_X2 U7489 ( .A(cv_next[135]), .B(N36), .S(n7168), .Z(cv_next_d[135]) );
  MUX2_X2 U7490 ( .A(cv_next[136]), .B(N37), .S(n7168), .Z(cv_next_d[136]) );
  MUX2_X2 U7491 ( .A(cv_next[137]), .B(N38), .S(n7168), .Z(cv_next_d[137]) );
  MUX2_X2 U7492 ( .A(cv_next[138]), .B(N39), .S(n7168), .Z(cv_next_d[138]) );
  MUX2_X2 U7493 ( .A(cv_next[139]), .B(N40), .S(n7168), .Z(cv_next_d[139]) );
  MUX2_X2 U7494 ( .A(cv_next[140]), .B(N41), .S(n7168), .Z(cv_next_d[140]) );
  MUX2_X2 U7495 ( .A(cv_next[141]), .B(N42), .S(n7168), .Z(cv_next_d[141]) );
  MUX2_X2 U7496 ( .A(cv_next[142]), .B(N43), .S(n7168), .Z(cv_next_d[142]) );
  MUX2_X2 U7497 ( .A(cv_next[143]), .B(N44), .S(n7168), .Z(cv_next_d[143]) );
  MUX2_X2 U7498 ( .A(cv_next[144]), .B(N45), .S(n7168), .Z(cv_next_d[144]) );
  MUX2_X2 U7499 ( .A(cv_next[145]), .B(N46), .S(n7168), .Z(cv_next_d[145]) );
  MUX2_X2 U7500 ( .A(cv_next[146]), .B(N47), .S(n7168), .Z(cv_next_d[146]) );
  MUX2_X2 U7501 ( .A(cv_next[147]), .B(N48), .S(n7167), .Z(cv_next_d[147]) );
  MUX2_X2 U7502 ( .A(cv_next[148]), .B(N49), .S(n7167), .Z(cv_next_d[148]) );
  MUX2_X2 U7503 ( .A(cv_next[149]), .B(N50), .S(n7167), .Z(cv_next_d[149]) );
  MUX2_X2 U7504 ( .A(cv_next[150]), .B(N51), .S(n7167), .Z(cv_next_d[150]) );
  MUX2_X2 U7505 ( .A(cv_next[151]), .B(N52), .S(n7167), .Z(cv_next_d[151]) );
  MUX2_X2 U7506 ( .A(cv_next[152]), .B(N53), .S(n7167), .Z(cv_next_d[152]) );
  MUX2_X2 U7507 ( .A(cv_next[153]), .B(N54), .S(n7167), .Z(cv_next_d[153]) );
  MUX2_X2 U7508 ( .A(cv_next[154]), .B(N55), .S(n7167), .Z(cv_next_d[154]) );
  MUX2_X2 U7509 ( .A(cv_next[155]), .B(N56), .S(n7167), .Z(cv_next_d[155]) );
  MUX2_X2 U7510 ( .A(cv_next[156]), .B(N57), .S(n7167), .Z(cv_next_d[156]) );
  MUX2_X2 U7511 ( .A(cv_next[157]), .B(N58), .S(n7167), .Z(cv_next_d[157]) );
  MUX2_X2 U7512 ( .A(cv_next[158]), .B(N59), .S(n7167), .Z(cv_next_d[158]) );
  MUX2_X2 U7513 ( .A(cv_next[159]), .B(N60), .S(n7167), .Z(cv_next_d[159]) );
  INV_X4 U7514 ( .A(state[1]), .ZN(n7281) );
  NAND2_X2 U7515 ( .A1(state[0]), .A2(n7281), .ZN(n7395) );
  INV_X4 U7516 ( .A(use_prev_cv), .ZN(n7282) );
  NAND2_X2 U7517 ( .A1(n7395), .A2(n7282), .ZN(n7283) );
  NAND2_X2 U7518 ( .A1(use_prev_cv), .A2(n7395), .ZN(n7284) );
  NAND2_X2 U7519 ( .A1(cv_next[138]), .A2(n7137), .ZN(n7285) );
  NAND2_X2 U7520 ( .A1(sha1_round_wire[138]), .A2(n7152), .ZN(n7288) );
  NAND2_X2 U7521 ( .A1(n7394), .A2(n7288), .ZN(rnd_d[138]) );
  NAND2_X2 U7522 ( .A1(cv_next[139]), .A2(n7137), .ZN(n7289) );
  NAND2_X2 U7523 ( .A1(sha1_round_wire[139]), .A2(n7162), .ZN(n7292) );
  NAND2_X2 U7524 ( .A1(n7393), .A2(n7292), .ZN(rnd_d[139]) );
  NAND2_X2 U7525 ( .A1(cv_next[140]), .A2(n7137), .ZN(n7293) );
  NAND2_X2 U7526 ( .A1(sha1_round_wire[140]), .A2(n7158), .ZN(n7296) );
  NAND2_X2 U7527 ( .A1(n7392), .A2(n7296), .ZN(rnd_d[140]) );
  NAND2_X2 U7528 ( .A1(cv_next[141]), .A2(n7137), .ZN(n7297) );
  NAND2_X2 U7529 ( .A1(sha1_round_wire[141]), .A2(n7158), .ZN(n7300) );
  NAND2_X2 U7530 ( .A1(n7391), .A2(n7300), .ZN(rnd_d[141]) );
  NAND2_X2 U7531 ( .A1(cv_next[142]), .A2(n7137), .ZN(n7301) );
  NAND2_X2 U7532 ( .A1(sha1_round_wire[142]), .A2(n7158), .ZN(n7304) );
  NAND2_X2 U7533 ( .A1(n7390), .A2(n7304), .ZN(rnd_d[142]) );
  NAND2_X2 U7534 ( .A1(cv_next[143]), .A2(n7137), .ZN(n7305) );
  NAND2_X2 U7535 ( .A1(sha1_round_wire[143]), .A2(n7158), .ZN(n7308) );
  NAND2_X2 U7536 ( .A1(n7389), .A2(n7308), .ZN(rnd_d[143]) );
  NAND2_X2 U7537 ( .A1(cv_next[144]), .A2(n7137), .ZN(n7309) );
  NAND2_X2 U7538 ( .A1(sha1_round_wire[144]), .A2(n7158), .ZN(n7312) );
  NAND2_X2 U7539 ( .A1(n7388), .A2(n7312), .ZN(rnd_d[144]) );
  NAND2_X2 U7540 ( .A1(cv_next[145]), .A2(n7137), .ZN(n7313) );
  NAND2_X2 U7541 ( .A1(sha1_round_wire[145]), .A2(n7158), .ZN(n7316) );
  NAND2_X2 U7542 ( .A1(n7387), .A2(n7316), .ZN(rnd_d[145]) );
  NAND2_X2 U7543 ( .A1(cv_next[146]), .A2(n7137), .ZN(n7317) );
  NAND2_X2 U7544 ( .A1(sha1_round_wire[146]), .A2(n7159), .ZN(n7320) );
  NAND2_X2 U7545 ( .A1(n7386), .A2(n7320), .ZN(rnd_d[146]) );
  NAND2_X2 U7546 ( .A1(cv_next[147]), .A2(n7137), .ZN(n7321) );
  NAND2_X2 U7547 ( .A1(sha1_round_wire[147]), .A2(n7159), .ZN(n7324) );
  NAND2_X2 U7548 ( .A1(n7385), .A2(n7324), .ZN(rnd_d[147]) );
  NAND2_X2 U7549 ( .A1(cv_next[148]), .A2(n7137), .ZN(n7325) );
  NAND2_X2 U7550 ( .A1(sha1_round_wire[148]), .A2(n7159), .ZN(n7328) );
  NAND2_X2 U7551 ( .A1(n7384), .A2(n7328), .ZN(rnd_d[148]) );
  NAND2_X2 U7552 ( .A1(cv_next[149]), .A2(n7138), .ZN(n7329) );
  NAND2_X2 U7553 ( .A1(sha1_round_wire[149]), .A2(n7159), .ZN(n7332) );
  NAND2_X2 U7554 ( .A1(n7332), .A2(n7383), .ZN(rnd_d[149]) );
  NAND2_X2 U7555 ( .A1(cv_next[150]), .A2(n7138), .ZN(n7333) );
  NAND2_X2 U7556 ( .A1(sha1_round_wire[150]), .A2(n7159), .ZN(n7336) );
  NAND2_X2 U7557 ( .A1(n7382), .A2(n7336), .ZN(rnd_d[150]) );
  NAND2_X2 U7558 ( .A1(cv_next[151]), .A2(n7138), .ZN(n7337) );
  NAND2_X2 U7559 ( .A1(cv_next[152]), .A2(n7138), .ZN(n7341) );
  NAND2_X2 U7560 ( .A1(sha1_round_wire[152]), .A2(n7159), .ZN(n7344) );
  NAND2_X2 U7561 ( .A1(n7380), .A2(n7344), .ZN(rnd_d[152]) );
  NAND2_X2 U7562 ( .A1(cv_next[153]), .A2(n7138), .ZN(n7345) );
  NAND2_X2 U7563 ( .A1(sha1_round_wire[153]), .A2(n7159), .ZN(n7348) );
  NAND2_X2 U7564 ( .A1(n7348), .A2(n7379), .ZN(rnd_d[153]) );
  NAND2_X2 U7565 ( .A1(cv_next[154]), .A2(n7138), .ZN(n7349) );
  NAND2_X2 U7566 ( .A1(sha1_round_wire[154]), .A2(n7159), .ZN(n7352) );
  NAND2_X2 U7567 ( .A1(n7352), .A2(n7378), .ZN(rnd_d[154]) );
  NAND2_X2 U7568 ( .A1(cv_next[155]), .A2(n7138), .ZN(n7353) );
  NAND2_X2 U7569 ( .A1(sha1_round_wire[155]), .A2(n7159), .ZN(n7356) );
  NAND2_X2 U7570 ( .A1(cv_next[156]), .A2(n7138), .ZN(n7357) );
  NAND2_X2 U7571 ( .A1(sha1_round_wire[156]), .A2(n7159), .ZN(n7360) );
  NAND2_X2 U7572 ( .A1(n7376), .A2(n7360), .ZN(rnd_d[156]) );
  NAND2_X2 U7573 ( .A1(cv_next[157]), .A2(n7138), .ZN(n7361) );
  NAND2_X2 U7574 ( .A1(n7375), .A2(n7364), .ZN(rnd_d[157]) );
  NAND2_X2 U7575 ( .A1(cv_next[158]), .A2(n7138), .ZN(n7365) );
  NAND2_X2 U7576 ( .A1(sha1_round_wire[158]), .A2(n7159), .ZN(n7368) );
  NAND2_X2 U7577 ( .A1(n7368), .A2(n7374), .ZN(rnd_d[158]) );
  NAND2_X2 U7578 ( .A1(cv_next[159]), .A2(n7138), .ZN(n7369) );
  INV_X4 U7579 ( .A(n6230), .ZN(n7396) );
  INV_X4 U7580 ( .A(rnd_cnt_d[0]), .ZN(n7397) );
  INV_X4 U7581 ( .A(rnd_cnt_q[1]), .ZN(n7401) );
  INV_X4 U7582 ( .A(n7116), .ZN(n7402) );
  INV_X4 U7583 ( .A(load_in), .ZN(n7403) );
  NAND2_X2 \sha1_round/U575  ( .A1(\sha1_round/n3200 ), .A2(\sha1_round/n821 ), 
        .ZN(\sha1_round/k[13] ) );
  INV_X4 \sha1_round/U574  ( .A(\sha1_round/k_23 ), .ZN(\sha1_round/n821 ) );
  NAND2_X2 \sha1_round/U573  ( .A1(\sha1_round/n819 ), .A2(\sha1_round/n510 ), 
        .ZN(\sha1_round/k_23 ) );
  INV_X4 \sha1_round/U572  ( .A(\sha1_round/n2 ), .ZN(\sha1_round/n818 ) );
  NAND2_X2 \sha1_round/U571  ( .A1(rnd_q[32]), .A2(\sha1_round/n812 ), .ZN(
        \sha1_round/n813 ) );
  NAND2_X2 \sha1_round/U570  ( .A1(\sha1_round/n811 ), .A2(\sha1_round/n810 ), 
        .ZN(\sha1_round/n812 ) );
  NAND2_X2 \sha1_round/U569  ( .A1(\sha1_round/n808 ), .A2(\sha1_round/n807 ), 
        .ZN(\sha1_round/n809 ) );
  INV_X4 \sha1_round/U568  ( .A(rnd_q[64]), .ZN(\sha1_round/n807 ) );
  NAND2_X2 \sha1_round/U567  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n808 ), 
        .ZN(\sha1_round/n811 ) );
  INV_X4 \sha1_round/U566  ( .A(rnd_q[32]), .ZN(\sha1_round/n804 ) );
  INV_X4 \sha1_round/U565  ( .A(\sha1_round/n806 ), .ZN(\sha1_round/n805 ) );
  XOR2_X2 \sha1_round/U564  ( .A(\sha1_round/n808 ), .B(rnd_q[64]), .Z(
        \sha1_round/n806 ) );
  INV_X4 \sha1_round/U563  ( .A(rnd_q[96]), .ZN(\sha1_round/n808 ) );
  NAND2_X2 \sha1_round/U562  ( .A1(\sha1_round/n798 ), .A2(\sha1_round/n797 ), 
        .ZN(\sha1_round/n799 ) );
  NAND2_X2 \sha1_round/U561  ( .A1(\sha1_round/n795 ), .A2(\sha1_round/n794 ), 
        .ZN(\sha1_round/n796 ) );
  INV_X4 \sha1_round/U560  ( .A(rnd_q[65]), .ZN(\sha1_round/n794 ) );
  NAND2_X2 \sha1_round/U559  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n795 ), 
        .ZN(\sha1_round/n798 ) );
  INV_X4 \sha1_round/U558  ( .A(\sha1_round/n793 ), .ZN(\sha1_round/n792 ) );
  XOR2_X2 \sha1_round/U557  ( .A(\sha1_round/n795 ), .B(rnd_q[65]), .Z(
        \sha1_round/n793 ) );
  INV_X4 \sha1_round/U556  ( .A(rnd_q[97]), .ZN(\sha1_round/n795 ) );
  NAND2_X2 \sha1_round/U555  ( .A1(rnd_q[34]), .A2(\sha1_round/n786 ), .ZN(
        \sha1_round/n787 ) );
  NAND2_X2 \sha1_round/U554  ( .A1(\sha1_round/n785 ), .A2(\sha1_round/n784 ), 
        .ZN(\sha1_round/n786 ) );
  NAND2_X2 \sha1_round/U553  ( .A1(\sha1_round/n782 ), .A2(\sha1_round/n781 ), 
        .ZN(\sha1_round/n783 ) );
  INV_X4 \sha1_round/U552  ( .A(rnd_q[66]), .ZN(\sha1_round/n781 ) );
  NAND2_X2 \sha1_round/U551  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n782 ), 
        .ZN(\sha1_round/n785 ) );
  INV_X4 \sha1_round/U550  ( .A(rnd_q[34]), .ZN(\sha1_round/n778 ) );
  INV_X4 \sha1_round/U549  ( .A(\sha1_round/n780 ), .ZN(\sha1_round/n779 ) );
  XOR2_X2 \sha1_round/U548  ( .A(\sha1_round/n782 ), .B(rnd_q[66]), .Z(
        \sha1_round/n780 ) );
  INV_X4 \sha1_round/U547  ( .A(rnd_q[98]), .ZN(\sha1_round/n782 ) );
  NAND2_X2 \sha1_round/U546  ( .A1(\sha1_round/n772 ), .A2(\sha1_round/n771 ), 
        .ZN(\sha1_round/n773 ) );
  NAND2_X2 \sha1_round/U545  ( .A1(\sha1_round/n769 ), .A2(\sha1_round/n768 ), 
        .ZN(\sha1_round/n770 ) );
  INV_X4 \sha1_round/U544  ( .A(rnd_q[67]), .ZN(\sha1_round/n768 ) );
  NAND2_X2 \sha1_round/U543  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n769 ), 
        .ZN(\sha1_round/n772 ) );
  INV_X4 \sha1_round/U542  ( .A(rnd_q[35]), .ZN(\sha1_round/n764 ) );
  INV_X4 \sha1_round/U541  ( .A(\sha1_round/n766 ), .ZN(\sha1_round/n765 ) );
  XOR2_X2 \sha1_round/U540  ( .A(\sha1_round/n769 ), .B(rnd_q[67]), .Z(
        \sha1_round/n766 ) );
  INV_X4 \sha1_round/U539  ( .A(rnd_q[99]), .ZN(\sha1_round/n769 ) );
  MUX2_X2 \sha1_round/U538  ( .A(\sha1_round/n761 ), .B(\sha1_round/n760 ), 
        .S(rnd_q[36]), .Z(\sha1_round/n762 ) );
  NOR3_X2 \sha1_round/U537  ( .A1(\sha1_round/n759 ), .A2(\sha1_round/n758 ), 
        .A3(\sha1_round/n757 ), .ZN(\sha1_round/n760 ) );
  NOR2_X2 \sha1_round/U536  ( .A1(\sha1_round/n755 ), .A2(\sha1_round/n3180 ), 
        .ZN(\sha1_round/n758 ) );
  NOR2_X2 \sha1_round/U535  ( .A1(rnd_q[68]), .A2(rnd_q[100]), .ZN(
        \sha1_round/n755 ) );
  NOR2_X2 \sha1_round/U534  ( .A1(rnd_q[100]), .A2(\sha1_round/n510 ), .ZN(
        \sha1_round/n759 ) );
  NAND2_X2 \sha1_round/U533  ( .A1(\sha1_round/n374 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n761 ) );
  NAND3_X2 \sha1_round/U532  ( .A1(rnd_q[68]), .A2(rnd_q[100]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n763 ) );
  NOR2_X2 \sha1_round/U531  ( .A1(rnd_q[69]), .A2(rnd_q[101]), .ZN(
        \sha1_round/n750 ) );
  NAND3_X2 \sha1_round/U530  ( .A1(rnd_q[69]), .A2(rnd_q[101]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n754 ) );
  NOR2_X2 \sha1_round/U529  ( .A1(rnd_q[70]), .A2(rnd_q[102]), .ZN(
        \sha1_round/n745 ) );
  NAND3_X2 \sha1_round/U528  ( .A1(rnd_q[70]), .A2(rnd_q[102]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n749 ) );
  NOR3_X2 \sha1_round/U527  ( .A1(\sha1_round/n740 ), .A2(\sha1_round/n739 ), 
        .A3(\sha1_round/n738 ), .ZN(\sha1_round/n741 ) );
  NOR2_X2 \sha1_round/U526  ( .A1(\sha1_round/n737 ), .A2(\sha1_round/n514 ), 
        .ZN(\sha1_round/n739 ) );
  NOR2_X2 \sha1_round/U525  ( .A1(rnd_q[71]), .A2(rnd_q[103]), .ZN(
        \sha1_round/n737 ) );
  NOR2_X2 \sha1_round/U524  ( .A1(rnd_q[103]), .A2(\sha1_round/n510 ), .ZN(
        \sha1_round/n740 ) );
  NAND3_X2 \sha1_round/U523  ( .A1(rnd_q[71]), .A2(rnd_q[103]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n744 ) );
  NOR2_X2 \sha1_round/U522  ( .A1(\sha1_round/n729 ), .A2(\sha1_round/n514 ), 
        .ZN(\sha1_round/n731 ) );
  NOR2_X2 \sha1_round/U521  ( .A1(rnd_q[72]), .A2(rnd_q[104]), .ZN(
        \sha1_round/n729 ) );
  NAND3_X2 \sha1_round/U520  ( .A1(rnd_q[72]), .A2(rnd_q[104]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n736 ) );
  NAND3_X2 \sha1_round/U519  ( .A1(rnd_q[73]), .A2(rnd_q[105]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n728 ) );
  NOR2_X2 \sha1_round/U518  ( .A1(\sha1_round/n714 ), .A2(\sha1_round/n3180 ), 
        .ZN(\sha1_round/n716 ) );
  NOR2_X2 \sha1_round/U517  ( .A1(rnd_q[74]), .A2(rnd_q[106]), .ZN(
        \sha1_round/n714 ) );
  NOR2_X2 \sha1_round/U516  ( .A1(rnd_q[106]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n717 ) );
  NAND3_X2 \sha1_round/U515  ( .A1(rnd_q[74]), .A2(rnd_q[106]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n721 ) );
  NOR2_X2 \sha1_round/U514  ( .A1(rnd_q[75]), .A2(rnd_q[107]), .ZN(
        \sha1_round/n706 ) );
  NAND3_X2 \sha1_round/U513  ( .A1(rnd_q[75]), .A2(rnd_q[107]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n713 ) );
  MUX2_X2 \sha1_round/U512  ( .A(\sha1_round/n703 ), .B(\sha1_round/n702 ), 
        .S(rnd_q[44]), .Z(\sha1_round/n704 ) );
  NOR3_X2 \sha1_round/U511  ( .A1(\sha1_round/n701 ), .A2(\sha1_round/n700 ), 
        .A3(\sha1_round/n699 ), .ZN(\sha1_round/n702 ) );
  NOR2_X2 \sha1_round/U510  ( .A1(\sha1_round/n698 ), .A2(\sha1_round/n3190 ), 
        .ZN(\sha1_round/n700 ) );
  NOR2_X2 \sha1_round/U509  ( .A1(rnd_q[76]), .A2(rnd_q[108]), .ZN(
        \sha1_round/n698 ) );
  NAND3_X2 \sha1_round/U508  ( .A1(rnd_q[76]), .A2(rnd_q[108]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n705 ) );
  MUX2_X2 \sha1_round/U507  ( .A(\sha1_round/n695 ), .B(\sha1_round/n694 ), 
        .S(rnd_q[45]), .Z(\sha1_round/n696 ) );
  NOR3_X2 \sha1_round/U506  ( .A1(\sha1_round/n693 ), .A2(\sha1_round/n692 ), 
        .A3(\sha1_round/n691 ), .ZN(\sha1_round/n694 ) );
  NOR2_X2 \sha1_round/U505  ( .A1(\sha1_round/n690 ), .A2(\sha1_round/n3160 ), 
        .ZN(\sha1_round/n692 ) );
  NOR2_X2 \sha1_round/U504  ( .A1(rnd_q[77]), .A2(rnd_q[109]), .ZN(
        \sha1_round/n690 ) );
  NAND3_X2 \sha1_round/U503  ( .A1(rnd_q[77]), .A2(rnd_q[109]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n697 ) );
  MUX2_X2 \sha1_round/U502  ( .A(\sha1_round/n687 ), .B(\sha1_round/n686 ), 
        .S(rnd_q[46]), .Z(\sha1_round/n688 ) );
  NOR3_X2 \sha1_round/U501  ( .A1(\sha1_round/n685 ), .A2(\sha1_round/n684 ), 
        .A3(\sha1_round/n683 ), .ZN(\sha1_round/n686 ) );
  NOR2_X2 \sha1_round/U500  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n368 ), 
        .ZN(\sha1_round/n683 ) );
  NOR2_X2 \sha1_round/U499  ( .A1(\sha1_round/n682 ), .A2(\sha1_round/n3160 ), 
        .ZN(\sha1_round/n684 ) );
  NOR2_X2 \sha1_round/U498  ( .A1(rnd_q[78]), .A2(rnd_q[110]), .ZN(
        \sha1_round/n682 ) );
  NAND3_X2 \sha1_round/U497  ( .A1(rnd_q[78]), .A2(rnd_q[110]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n689 ) );
  NAND2_X2 \sha1_round/U496  ( .A1(\sha1_round/n681 ), .A2(\sha1_round/n680 ), 
        .ZN(\sha1_round/f [15]) );
  MUX2_X2 \sha1_round/U495  ( .A(\sha1_round/n679 ), .B(\sha1_round/n678 ), 
        .S(rnd_q[47]), .Z(\sha1_round/n680 ) );
  NOR3_X2 \sha1_round/U494  ( .A1(\sha1_round/n677 ), .A2(\sha1_round/n676 ), 
        .A3(\sha1_round/n675 ), .ZN(\sha1_round/n678 ) );
  NOR2_X2 \sha1_round/U493  ( .A1(\sha1_round/n674 ), .A2(\sha1_round/n3120 ), 
        .ZN(\sha1_round/n676 ) );
  NOR2_X2 \sha1_round/U492  ( .A1(rnd_q[79]), .A2(rnd_q[111]), .ZN(
        \sha1_round/n674 ) );
  NAND3_X2 \sha1_round/U491  ( .A1(rnd_q[79]), .A2(rnd_q[111]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n681 ) );
  NAND2_X2 \sha1_round/U490  ( .A1(\sha1_round/n673 ), .A2(\sha1_round/n672 ), 
        .ZN(\sha1_round/f [16]) );
  MUX2_X2 \sha1_round/U489  ( .A(\sha1_round/n671 ), .B(\sha1_round/n670 ), 
        .S(rnd_q[48]), .Z(\sha1_round/n672 ) );
  NOR3_X2 \sha1_round/U488  ( .A1(\sha1_round/n669 ), .A2(\sha1_round/n668 ), 
        .A3(\sha1_round/n667 ), .ZN(\sha1_round/n670 ) );
  NOR2_X2 \sha1_round/U487  ( .A1(\sha1_round/n666 ), .A2(\sha1_round/n3160 ), 
        .ZN(\sha1_round/n668 ) );
  NOR2_X2 \sha1_round/U486  ( .A1(rnd_q[80]), .A2(rnd_q[112]), .ZN(
        \sha1_round/n666 ) );
  NAND3_X2 \sha1_round/U485  ( .A1(rnd_q[80]), .A2(rnd_q[112]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n673 ) );
  NAND2_X2 \sha1_round/U484  ( .A1(\sha1_round/n665 ), .A2(\sha1_round/n664 ), 
        .ZN(\sha1_round/f [17]) );
  MUX2_X2 \sha1_round/U483  ( .A(\sha1_round/n663 ), .B(\sha1_round/n662 ), 
        .S(rnd_q[49]), .Z(\sha1_round/n664 ) );
  NOR3_X2 \sha1_round/U482  ( .A1(\sha1_round/n661 ), .A2(\sha1_round/n660 ), 
        .A3(\sha1_round/n659 ), .ZN(\sha1_round/n662 ) );
  NOR2_X2 \sha1_round/U481  ( .A1(\sha1_round/n658 ), .A2(\sha1_round/n3200 ), 
        .ZN(\sha1_round/n660 ) );
  NOR2_X2 \sha1_round/U480  ( .A1(rnd_q[81]), .A2(rnd_q[113]), .ZN(
        \sha1_round/n658 ) );
  NAND3_X2 \sha1_round/U479  ( .A1(rnd_q[81]), .A2(rnd_q[113]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n665 ) );
  NAND2_X2 \sha1_round/U478  ( .A1(\sha1_round/n657 ), .A2(\sha1_round/n656 ), 
        .ZN(\sha1_round/f [18]) );
  MUX2_X2 \sha1_round/U477  ( .A(\sha1_round/n655 ), .B(\sha1_round/n654 ), 
        .S(rnd_q[50]), .Z(\sha1_round/n656 ) );
  NOR3_X2 \sha1_round/U476  ( .A1(\sha1_round/n653 ), .A2(\sha1_round/n652 ), 
        .A3(\sha1_round/n651 ), .ZN(\sha1_round/n654 ) );
  NOR2_X2 \sha1_round/U475  ( .A1(\sha1_round/n650 ), .A2(\sha1_round/n513 ), 
        .ZN(\sha1_round/n652 ) );
  NOR2_X2 \sha1_round/U474  ( .A1(rnd_q[82]), .A2(rnd_q[114]), .ZN(
        \sha1_round/n650 ) );
  NAND3_X2 \sha1_round/U473  ( .A1(rnd_q[82]), .A2(rnd_q[114]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n657 ) );
  NAND2_X2 \sha1_round/U472  ( .A1(\sha1_round/n649 ), .A2(\sha1_round/n648 ), 
        .ZN(\sha1_round/f [19]) );
  MUX2_X2 \sha1_round/U471  ( .A(\sha1_round/n647 ), .B(\sha1_round/n646 ), 
        .S(rnd_q[51]), .Z(\sha1_round/n648 ) );
  NOR3_X2 \sha1_round/U470  ( .A1(\sha1_round/n645 ), .A2(\sha1_round/n644 ), 
        .A3(\sha1_round/n643 ), .ZN(\sha1_round/n646 ) );
  NOR2_X2 \sha1_round/U469  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n371 ), 
        .ZN(\sha1_round/n643 ) );
  NOR2_X2 \sha1_round/U468  ( .A1(\sha1_round/n642 ), .A2(\sha1_round/n3180 ), 
        .ZN(\sha1_round/n644 ) );
  NOR2_X2 \sha1_round/U467  ( .A1(rnd_q[83]), .A2(rnd_q[115]), .ZN(
        \sha1_round/n642 ) );
  NAND3_X2 \sha1_round/U466  ( .A1(rnd_q[83]), .A2(rnd_q[115]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n649 ) );
  MUX2_X2 \sha1_round/U465  ( .A(\sha1_round/n639 ), .B(\sha1_round/n638 ), 
        .S(rnd_q[52]), .Z(\sha1_round/n640 ) );
  NOR3_X2 \sha1_round/U464  ( .A1(\sha1_round/n637 ), .A2(\sha1_round/n636 ), 
        .A3(\sha1_round/n635 ), .ZN(\sha1_round/n638 ) );
  NOR2_X2 \sha1_round/U463  ( .A1(\sha1_round/n634 ), .A2(\sha1_round/n3180 ), 
        .ZN(\sha1_round/n636 ) );
  NOR2_X2 \sha1_round/U462  ( .A1(rnd_q[84]), .A2(rnd_q[116]), .ZN(
        \sha1_round/n634 ) );
  NAND3_X2 \sha1_round/U461  ( .A1(rnd_q[84]), .A2(rnd_q[116]), .A3(
        \sha1_round/n517 ), .ZN(\sha1_round/n641 ) );
  NAND2_X2 \sha1_round/U460  ( .A1(\sha1_round/n633 ), .A2(\sha1_round/n632 ), 
        .ZN(\sha1_round/f [21]) );
  MUX2_X2 \sha1_round/U459  ( .A(\sha1_round/n631 ), .B(\sha1_round/n630 ), 
        .S(rnd_q[53]), .Z(\sha1_round/n632 ) );
  NOR3_X2 \sha1_round/U458  ( .A1(\sha1_round/n629 ), .A2(\sha1_round/n628 ), 
        .A3(\sha1_round/n627 ), .ZN(\sha1_round/n630 ) );
  NOR2_X2 \sha1_round/U457  ( .A1(\sha1_round/n626 ), .A2(\sha1_round/n514 ), 
        .ZN(\sha1_round/n628 ) );
  NOR2_X2 \sha1_round/U456  ( .A1(rnd_q[85]), .A2(rnd_q[117]), .ZN(
        \sha1_round/n626 ) );
  NAND3_X2 \sha1_round/U455  ( .A1(rnd_q[85]), .A2(rnd_q[117]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n633 ) );
  NAND2_X2 \sha1_round/U454  ( .A1(\sha1_round/n625 ), .A2(\sha1_round/n624 ), 
        .ZN(\sha1_round/f [22]) );
  MUX2_X2 \sha1_round/U453  ( .A(\sha1_round/n623 ), .B(\sha1_round/n622 ), 
        .S(rnd_q[54]), .Z(\sha1_round/n624 ) );
  NOR3_X2 \sha1_round/U452  ( .A1(\sha1_round/n621 ), .A2(\sha1_round/n620 ), 
        .A3(\sha1_round/n619 ), .ZN(\sha1_round/n622 ) );
  NOR2_X2 \sha1_round/U451  ( .A1(\sha1_round/n618 ), .A2(\sha1_round/n514 ), 
        .ZN(\sha1_round/n620 ) );
  NOR2_X2 \sha1_round/U450  ( .A1(rnd_q[86]), .A2(rnd_q[118]), .ZN(
        \sha1_round/n618 ) );
  NAND3_X2 \sha1_round/U449  ( .A1(rnd_q[86]), .A2(rnd_q[118]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n625 ) );
  NAND2_X2 \sha1_round/U448  ( .A1(\sha1_round/n617 ), .A2(\sha1_round/n616 ), 
        .ZN(\sha1_round/f [23]) );
  MUX2_X2 \sha1_round/U447  ( .A(\sha1_round/n615 ), .B(\sha1_round/n614 ), 
        .S(rnd_q[55]), .Z(\sha1_round/n616 ) );
  AND3_X2 \sha1_round/U446  ( .A1(\sha1_round/n613 ), .A2(\sha1_round/n612 ), 
        .A3(\sha1_round/n611 ), .ZN(\sha1_round/n614 ) );
  NAND2_X2 \sha1_round/U445  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n610 ), 
        .ZN(\sha1_round/n611 ) );
  INV_X4 \sha1_round/U444  ( .A(rnd_q[119]), .ZN(\sha1_round/n610 ) );
  NAND2_X2 \sha1_round/U443  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n609 ), 
        .ZN(\sha1_round/n615 ) );
  INV_X4 \sha1_round/U442  ( .A(\sha1_round/n168 ), .ZN(\sha1_round/n609 ) );
  NAND3_X2 \sha1_round/U441  ( .A1(rnd_q[87]), .A2(rnd_q[119]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n617 ) );
  NAND2_X2 \sha1_round/U440  ( .A1(\sha1_round/n608 ), .A2(\sha1_round/n607 ), 
        .ZN(\sha1_round/f [24]) );
  MUX2_X2 \sha1_round/U439  ( .A(\sha1_round/n606 ), .B(\sha1_round/n605 ), 
        .S(rnd_q[56]), .Z(\sha1_round/n607 ) );
  AND3_X2 \sha1_round/U438  ( .A1(\sha1_round/n604 ), .A2(\sha1_round/n603 ), 
        .A3(\sha1_round/n602 ), .ZN(\sha1_round/n605 ) );
  NAND2_X2 \sha1_round/U437  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n601 ), 
        .ZN(\sha1_round/n602 ) );
  INV_X4 \sha1_round/U436  ( .A(rnd_q[120]), .ZN(\sha1_round/n601 ) );
  NAND2_X2 \sha1_round/U435  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n600 ), 
        .ZN(\sha1_round/n606 ) );
  INV_X4 \sha1_round/U434  ( .A(\sha1_round/n159 ), .ZN(\sha1_round/n600 ) );
  NAND3_X2 \sha1_round/U433  ( .A1(rnd_q[88]), .A2(rnd_q[120]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n608 ) );
  NAND2_X2 \sha1_round/U432  ( .A1(\sha1_round/n599 ), .A2(\sha1_round/n598 ), 
        .ZN(\sha1_round/f [25]) );
  MUX2_X2 \sha1_round/U431  ( .A(\sha1_round/n597 ), .B(\sha1_round/n596 ), 
        .S(rnd_q[57]), .Z(\sha1_round/n598 ) );
  AND3_X2 \sha1_round/U430  ( .A1(\sha1_round/n595 ), .A2(\sha1_round/n594 ), 
        .A3(\sha1_round/n593 ), .ZN(\sha1_round/n596 ) );
  NAND2_X2 \sha1_round/U429  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n592 ), 
        .ZN(\sha1_round/n593 ) );
  INV_X4 \sha1_round/U428  ( .A(rnd_q[121]), .ZN(\sha1_round/n592 ) );
  NAND2_X2 \sha1_round/U427  ( .A1(\sha1_round/n150 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n594 ) );
  NAND2_X2 \sha1_round/U426  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n591 ), 
        .ZN(\sha1_round/n597 ) );
  INV_X4 \sha1_round/U425  ( .A(\sha1_round/n150 ), .ZN(\sha1_round/n591 ) );
  NAND3_X2 \sha1_round/U424  ( .A1(rnd_q[89]), .A2(rnd_q[121]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n599 ) );
  NAND2_X2 \sha1_round/U423  ( .A1(\sha1_round/n590 ), .A2(\sha1_round/n589 ), 
        .ZN(\sha1_round/f [26]) );
  MUX2_X2 \sha1_round/U422  ( .A(\sha1_round/n588 ), .B(\sha1_round/n587 ), 
        .S(rnd_q[58]), .Z(\sha1_round/n589 ) );
  AND3_X2 \sha1_round/U421  ( .A1(\sha1_round/n586 ), .A2(\sha1_round/n585 ), 
        .A3(\sha1_round/n584 ), .ZN(\sha1_round/n587 ) );
  NAND2_X2 \sha1_round/U420  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n583 ), 
        .ZN(\sha1_round/n584 ) );
  INV_X4 \sha1_round/U419  ( .A(rnd_q[122]), .ZN(\sha1_round/n583 ) );
  NAND2_X2 \sha1_round/U418  ( .A1(\sha1_round/n141 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n585 ) );
  NAND2_X2 \sha1_round/U417  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n582 ), 
        .ZN(\sha1_round/n588 ) );
  INV_X4 \sha1_round/U416  ( .A(\sha1_round/n141 ), .ZN(\sha1_round/n582 ) );
  NAND3_X2 \sha1_round/U415  ( .A1(rnd_q[90]), .A2(rnd_q[122]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n590 ) );
  NAND2_X2 \sha1_round/U414  ( .A1(\sha1_round/n581 ), .A2(\sha1_round/n580 ), 
        .ZN(\sha1_round/f [27]) );
  MUX2_X2 \sha1_round/U413  ( .A(\sha1_round/n579 ), .B(\sha1_round/n578 ), 
        .S(rnd_q[59]), .Z(\sha1_round/n580 ) );
  AND3_X2 \sha1_round/U412  ( .A1(\sha1_round/n577 ), .A2(\sha1_round/n576 ), 
        .A3(\sha1_round/n575 ), .ZN(\sha1_round/n578 ) );
  NAND2_X2 \sha1_round/U411  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n574 ), 
        .ZN(\sha1_round/n575 ) );
  INV_X4 \sha1_round/U410  ( .A(rnd_q[123]), .ZN(\sha1_round/n574 ) );
  NAND2_X2 \sha1_round/U409  ( .A1(\sha1_round/n132 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n576 ) );
  NAND2_X2 \sha1_round/U408  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n573 ), 
        .ZN(\sha1_round/n579 ) );
  INV_X4 \sha1_round/U407  ( .A(\sha1_round/n132 ), .ZN(\sha1_round/n573 ) );
  NAND3_X2 \sha1_round/U406  ( .A1(rnd_q[91]), .A2(rnd_q[123]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n581 ) );
  NAND2_X2 \sha1_round/U405  ( .A1(\sha1_round/n572 ), .A2(\sha1_round/n571 ), 
        .ZN(\sha1_round/f [28]) );
  MUX2_X2 \sha1_round/U404  ( .A(\sha1_round/n570 ), .B(\sha1_round/n569 ), 
        .S(rnd_q[60]), .Z(\sha1_round/n571 ) );
  AND3_X2 \sha1_round/U403  ( .A1(\sha1_round/n568 ), .A2(\sha1_round/n567 ), 
        .A3(\sha1_round/n566 ), .ZN(\sha1_round/n569 ) );
  NAND2_X2 \sha1_round/U402  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n565 ), 
        .ZN(\sha1_round/n566 ) );
  INV_X4 \sha1_round/U401  ( .A(rnd_q[124]), .ZN(\sha1_round/n565 ) );
  NAND2_X2 \sha1_round/U400  ( .A1(\sha1_round/n123 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n567 ) );
  NAND2_X2 \sha1_round/U399  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n564 ), 
        .ZN(\sha1_round/n570 ) );
  INV_X4 \sha1_round/U398  ( .A(\sha1_round/n123 ), .ZN(\sha1_round/n564 ) );
  NAND3_X2 \sha1_round/U397  ( .A1(rnd_q[92]), .A2(rnd_q[124]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n572 ) );
  NAND2_X2 \sha1_round/U396  ( .A1(\sha1_round/n563 ), .A2(\sha1_round/n562 ), 
        .ZN(\sha1_round/f [29]) );
  MUX2_X2 \sha1_round/U395  ( .A(\sha1_round/n561 ), .B(\sha1_round/n560 ), 
        .S(rnd_q[61]), .Z(\sha1_round/n562 ) );
  AND3_X2 \sha1_round/U394  ( .A1(\sha1_round/n559 ), .A2(\sha1_round/n558 ), 
        .A3(\sha1_round/n557 ), .ZN(\sha1_round/n560 ) );
  NAND2_X2 \sha1_round/U393  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n556 ), 
        .ZN(\sha1_round/n557 ) );
  INV_X4 \sha1_round/U392  ( .A(rnd_q[125]), .ZN(\sha1_round/n556 ) );
  NAND2_X2 \sha1_round/U391  ( .A1(\sha1_round/n114 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n558 ) );
  NAND2_X2 \sha1_round/U390  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n555 ), 
        .ZN(\sha1_round/n561 ) );
  INV_X4 \sha1_round/U389  ( .A(\sha1_round/n114 ), .ZN(\sha1_round/n555 ) );
  NAND3_X2 \sha1_round/U388  ( .A1(rnd_q[93]), .A2(rnd_q[125]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n563 ) );
  NAND2_X2 \sha1_round/U387  ( .A1(\sha1_round/n554 ), .A2(\sha1_round/n553 ), 
        .ZN(\sha1_round/f [30]) );
  MUX2_X2 \sha1_round/U386  ( .A(\sha1_round/n552 ), .B(\sha1_round/n551 ), 
        .S(rnd_q[62]), .Z(\sha1_round/n553 ) );
  AND3_X2 \sha1_round/U385  ( .A1(\sha1_round/n550 ), .A2(\sha1_round/n549 ), 
        .A3(\sha1_round/n548 ), .ZN(\sha1_round/n551 ) );
  NAND2_X2 \sha1_round/U384  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n547 ), 
        .ZN(\sha1_round/n548 ) );
  INV_X4 \sha1_round/U383  ( .A(rnd_q[126]), .ZN(\sha1_round/n547 ) );
  NAND2_X2 \sha1_round/U382  ( .A1(\sha1_round/n96 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n549 ) );
  NAND2_X2 \sha1_round/U381  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n546 ), 
        .ZN(\sha1_round/n552 ) );
  INV_X4 \sha1_round/U380  ( .A(\sha1_round/n96 ), .ZN(\sha1_round/n546 ) );
  NAND3_X2 \sha1_round/U379  ( .A1(rnd_q[94]), .A2(rnd_q[126]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n554 ) );
  NAND2_X2 \sha1_round/U378  ( .A1(\sha1_round/n545 ), .A2(\sha1_round/n544 ), 
        .ZN(\sha1_round/f [31]) );
  MUX2_X2 \sha1_round/U377  ( .A(\sha1_round/n543 ), .B(\sha1_round/n542 ), 
        .S(rnd_q[63]), .Z(\sha1_round/n544 ) );
  AND3_X2 \sha1_round/U376  ( .A1(\sha1_round/n541 ), .A2(\sha1_round/n540 ), 
        .A3(\sha1_round/n539 ), .ZN(\sha1_round/n542 ) );
  NAND2_X2 \sha1_round/U375  ( .A1(\sha1_round/n511 ), .A2(\sha1_round/n538 ), 
        .ZN(\sha1_round/n539 ) );
  INV_X4 \sha1_round/U374  ( .A(rnd_q[127]), .ZN(\sha1_round/n538 ) );
  NAND2_X2 \sha1_round/U373  ( .A1(\sha1_round/n87 ), .A2(\sha1_round/n3370 ), 
        .ZN(\sha1_round/n540 ) );
  NAND2_X2 \sha1_round/U372  ( .A1(\sha1_round/n3370 ), .A2(\sha1_round/n537 ), 
        .ZN(\sha1_round/n543 ) );
  INV_X4 \sha1_round/U371  ( .A(\sha1_round/n87 ), .ZN(\sha1_round/n537 ) );
  NAND3_X2 \sha1_round/U370  ( .A1(rnd_q[95]), .A2(rnd_q[127]), .A3(
        \sha1_round/n3300 ), .ZN(\sha1_round/n545 ) );
  NAND2_X2 \sha1_round/U369  ( .A1(\sha1_round/n533 ), .A2(\sha1_round/n534 ), 
        .ZN(\sha1_round/n536 ) );
  INV_X4 \sha1_round/U368  ( .A(\sha1_round/n520 ), .ZN(\sha1_round/n532 ) );
  INV_X32 \sha1_round/U367  ( .A(\sha1_round/n516 ), .ZN(\sha1_round/n515 ) );
  NAND2_X4 \sha1_round/U366  ( .A1(\sha1_round/n510 ), .A2(\sha1_round/n3120 ), 
        .ZN(\sha1_round/k[3] ) );
  NAND2_X4 \sha1_round/U365  ( .A1(\sha1_round/n530 ), .A2(\sha1_round/n529 ), 
        .ZN(\sha1_round/n819 ) );
  NAND2_X4 \sha1_round/U364  ( .A1(\sha1_round/n819 ), .A2(\sha1_round/n820 ), 
        .ZN(\sha1_round/n823 ) );
  NAND2_X4 \sha1_round/U363  ( .A1(\sha1_round/n748 ), .A2(\sha1_round/n749 ), 
        .ZN(\sha1_round/f [6]) );
  NAND2_X1 \sha1_round/U362  ( .A1(rnd_cnt_q[6]), .A2(\sha1_round/n531 ), .ZN(
        \sha1_round/n534 ) );
  NAND2_X4 \sha1_round/U361  ( .A1(\sha1_round/n536 ), .A2(\sha1_round/n535 ), 
        .ZN(\sha1_round/n820 ) );
  NAND3_X1 \sha1_round/U360  ( .A1(rnd_q[35]), .A2(\sha1_round/n767 ), .A3(
        \sha1_round/n766 ), .ZN(\sha1_round/n775 ) );
  INV_X16 \sha1_round/U359  ( .A(\sha1_round/n823 ), .ZN(\sha1_round/n516 ) );
  NAND2_X1 \sha1_round/U358  ( .A1(\sha1_round/n819 ), .A2(\sha1_round/n514 ), 
        .ZN(\sha1_round/k_26 ) );
  NAND2_X2 \sha1_round/U357  ( .A1(\sha1_round/n818 ), .A2(\sha1_round/n819 ), 
        .ZN(\sha1_round/k_27 ) );
  NAND2_X4 \sha1_round/U356  ( .A1(\sha1_round/n727 ), .A2(\sha1_round/n728 ), 
        .ZN(\sha1_round/f [9]) );
  INV_X1 \sha1_round/U355  ( .A(\sha1_round/n820 ), .ZN(\sha1_round/n824 ) );
  INV_X4 \sha1_round/U354  ( .A(\sha1_round/N332 ), .ZN(\sha1_round/n508 ) );
  NOR2_X1 \sha1_round/U353  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n378 ), 
        .ZN(\sha1_round/n699 ) );
  NOR2_X1 \sha1_round/U352  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n376 ), 
        .ZN(\sha1_round/n659 ) );
  NOR2_X1 \sha1_round/U351  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n380 ), 
        .ZN(\sha1_round/n619 ) );
  NAND2_X1 \sha1_round/U350  ( .A1(\sha1_round/n510 ), .A2(\sha1_round/n516 ), 
        .ZN(\sha1_round/k_30 ) );
  NAND2_X1 \sha1_round/U349  ( .A1(\sha1_round/n363 ), .A2(\sha1_round/n516 ), 
        .ZN(\sha1_round/k[15] ) );
  NAND3_X1 \sha1_round/U348  ( .A1(\sha1_round/n765 ), .A2(\sha1_round/n764 ), 
        .A3(\sha1_round/n767 ), .ZN(\sha1_round/n777 ) );
  NAND2_X1 \sha1_round/U347  ( .A1(\sha1_round/n3150 ), .A2(\sha1_round/n783 ), 
        .ZN(\sha1_round/n784 ) );
  NAND2_X1 \sha1_round/U346  ( .A1(\sha1_round/n3150 ), .A2(\sha1_round/n809 ), 
        .ZN(\sha1_round/n810 ) );
  NAND2_X1 \sha1_round/U345  ( .A1(\sha1_round/n167 ), .A2(\sha1_round/n360 ), 
        .ZN(\sha1_round/n613 ) );
  NAND2_X1 \sha1_round/U344  ( .A1(\sha1_round/n149 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n595 ) );
  NAND2_X1 \sha1_round/U343  ( .A1(\sha1_round/n158 ), .A2(\sha1_round/n360 ), 
        .ZN(\sha1_round/n604 ) );
  NAND2_X1 \sha1_round/U342  ( .A1(\sha1_round/n140 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n586 ) );
  NAND2_X1 \sha1_round/U341  ( .A1(\sha1_round/n131 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n577 ) );
  NAND2_X1 \sha1_round/U340  ( .A1(\sha1_round/n122 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n568 ) );
  NAND2_X1 \sha1_round/U339  ( .A1(\sha1_round/n113 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n559 ) );
  NAND2_X1 \sha1_round/U338  ( .A1(\sha1_round/n95 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n550 ) );
  NAND2_X1 \sha1_round/U337  ( .A1(\sha1_round/n86 ), .A2(\sha1_round/n364 ), 
        .ZN(\sha1_round/n541 ) );
  BUF_X4 \sha1_round/U336  ( .A(rnd_q[137]), .Z(sha1_round_wire[105]) );
  BUF_X4 \sha1_round/U335  ( .A(rnd_q[138]), .Z(sha1_round_wire[106]) );
  BUF_X4 \sha1_round/U334  ( .A(rnd_q[139]), .Z(sha1_round_wire[107]) );
  BUF_X4 \sha1_round/U333  ( .A(rnd_q[140]), .Z(sha1_round_wire[108]) );
  BUF_X4 \sha1_round/U332  ( .A(rnd_q[141]), .Z(sha1_round_wire[109]) );
  BUF_X4 \sha1_round/U331  ( .A(rnd_q[142]), .Z(sha1_round_wire[110]) );
  BUF_X4 \sha1_round/U330  ( .A(rnd_q[143]), .Z(sha1_round_wire[111]) );
  BUF_X4 \sha1_round/U329  ( .A(rnd_q[144]), .Z(sha1_round_wire[112]) );
  BUF_X4 \sha1_round/U328  ( .A(rnd_q[145]), .Z(sha1_round_wire[113]) );
  BUF_X4 \sha1_round/U327  ( .A(rnd_q[146]), .Z(sha1_round_wire[114]) );
  BUF_X4 \sha1_round/U326  ( .A(rnd_q[147]), .Z(sha1_round_wire[115]) );
  BUF_X4 \sha1_round/U325  ( .A(rnd_q[148]), .Z(sha1_round_wire[116]) );
  BUF_X4 \sha1_round/U324  ( .A(rnd_q[149]), .Z(sha1_round_wire[117]) );
  BUF_X4 \sha1_round/U323  ( .A(rnd_q[150]), .Z(sha1_round_wire[118]) );
  BUF_X4 \sha1_round/U322  ( .A(rnd_q[151]), .Z(sha1_round_wire[119]) );
  BUF_X4 \sha1_round/U321  ( .A(rnd_q[152]), .Z(sha1_round_wire[120]) );
  BUF_X4 \sha1_round/U320  ( .A(rnd_q[153]), .Z(sha1_round_wire[121]) );
  BUF_X4 \sha1_round/U319  ( .A(rnd_q[154]), .Z(sha1_round_wire[122]) );
  BUF_X4 \sha1_round/U318  ( .A(rnd_q[155]), .Z(sha1_round_wire[123]) );
  BUF_X4 \sha1_round/U317  ( .A(rnd_q[156]), .Z(sha1_round_wire[124]) );
  BUF_X4 \sha1_round/U316  ( .A(rnd_q[157]), .Z(sha1_round_wire[125]) );
  BUF_X4 \sha1_round/U315  ( .A(rnd_q[158]), .Z(sha1_round_wire[126]) );
  BUF_X4 \sha1_round/U314  ( .A(rnd_q[159]), .Z(sha1_round_wire[127]) );
  INV_X4 \sha1_round/U313  ( .A(rnd_cnt_q[3]), .ZN(\sha1_round/n524 ) );
  BUF_X4 \sha1_round/U312  ( .A(rnd_q[134]), .Z(sha1_round_wire[102]) );
  BUF_X4 \sha1_round/U311  ( .A(rnd_q[133]), .Z(sha1_round_wire[101]) );
  BUF_X4 \sha1_round/U310  ( .A(rnd_q[131]), .Z(sha1_round_wire[99]) );
  BUF_X4 \sha1_round/U309  ( .A(rnd_q[130]), .Z(sha1_round_wire[98]) );
  BUF_X4 \sha1_round/U308  ( .A(rnd_q[129]), .Z(sha1_round_wire[97]) );
  BUF_X4 \sha1_round/U307  ( .A(rnd_q[128]), .Z(sha1_round_wire[96]) );
  BUF_X4 \sha1_round/U306  ( .A(rnd_q[96]), .Z(sha1_round_wire[94]) );
  BUF_X4 \sha1_round/U305  ( .A(rnd_q[117]), .Z(sha1_round_wire[83]) );
  BUF_X4 \sha1_round/U304  ( .A(rnd_q[116]), .Z(sha1_round_wire[82]) );
  BUF_X4 \sha1_round/U303  ( .A(rnd_q[113]), .Z(sha1_round_wire[79]) );
  BUF_X4 \sha1_round/U302  ( .A(rnd_q[112]), .Z(sha1_round_wire[78]) );
  BUF_X4 \sha1_round/U301  ( .A(rnd_q[110]), .Z(sha1_round_wire[76]) );
  BUF_X4 \sha1_round/U300  ( .A(rnd_q[109]), .Z(sha1_round_wire[75]) );
  BUF_X4 \sha1_round/U299  ( .A(rnd_q[106]), .Z(sha1_round_wire[72]) );
  BUF_X4 \sha1_round/U298  ( .A(rnd_q[105]), .Z(sha1_round_wire[71]) );
  BUF_X4 \sha1_round/U297  ( .A(rnd_q[104]), .Z(sha1_round_wire[70]) );
  BUF_X4 \sha1_round/U296  ( .A(rnd_q[103]), .Z(sha1_round_wire[69]) );
  BUF_X4 \sha1_round/U295  ( .A(rnd_q[99]), .Z(sha1_round_wire[65]) );
  BUF_X4 \sha1_round/U294  ( .A(rnd_q[95]), .Z(sha1_round_wire[63]) );
  BUF_X4 \sha1_round/U293  ( .A(rnd_q[91]), .Z(sha1_round_wire[59]) );
  BUF_X4 \sha1_round/U292  ( .A(rnd_q[90]), .Z(sha1_round_wire[58]) );
  BUF_X4 \sha1_round/U291  ( .A(rnd_q[89]), .Z(sha1_round_wire[57]) );
  BUF_X4 \sha1_round/U290  ( .A(rnd_q[88]), .Z(sha1_round_wire[56]) );
  BUF_X4 \sha1_round/U289  ( .A(rnd_q[87]), .Z(sha1_round_wire[55]) );
  BUF_X4 \sha1_round/U288  ( .A(rnd_q[85]), .Z(sha1_round_wire[53]) );
  BUF_X4 \sha1_round/U287  ( .A(rnd_q[81]), .Z(sha1_round_wire[49]) );
  BUF_X4 \sha1_round/U286  ( .A(rnd_q[80]), .Z(sha1_round_wire[48]) );
  BUF_X4 \sha1_round/U285  ( .A(rnd_q[78]), .Z(sha1_round_wire[46]) );
  BUF_X4 \sha1_round/U284  ( .A(rnd_q[76]), .Z(sha1_round_wire[44]) );
  BUF_X4 \sha1_round/U283  ( .A(rnd_q[74]), .Z(sha1_round_wire[42]) );
  BUF_X4 \sha1_round/U282  ( .A(rnd_q[72]), .Z(sha1_round_wire[40]) );
  BUF_X4 \sha1_round/U281  ( .A(rnd_q[71]), .Z(sha1_round_wire[39]) );
  BUF_X4 \sha1_round/U280  ( .A(rnd_q[67]), .Z(sha1_round_wire[35]) );
  BUF_X4 \sha1_round/U279  ( .A(rnd_q[66]), .Z(sha1_round_wire[34]) );
  BUF_X4 \sha1_round/U278  ( .A(rnd_q[65]), .Z(sha1_round_wire[33]) );
  BUF_X4 \sha1_round/U277  ( .A(rnd_q[62]), .Z(sha1_round_wire[30]) );
  BUF_X4 \sha1_round/U276  ( .A(rnd_q[61]), .Z(sha1_round_wire[29]) );
  BUF_X4 \sha1_round/U275  ( .A(rnd_q[60]), .Z(sha1_round_wire[28]) );
  BUF_X4 \sha1_round/U274  ( .A(rnd_q[59]), .Z(sha1_round_wire[27]) );
  BUF_X4 \sha1_round/U273  ( .A(rnd_q[58]), .Z(sha1_round_wire[26]) );
  BUF_X4 \sha1_round/U272  ( .A(rnd_q[57]), .Z(sha1_round_wire[25]) );
  BUF_X4 \sha1_round/U271  ( .A(rnd_q[55]), .Z(sha1_round_wire[23]) );
  BUF_X4 \sha1_round/U270  ( .A(rnd_q[54]), .Z(sha1_round_wire[22]) );
  BUF_X4 \sha1_round/U269  ( .A(rnd_q[53]), .Z(sha1_round_wire[21]) );
  BUF_X4 \sha1_round/U268  ( .A(rnd_q[51]), .Z(sha1_round_wire[19]) );
  BUF_X4 \sha1_round/U267  ( .A(rnd_q[50]), .Z(sha1_round_wire[18]) );
  BUF_X4 \sha1_round/U266  ( .A(rnd_q[49]), .Z(sha1_round_wire[17]) );
  BUF_X4 \sha1_round/U265  ( .A(rnd_q[47]), .Z(sha1_round_wire[15]) );
  BUF_X4 \sha1_round/U264  ( .A(rnd_q[46]), .Z(sha1_round_wire[14]) );
  BUF_X4 \sha1_round/U263  ( .A(rnd_q[43]), .Z(sha1_round_wire[11]) );
  BUF_X4 \sha1_round/U262  ( .A(rnd_q[42]), .Z(sha1_round_wire[10]) );
  BUF_X4 \sha1_round/U261  ( .A(rnd_q[41]), .Z(sha1_round_wire[9]) );
  BUF_X4 \sha1_round/U260  ( .A(rnd_q[38]), .Z(sha1_round_wire[6]) );
  BUF_X4 \sha1_round/U259  ( .A(rnd_q[37]), .Z(sha1_round_wire[5]) );
  BUF_X4 \sha1_round/U258  ( .A(rnd_q[36]), .Z(sha1_round_wire[4]) );
  BUF_X4 \sha1_round/U257  ( .A(rnd_q[35]), .Z(sha1_round_wire[3]) );
  BUF_X4 \sha1_round/U256  ( .A(rnd_q[34]), .Z(sha1_round_wire[2]) );
  BUF_X4 \sha1_round/U255  ( .A(rnd_q[33]), .Z(sha1_round_wire[1]) );
  BUF_X4 \sha1_round/U254  ( .A(rnd_q[32]), .Z(sha1_round_wire[0]) );
  BUF_X4 \sha1_round/U253  ( .A(rnd_q[136]), .Z(sha1_round_wire[104]) );
  BUF_X4 \sha1_round/U252  ( .A(rnd_q[135]), .Z(sha1_round_wire[103]) );
  BUF_X4 \sha1_round/U251  ( .A(rnd_q[132]), .Z(sha1_round_wire[100]) );
  BUF_X4 \sha1_round/U250  ( .A(rnd_q[127]), .Z(sha1_round_wire[93]) );
  BUF_X4 \sha1_round/U249  ( .A(rnd_q[126]), .Z(sha1_round_wire[92]) );
  BUF_X4 \sha1_round/U248  ( .A(rnd_q[125]), .Z(sha1_round_wire[91]) );
  BUF_X4 \sha1_round/U247  ( .A(rnd_q[124]), .Z(sha1_round_wire[90]) );
  BUF_X4 \sha1_round/U246  ( .A(rnd_q[123]), .Z(sha1_round_wire[89]) );
  BUF_X4 \sha1_round/U245  ( .A(rnd_q[122]), .Z(sha1_round_wire[88]) );
  BUF_X4 \sha1_round/U244  ( .A(rnd_q[121]), .Z(sha1_round_wire[87]) );
  BUF_X4 \sha1_round/U243  ( .A(rnd_q[119]), .Z(sha1_round_wire[85]) );
  BUF_X4 \sha1_round/U242  ( .A(rnd_q[118]), .Z(sha1_round_wire[84]) );
  BUF_X4 \sha1_round/U241  ( .A(rnd_q[115]), .Z(sha1_round_wire[81]) );
  BUF_X4 \sha1_round/U240  ( .A(rnd_q[114]), .Z(sha1_round_wire[80]) );
  BUF_X4 \sha1_round/U239  ( .A(rnd_q[111]), .Z(sha1_round_wire[77]) );
  BUF_X4 \sha1_round/U238  ( .A(rnd_q[107]), .Z(sha1_round_wire[73]) );
  BUF_X4 \sha1_round/U237  ( .A(rnd_q[100]), .Z(sha1_round_wire[66]) );
  BUF_X4 \sha1_round/U236  ( .A(rnd_q[94]), .Z(sha1_round_wire[62]) );
  BUF_X4 \sha1_round/U235  ( .A(rnd_q[93]), .Z(sha1_round_wire[61]) );
  BUF_X4 \sha1_round/U234  ( .A(rnd_q[92]), .Z(sha1_round_wire[60]) );
  BUF_X4 \sha1_round/U233  ( .A(rnd_q[86]), .Z(sha1_round_wire[54]) );
  BUF_X4 \sha1_round/U232  ( .A(rnd_q[83]), .Z(sha1_round_wire[51]) );
  BUF_X4 \sha1_round/U231  ( .A(rnd_q[82]), .Z(sha1_round_wire[50]) );
  BUF_X4 \sha1_round/U230  ( .A(rnd_q[79]), .Z(sha1_round_wire[47]) );
  BUF_X4 \sha1_round/U229  ( .A(rnd_q[75]), .Z(sha1_round_wire[43]) );
  BUF_X4 \sha1_round/U228  ( .A(rnd_q[68]), .Z(sha1_round_wire[36]) );
  BUF_X4 \sha1_round/U227  ( .A(rnd_q[64]), .Z(sha1_round_wire[32]) );
  BUF_X4 \sha1_round/U226  ( .A(rnd_q[63]), .Z(sha1_round_wire[31]) );
  BUF_X4 \sha1_round/U225  ( .A(rnd_q[56]), .Z(sha1_round_wire[24]) );
  BUF_X4 \sha1_round/U224  ( .A(rnd_q[48]), .Z(sha1_round_wire[16]) );
  BUF_X4 \sha1_round/U223  ( .A(rnd_q[45]), .Z(sha1_round_wire[13]) );
  BUF_X4 \sha1_round/U222  ( .A(rnd_q[44]), .Z(sha1_round_wire[12]) );
  BUF_X4 \sha1_round/U221  ( .A(rnd_q[40]), .Z(sha1_round_wire[8]) );
  BUF_X4 \sha1_round/U220  ( .A(rnd_q[120]), .Z(sha1_round_wire[86]) );
  BUF_X4 \sha1_round/U219  ( .A(rnd_q[108]), .Z(sha1_round_wire[74]) );
  BUF_X4 \sha1_round/U218  ( .A(rnd_q[98]), .Z(sha1_round_wire[64]) );
  BUF_X4 \sha1_round/U217  ( .A(rnd_q[52]), .Z(sha1_round_wire[20]) );
  BUF_X4 \sha1_round/U216  ( .A(rnd_q[97]), .Z(sha1_round_wire[95]) );
  BUF_X4 \sha1_round/U215  ( .A(rnd_q[77]), .Z(sha1_round_wire[45]) );
  BUF_X4 \sha1_round/U214  ( .A(rnd_q[73]), .Z(sha1_round_wire[41]) );
  BUF_X4 \sha1_round/U213  ( .A(rnd_q[84]), .Z(sha1_round_wire[52]) );
  BUF_X4 \sha1_round/U212  ( .A(rnd_q[70]), .Z(sha1_round_wire[38]) );
  BUF_X4 \sha1_round/U211  ( .A(rnd_q[102]), .Z(sha1_round_wire[68]) );
  BUF_X4 \sha1_round/U210  ( .A(rnd_q[69]), .Z(sha1_round_wire[37]) );
  BUF_X4 \sha1_round/U209  ( .A(rnd_q[101]), .Z(sha1_round_wire[67]) );
  XOR2_X2 \sha1_round/U208  ( .A(rnd_q[118]), .B(rnd_q[86]), .Z(
        \sha1_round/n380 ) );
  XOR2_X2 \sha1_round/U207  ( .A(rnd_q[112]), .B(rnd_q[80]), .Z(
        \sha1_round/n379 ) );
  XOR2_X2 \sha1_round/U206  ( .A(rnd_q[108]), .B(rnd_q[76]), .Z(
        \sha1_round/n378 ) );
  XOR2_X2 \sha1_round/U205  ( .A(rnd_q[109]), .B(rnd_q[77]), .Z(
        \sha1_round/n377 ) );
  XOR2_X2 \sha1_round/U204  ( .A(rnd_q[113]), .B(rnd_q[81]), .Z(
        \sha1_round/n376 ) );
  XOR2_X2 \sha1_round/U203  ( .A(rnd_q[111]), .B(rnd_q[79]), .Z(
        \sha1_round/n375 ) );
  XOR2_X2 \sha1_round/U202  ( .A(rnd_q[100]), .B(rnd_q[68]), .Z(
        \sha1_round/n374 ) );
  XOR2_X2 \sha1_round/U201  ( .A(rnd_q[114]), .B(rnd_q[82]), .Z(
        \sha1_round/n373 ) );
  XOR2_X2 \sha1_round/U200  ( .A(rnd_q[107]), .B(rnd_q[75]), .Z(
        \sha1_round/n372 ) );
  XOR2_X2 \sha1_round/U199  ( .A(rnd_q[115]), .B(rnd_q[83]), .Z(
        \sha1_round/n371 ) );
  XOR2_X2 \sha1_round/U198  ( .A(rnd_q[104]), .B(rnd_q[72]), .Z(
        \sha1_round/n370 ) );
  XOR2_X2 \sha1_round/U197  ( .A(rnd_q[117]), .B(rnd_q[85]), .Z(
        \sha1_round/n369 ) );
  XOR2_X2 \sha1_round/U196  ( .A(rnd_q[110]), .B(rnd_q[78]), .Z(
        \sha1_round/n368 ) );
  XOR2_X2 \sha1_round/U195  ( .A(rnd_q[106]), .B(rnd_q[74]), .Z(
        \sha1_round/n367 ) );
  XOR2_X2 \sha1_round/U194  ( .A(rnd_q[116]), .B(rnd_q[84]), .Z(
        \sha1_round/n366 ) );
  XOR2_X2 \sha1_round/U193  ( .A(rnd_q[101]), .B(rnd_q[69]), .Z(
        \sha1_round/n365 ) );
  NAND2_X1 \sha1_round/U192  ( .A1(\sha1_round/n365 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n752 ) );
  NAND2_X4 \sha1_round/U191  ( .A1(\sha1_round/n819 ), .A2(\sha1_round/n820 ), 
        .ZN(\sha1_round/n767 ) );
  NAND2_X1 \sha1_round/U190  ( .A1(\sha1_round/n3120 ), .A2(\sha1_round/n820 ), 
        .ZN(\sha1_round/n3170 ) );
  INV_X2 \sha1_round/U189  ( .A(\sha1_round/n360 ), .ZN(\sha1_round/n363 ) );
  INV_X4 \sha1_round/U188  ( .A(\sha1_round/n3140 ), .ZN(\sha1_round/n510 ) );
  INV_X4 \sha1_round/U187  ( .A(\sha1_round/n363 ), .ZN(\sha1_round/n364 ) );
  NAND3_X1 \sha1_round/U186  ( .A1(rnd_q[64]), .A2(rnd_q[96]), .A3(
        \sha1_round/k[3] ), .ZN(\sha1_round/n815 ) );
  OR2_X4 \sha1_round/U185  ( .A1(rnd_q[73]), .A2(rnd_q[105]), .ZN(
        \sha1_round/n362 ) );
  NAND2_X4 \sha1_round/U184  ( .A1(\sha1_round/n712 ), .A2(\sha1_round/n713 ), 
        .ZN(\sha1_round/f [11]) );
  NAND2_X4 \sha1_round/U183  ( .A1(\sha1_round/n721 ), .A2(\sha1_round/n720 ), 
        .ZN(\sha1_round/f [10]) );
  NAND2_X4 \sha1_round/U182  ( .A1(\sha1_round/n753 ), .A2(\sha1_round/n754 ), 
        .ZN(\sha1_round/f [5]) );
  NOR2_X1 \sha1_round/U180  ( .A1(\sha1_round/n706 ), .A2(\sha1_round/n3120 ), 
        .ZN(\sha1_round/n708 ) );
  NOR2_X1 \sha1_round/U179  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n3210 ), 
        .ZN(\sha1_round/n722 ) );
  NOR2_X1 \sha1_round/U177  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n3240 ), 
        .ZN(\sha1_round/n738 ) );
  NAND2_X1 \sha1_round/U176  ( .A1(\sha1_round/n372 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n711 ) );
  INV_X4 \sha1_round/U175  ( .A(rnd_q[43]), .ZN(\sha1_round/n357 ) );
  NAND2_X2 \sha1_round/U174  ( .A1(\sha1_round/n711 ), .A2(\sha1_round/n357 ), 
        .ZN(\sha1_round/n358 ) );
  NAND2_X2 \sha1_round/U173  ( .A1(\sha1_round/n3230 ), .A2(\sha1_round/n532 ), 
        .ZN(\sha1_round/n533 ) );
  NAND2_X2 \sha1_round/U172  ( .A1(\sha1_round/n367 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n719 ) );
  INV_X1 \sha1_round/U170  ( .A(rnd_q[42]), .ZN(\sha1_round/n354 ) );
  NAND2_X2 \sha1_round/U169  ( .A1(\sha1_round/n719 ), .A2(\sha1_round/n354 ), 
        .ZN(\sha1_round/n355 ) );
  NAND2_X1 \sha1_round/U167  ( .A1(\sha1_round/n3220 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n747 ) );
  INV_X1 \sha1_round/U166  ( .A(rnd_q[38]), .ZN(\sha1_round/n351 ) );
  NAND2_X2 \sha1_round/U165  ( .A1(\sha1_round/n747 ), .A2(\sha1_round/n351 ), 
        .ZN(\sha1_round/n352 ) );
  INV_X1 \sha1_round/U164  ( .A(rnd_q[41]), .ZN(\sha1_round/n348 ) );
  NAND2_X2 \sha1_round/U163  ( .A1(\sha1_round/n726 ), .A2(\sha1_round/n348 ), 
        .ZN(\sha1_round/n349 ) );
  INV_X1 \sha1_round/U162  ( .A(rnd_q[37]), .ZN(\sha1_round/n3450 ) );
  NAND2_X2 \sha1_round/U160  ( .A1(\sha1_round/n752 ), .A2(\sha1_round/n3450 ), 
        .ZN(\sha1_round/n3460 ) );
  NAND3_X1 \sha1_round/U159  ( .A1(rnd_q[65]), .A2(rnd_q[97]), .A3(
        \sha1_round/k[3] ), .ZN(\sha1_round/n802 ) );
  NAND2_X4 \sha1_round/U157  ( .A1(\sha1_round/n3250 ), .A2(\sha1_round/n800 ), 
        .ZN(\sha1_round/f [1]) );
  NOR2_X1 \sha1_round/U156  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n369 ), 
        .ZN(\sha1_round/n627 ) );
  NOR2_X1 \sha1_round/U155  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n373 ), 
        .ZN(\sha1_round/n651 ) );
  NAND3_X1 \sha1_round/U154  ( .A1(rnd_q[67]), .A2(rnd_q[99]), .A3(
        \sha1_round/k[3] ), .ZN(\sha1_round/n776 ) );
  NAND3_X1 \sha1_round/U153  ( .A1(rnd_q[66]), .A2(rnd_q[98]), .A3(
        \sha1_round/k[3] ), .ZN(\sha1_round/n789 ) );
  AND2_X2 \sha1_round/U152  ( .A1(\sha1_round/n3150 ), .A2(\sha1_round/n362 ), 
        .ZN(\sha1_round/n723 ) );
  NAND2_X1 \sha1_round/U150  ( .A1(\sha1_round/n3150 ), .A2(\sha1_round/n796 ), 
        .ZN(\sha1_round/n797 ) );
  NOR2_X2 \sha1_round/U149  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n367 ), 
        .ZN(\sha1_round/n715 ) );
  NOR2_X2 \sha1_round/U147  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n372 ), 
        .ZN(\sha1_round/n707 ) );
  INV_X2 \sha1_round/U146  ( .A(\sha1_round/n3170 ), .ZN(\sha1_round/n817 ) );
  NAND2_X4 \sha1_round/U145  ( .A1(\sha1_round/n736 ), .A2(\sha1_round/n735 ), 
        .ZN(\sha1_round/f [8]) );
  OR2_X2 \sha1_round/U144  ( .A1(\sha1_round/n750 ), .A2(\sha1_round/n3120 ), 
        .ZN(\sha1_round/n3420 ) );
  OR2_X4 \sha1_round/U143  ( .A1(rnd_q[101]), .A2(\sha1_round/n510 ), .ZN(
        \sha1_round/n3410 ) );
  AND3_X4 \sha1_round/U142  ( .A1(\sha1_round/n3410 ), .A2(\sha1_round/n3420 ), 
        .A3(\sha1_round/n3430 ), .ZN(\sha1_round/n751 ) );
  NAND2_X4 \sha1_round/U140  ( .A1(\sha1_round/n697 ), .A2(\sha1_round/n696 ), 
        .ZN(\sha1_round/f [13]) );
  NAND2_X2 \sha1_round/U139  ( .A1(\sha1_round/n531 ), .A2(\sha1_round/n524 ), 
        .ZN(\sha1_round/n522 ) );
  NAND2_X2 \sha1_round/U137  ( .A1(\sha1_round/n524 ), .A2(\sha1_round/n523 ), 
        .ZN(\sha1_round/n526 ) );
  OR2_X1 \sha1_round/U136  ( .A1(\sha1_round/n745 ), .A2(\sha1_round/n3160 ), 
        .ZN(\sha1_round/n3390 ) );
  OR2_X1 \sha1_round/U135  ( .A1(rnd_q[102]), .A2(\sha1_round/n510 ), .ZN(
        \sha1_round/n3380 ) );
  AND3_X4 \sha1_round/U134  ( .A1(\sha1_round/n3380 ), .A2(\sha1_round/n3390 ), 
        .A3(\sha1_round/n3400 ), .ZN(\sha1_round/n746 ) );
  NAND2_X2 \sha1_round/U133  ( .A1(\sha1_round/n3150 ), .A2(\sha1_round/n770 ), 
        .ZN(\sha1_round/n771 ) );
  INV_X2 \sha1_round/U132  ( .A(rnd_q[33]), .ZN(\sha1_round/n791 ) );
  NOR2_X2 \sha1_round/U130  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n374 ), 
        .ZN(\sha1_round/n757 ) );
  NOR2_X2 \sha1_round/U129  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n379 ), 
        .ZN(\sha1_round/n667 ) );
  NOR2_X2 \sha1_round/U127  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n375 ), 
        .ZN(\sha1_round/n675 ) );
  INV_X1 \sha1_round/U126  ( .A(\sha1_round/n819 ), .ZN(\sha1_round/n825 ) );
  OR2_X2 \sha1_round/U125  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n3220 ), 
        .ZN(\sha1_round/n3400 ) );
  OR2_X2 \sha1_round/U124  ( .A1(\sha1_round/n756 ), .A2(\sha1_round/n365 ), 
        .ZN(\sha1_round/n3430 ) );
  NAND2_X1 \sha1_round/U123  ( .A1(rnd_cnt_q[6]), .A2(rnd_cnt_q[5]), .ZN(
        \sha1_round/n535 ) );
  NAND3_X2 \sha1_round/U122  ( .A1(rnd_cnt_q[5]), .A2(\sha1_round/n531 ), .A3(
        \sha1_round/n524 ), .ZN(\sha1_round/n528 ) );
  NAND2_X1 \sha1_round/U120  ( .A1(\sha1_round/n370 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n734 ) );
  NAND2_X1 \sha1_round/U119  ( .A1(\sha1_round/n366 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n639 ) );
  NAND2_X2 \sha1_round/U117  ( .A1(\sha1_round/n3210 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n726 ) );
  NAND2_X1 \sha1_round/U116  ( .A1(\sha1_round/n368 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n687 ) );
  NAND2_X1 \sha1_round/U115  ( .A1(\sha1_round/n371 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n647 ) );
  NAND2_X1 \sha1_round/U114  ( .A1(\sha1_round/n379 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n671 ) );
  NAND2_X1 \sha1_round/U113  ( .A1(\sha1_round/n375 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n679 ) );
  NAND2_X1 \sha1_round/U112  ( .A1(\sha1_round/n378 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n703 ) );
  NAND3_X1 \sha1_round/U111  ( .A1(rnd_q[34]), .A2(\sha1_round/n515 ), .A3(
        \sha1_round/n780 ), .ZN(\sha1_round/n788 ) );
  NAND2_X1 \sha1_round/U110  ( .A1(\sha1_round/n377 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n695 ) );
  NAND3_X1 \sha1_round/U109  ( .A1(\sha1_round/n779 ), .A2(\sha1_round/n778 ), 
        .A3(\sha1_round/n515 ), .ZN(\sha1_round/n790 ) );
  NAND2_X1 \sha1_round/U108  ( .A1(\sha1_round/n369 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n631 ) );
  NAND2_X1 \sha1_round/U107  ( .A1(\sha1_round/n168 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n612 ) );
  NAND2_X1 \sha1_round/U106  ( .A1(\sha1_round/n373 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n655 ) );
  NAND2_X1 \sha1_round/U105  ( .A1(\sha1_round/n159 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n603 ) );
  NAND2_X1 \sha1_round/U104  ( .A1(\sha1_round/n376 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n663 ) );
  NAND2_X1 \sha1_round/U103  ( .A1(\sha1_round/n380 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n623 ) );
  INV_X1 \sha1_round/U102  ( .A(rnd_q[40]), .ZN(\sha1_round/n3340 ) );
  NAND2_X2 \sha1_round/U100  ( .A1(\sha1_round/n734 ), .A2(\sha1_round/n3340 ), 
        .ZN(\sha1_round/n3350 ) );
  NAND2_X4 \sha1_round/U99  ( .A1(\sha1_round/n705 ), .A2(\sha1_round/n704 ), 
        .ZN(\sha1_round/f [12]) );
  NOR2_X2 \sha1_round/U97  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n377 ), 
        .ZN(\sha1_round/n691 ) );
  NAND2_X2 \sha1_round/U96  ( .A1(\sha1_round/n3270 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n814 ) );
  INV_X4 \sha1_round/U95  ( .A(rnd_q[39]), .ZN(\sha1_round/n3440 ) );
  NAND2_X1 \sha1_round/U94  ( .A1(\sha1_round/n3240 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n742 ) );
  INV_X4 \sha1_round/U93  ( .A(\sha1_round/n3440 ), .ZN(sha1_round_wire[7]) );
  NAND2_X2 \sha1_round/U92  ( .A1(\sha1_round/n742 ), .A2(\sha1_round/n3440 ), 
        .ZN(\sha1_round/n3330 ) );
  NAND2_X2 \sha1_round/U90  ( .A1(\sha1_round/n741 ), .A2(sha1_round_wire[7]), 
        .ZN(\sha1_round/n3320 ) );
  INV_X4 \sha1_round/U89  ( .A(\sha1_round/k[3] ), .ZN(\sha1_round/n518 ) );
  INV_X2 \sha1_round/U87  ( .A(\sha1_round/n518 ), .ZN(\sha1_round/n3300 ) );
  INV_X4 \sha1_round/U86  ( .A(rnd_cnt_q[5]), .ZN(\sha1_round/n525 ) );
  AND2_X4 \sha1_round/U85  ( .A1(\sha1_round/n804 ), .A2(\sha1_round/n805 ), 
        .ZN(\sha1_round/n3290 ) );
  AND2_X4 \sha1_round/U84  ( .A1(\sha1_round/n791 ), .A2(\sha1_round/n792 ), 
        .ZN(\sha1_round/n3280 ) );
  AND2_X4 \sha1_round/U83  ( .A1(rnd_q[32]), .A2(\sha1_round/n806 ), .ZN(
        \sha1_round/n3270 ) );
  OR2_X2 \sha1_round/U82  ( .A1(\sha1_round/n723 ), .A2(\sha1_round/n724 ), 
        .ZN(\sha1_round/n3260 ) );
  XOR2_X2 \sha1_round/U81  ( .A(rnd_q[103]), .B(rnd_q[71]), .Z(
        \sha1_round/n3240 ) );
  AND2_X4 \sha1_round/U80  ( .A1(n7119), .A2(rnd_cnt_q[5]), .ZN(
        \sha1_round/n3230 ) );
  XOR2_X2 \sha1_round/U79  ( .A(rnd_q[102]), .B(rnd_q[70]), .Z(
        \sha1_round/n3220 ) );
  XOR2_X2 \sha1_round/U78  ( .A(rnd_q[105]), .B(rnd_q[73]), .Z(
        \sha1_round/n3210 ) );
  BUF_X4 \sha1_round/U77  ( .A(\sha1_round/n515 ), .Z(\sha1_round/n3370 ) );
  NAND2_X1 \sha1_round/U76  ( .A1(n7119), .A2(rnd_cnt_q[4]), .ZN(
        \sha1_round/n519 ) );
  NAND2_X4 \sha1_round/U75  ( .A1(\sha1_round/n358 ), .A2(\sha1_round/n359 ), 
        .ZN(\sha1_round/n712 ) );
  NAND2_X2 \sha1_round/U74  ( .A1(\sha1_round/n532 ), .A2(n7119), .ZN(
        \sha1_round/n521 ) );
  NAND3_X2 \sha1_round/U73  ( .A1(rnd_q[33]), .A2(\sha1_round/n515 ), .A3(
        \sha1_round/n793 ), .ZN(\sha1_round/n801 ) );
  NAND2_X2 \sha1_round/U72  ( .A1(\sha1_round/n641 ), .A2(\sha1_round/n640 ), 
        .ZN(\sha1_round/f [20]) );
  NAND2_X2 \sha1_round/U71  ( .A1(\sha1_round/n689 ), .A2(\sha1_round/n688 ), 
        .ZN(\sha1_round/f [14]) );
  NAND2_X2 \sha1_round/U70  ( .A1(\sha1_round/n510 ), .A2(\sha1_round/n817 ), 
        .ZN(\sha1_round/n2 ) );
  NAND2_X2 \sha1_round/U69  ( .A1(rnd_q[33]), .A2(\sha1_round/n799 ), .ZN(
        \sha1_round/n800 ) );
  NAND2_X2 \sha1_round/U68  ( .A1(rnd_q[35]), .A2(\sha1_round/n773 ), .ZN(
        \sha1_round/n774 ) );
  NAND2_X2 \sha1_round/U67  ( .A1(\sha1_round/n718 ), .A2(rnd_q[42]), .ZN(
        \sha1_round/n356 ) );
  NAND2_X2 \sha1_round/U66  ( .A1(\sha1_round/n733 ), .A2(rnd_q[40]), .ZN(
        \sha1_round/n3360 ) );
  NOR2_X2 \sha1_round/U65  ( .A1(\sha1_round/n722 ), .A2(\sha1_round/n3260 ), 
        .ZN(\sha1_round/n725 ) );
  NAND2_X2 \sha1_round/U64  ( .A1(\sha1_round/n725 ), .A2(rnd_q[41]), .ZN(
        \sha1_round/n350 ) );
  NAND2_X2 \sha1_round/U63  ( .A1(\sha1_round/n746 ), .A2(rnd_q[38]), .ZN(
        \sha1_round/n353 ) );
  NOR3_X2 \sha1_round/U62  ( .A1(\sha1_round/n709 ), .A2(\sha1_round/n708 ), 
        .A3(\sha1_round/n707 ), .ZN(\sha1_round/n710 ) );
  NAND2_X2 \sha1_round/U61  ( .A1(\sha1_round/n349 ), .A2(\sha1_round/n350 ), 
        .ZN(\sha1_round/n727 ) );
  NOR2_X2 \sha1_round/U60  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n366 ), 
        .ZN(\sha1_round/n635 ) );
  INV_X1 \sha1_round/U59  ( .A(\sha1_round/n514 ), .ZN(\sha1_round/n360 ) );
  INV_X8 \sha1_round/U58  ( .A(\sha1_round/n512 ), .ZN(\sha1_round/n514 ) );
  NAND4_X4 \sha1_round/U57  ( .A1(\sha1_round/n777 ), .A2(\sha1_round/n776 ), 
        .A3(\sha1_round/n775 ), .A4(\sha1_round/n774 ), .ZN(\sha1_round/f [3])
         );
  NOR2_X1 \sha1_round/U56  ( .A1(rnd_q[107]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n709 ) );
  NOR2_X1 \sha1_round/U55  ( .A1(rnd_q[116]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n637 ) );
  NOR2_X1 \sha1_round/U54  ( .A1(rnd_q[104]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n732 ) );
  NOR2_X1 \sha1_round/U53  ( .A1(rnd_q[115]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n645 ) );
  NOR2_X1 \sha1_round/U52  ( .A1(rnd_q[108]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n701 ) );
  NOR2_X1 \sha1_round/U51  ( .A1(rnd_q[117]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n629 ) );
  NOR2_X1 \sha1_round/U50  ( .A1(rnd_q[113]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n661 ) );
  NOR2_X1 \sha1_round/U49  ( .A1(rnd_q[118]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n621 ) );
  NOR2_X1 \sha1_round/U48  ( .A1(rnd_q[114]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n653 ) );
  NAND2_X4 \sha1_round/U47  ( .A1(\sha1_round/n352 ), .A2(\sha1_round/n353 ), 
        .ZN(\sha1_round/n748 ) );
  INV_X8 \sha1_round/U46  ( .A(\sha1_round/n767 ), .ZN(\sha1_round/n756 ) );
  INV_X4 \sha1_round/U45  ( .A(n7119), .ZN(\sha1_round/n523 ) );
  NAND4_X2 \sha1_round/U44  ( .A1(\sha1_round/n521 ), .A2(\sha1_round/n529 ), 
        .A3(\sha1_round/n522 ), .A4(rnd_cnt_q[5]), .ZN(\sha1_round/n822 ) );
  NAND3_X2 \sha1_round/U43  ( .A1(\sha1_round/n525 ), .A2(\sha1_round/n526 ), 
        .A3(rnd_cnt_q[4]), .ZN(\sha1_round/n527 ) );
  NAND2_X2 \sha1_round/U42  ( .A1(\sha1_round/n528 ), .A2(\sha1_round/n527 ), 
        .ZN(\sha1_round/n530 ) );
  AND4_X4 \sha1_round/U41  ( .A1(\sha1_round/n520 ), .A2(\sha1_round/n529 ), 
        .A3(\sha1_round/n519 ), .A4(\sha1_round/n525 ), .ZN(\sha1_round/n3140 ) );
  INV_X4 \sha1_round/U40  ( .A(\sha1_round/n508 ), .ZN(\sha1_round/n509 ) );
  NAND3_X2 \sha1_round/U39  ( .A1(\sha1_round/n3130 ), .A2(\sha1_round/n815 ), 
        .A3(\sha1_round/n813 ), .ZN(\sha1_round/f [0]) );
  INV_X4 \sha1_round/U38  ( .A(rnd_cnt_q[6]), .ZN(\sha1_round/n529 ) );
  INV_X4 \sha1_round/U37  ( .A(\sha1_round/n3150 ), .ZN(\sha1_round/n3160 ) );
  INV_X8 \sha1_round/U36  ( .A(\sha1_round/n3160 ), .ZN(\sha1_round/n512 ) );
  INV_X8 \sha1_round/U35  ( .A(\sha1_round/n518 ), .ZN(\sha1_round/n517 ) );
  NAND2_X2 \sha1_round/U34  ( .A1(\sha1_round/n762 ), .A2(\sha1_round/n763 ), 
        .ZN(\sha1_round/f [4]) );
  NAND4_X2 \sha1_round/U33  ( .A1(\sha1_round/n790 ), .A2(\sha1_round/n788 ), 
        .A3(\sha1_round/n789 ), .A4(\sha1_round/n787 ), .ZN(\sha1_round/f [2])
         );
  NAND2_X2 \sha1_round/U32  ( .A1(\sha1_round/n355 ), .A2(\sha1_round/n356 ), 
        .ZN(\sha1_round/n720 ) );
  NAND2_X2 \sha1_round/U31  ( .A1(\sha1_round/n3320 ), .A2(\sha1_round/n3330 ), 
        .ZN(\sha1_round/n743 ) );
  NAND2_X2 \sha1_round/U30  ( .A1(\sha1_round/n744 ), .A2(\sha1_round/n743 ), 
        .ZN(\sha1_round/f [7]) );
  NAND2_X2 \sha1_round/U29  ( .A1(\sha1_round/n710 ), .A2(rnd_q[43]), .ZN(
        \sha1_round/n359 ) );
  NOR2_X2 \sha1_round/U28  ( .A1(\sha1_round/n516 ), .A2(\sha1_round/n370 ), 
        .ZN(\sha1_round/n730 ) );
  INV_X8 \sha1_round/U27  ( .A(\sha1_round/n3140 ), .ZN(\sha1_round/n361 ) );
  NOR2_X2 \sha1_round/U26  ( .A1(rnd_q[109]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n693 ) );
  NOR2_X2 \sha1_round/U25  ( .A1(rnd_q[110]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n685 ) );
  NOR2_X2 \sha1_round/U24  ( .A1(rnd_q[111]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n677 ) );
  NOR2_X1 \sha1_round/U23  ( .A1(rnd_q[105]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n724 ) );
  NOR2_X2 \sha1_round/U22  ( .A1(rnd_q[112]), .A2(\sha1_round/n361 ), .ZN(
        \sha1_round/n669 ) );
  INV_X16 \sha1_round/U21  ( .A(\sha1_round/n361 ), .ZN(\sha1_round/n511 ) );
  INV_X8 \sha1_round/U20  ( .A(\sha1_round/n822 ), .ZN(\sha1_round/n3150 ) );
  INV_X2 \sha1_round/U19  ( .A(\sha1_round/n512 ), .ZN(\sha1_round/n3200 ) );
  INV_X2 \sha1_round/U18  ( .A(\sha1_round/n512 ), .ZN(\sha1_round/n513 ) );
  INV_X2 \sha1_round/U17  ( .A(\sha1_round/n512 ), .ZN(\sha1_round/n3190 ) );
  INV_X4 \sha1_round/U16  ( .A(\sha1_round/n3150 ), .ZN(\sha1_round/n3180 ) );
  NAND4_X2 \sha1_round/U15  ( .A1(\sha1_round/n521 ), .A2(\sha1_round/n529 ), 
        .A3(\sha1_round/n522 ), .A4(rnd_cnt_q[5]), .ZN(\sha1_round/n3120 ) );
  INV_X8 \sha1_round/U14  ( .A(rnd_cnt_q[4]), .ZN(\sha1_round/n531 ) );
  NAND2_X4 \sha1_round/U13  ( .A1(rnd_cnt_q[3]), .A2(rnd_cnt_q[4]), .ZN(
        \sha1_round/n520 ) );
  NOR3_X4 \sha1_round/U12  ( .A1(\sha1_round/n717 ), .A2(\sha1_round/n716 ), 
        .A3(\sha1_round/n715 ), .ZN(\sha1_round/n718 ) );
  NAND2_X2 \sha1_round/U11  ( .A1(\sha1_round/n3280 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n803 ) );
  NOR3_X4 \sha1_round/U10  ( .A1(\sha1_round/n732 ), .A2(\sha1_round/n731 ), 
        .A3(\sha1_round/n730 ), .ZN(\sha1_round/n733 ) );
  NAND2_X2 \sha1_round/U9  ( .A1(\sha1_round/n3350 ), .A2(\sha1_round/n3360 ), 
        .ZN(\sha1_round/n735 ) );
  AND3_X4 \sha1_round/U8  ( .A1(\sha1_round/n801 ), .A2(\sha1_round/n803 ), 
        .A3(\sha1_round/n802 ), .ZN(\sha1_round/n3250 ) );
  NAND2_X2 \sha1_round/U7  ( .A1(\sha1_round/n3290 ), .A2(\sha1_round/n515 ), 
        .ZN(\sha1_round/n816 ) );
  AND2_X2 \sha1_round/U6  ( .A1(\sha1_round/n816 ), .A2(\sha1_round/n814 ), 
        .ZN(\sha1_round/n3130 ) );
  NAND2_X4 \sha1_round/U5  ( .A1(\sha1_round/n751 ), .A2(rnd_q[37]), .ZN(
        \sha1_round/n3470 ) );
  NAND2_X4 \sha1_round/U3  ( .A1(\sha1_round/n3470 ), .A2(\sha1_round/n3460 ), 
        .ZN(\sha1_round/n753 ) );
  XNOR2_X2 \sha1_round/U181  ( .A(rnd_q[87]), .B(rnd_q[119]), .ZN(
        \sha1_round/n168 ) );
  OR2_X2 \sha1_round/U178  ( .A1(rnd_q[87]), .A2(rnd_q[119]), .ZN(
        \sha1_round/n167 ) );
  XNOR2_X2 \sha1_round/U171  ( .A(rnd_q[88]), .B(rnd_q[120]), .ZN(
        \sha1_round/n159 ) );
  OR2_X2 \sha1_round/U168  ( .A1(rnd_q[88]), .A2(rnd_q[120]), .ZN(
        \sha1_round/n158 ) );
  XNOR2_X2 \sha1_round/U161  ( .A(rnd_q[89]), .B(rnd_q[121]), .ZN(
        \sha1_round/n150 ) );
  OR2_X2 \sha1_round/U158  ( .A1(rnd_q[89]), .A2(rnd_q[121]), .ZN(
        \sha1_round/n149 ) );
  XNOR2_X2 \sha1_round/U151  ( .A(rnd_q[90]), .B(rnd_q[122]), .ZN(
        \sha1_round/n141 ) );
  OR2_X2 \sha1_round/U148  ( .A1(rnd_q[90]), .A2(rnd_q[122]), .ZN(
        \sha1_round/n140 ) );
  XNOR2_X2 \sha1_round/U141  ( .A(rnd_q[91]), .B(rnd_q[123]), .ZN(
        \sha1_round/n132 ) );
  OR2_X2 \sha1_round/U138  ( .A1(rnd_q[91]), .A2(rnd_q[123]), .ZN(
        \sha1_round/n131 ) );
  XNOR2_X2 \sha1_round/U131  ( .A(rnd_q[92]), .B(rnd_q[124]), .ZN(
        \sha1_round/n123 ) );
  OR2_X2 \sha1_round/U128  ( .A1(rnd_q[92]), .A2(rnd_q[124]), .ZN(
        \sha1_round/n122 ) );
  XNOR2_X2 \sha1_round/U121  ( .A(rnd_q[93]), .B(rnd_q[125]), .ZN(
        \sha1_round/n114 ) );
  OR2_X2 \sha1_round/U118  ( .A1(rnd_q[93]), .A2(rnd_q[125]), .ZN(
        \sha1_round/n113 ) );
  XNOR2_X2 \sha1_round/U101  ( .A(rnd_q[94]), .B(rnd_q[126]), .ZN(
        \sha1_round/n96 ) );
  OR2_X2 \sha1_round/U98  ( .A1(rnd_q[94]), .A2(rnd_q[126]), .ZN(
        \sha1_round/n95 ) );
  XNOR2_X2 \sha1_round/U91  ( .A(rnd_q[95]), .B(rnd_q[127]), .ZN(
        \sha1_round/n87 ) );
  OR2_X2 \sha1_round/U88  ( .A1(rnd_q[95]), .A2(rnd_q[127]), .ZN(
        \sha1_round/n86 ) );
  NAND2_X2 \sha1_round/add_79_4/U377  ( .A1(\sha1_round/N316 ), .A2(rnd_q[155]), .ZN(\sha1_round/add_79_4/n243 ) );
  INV_X4 \sha1_round/add_79_4/U376  ( .A(\sha1_round/add_79_4/n56 ), .ZN(
        \sha1_round/add_79_4/n311 ) );
  NAND4_X2 \sha1_round/add_79_4/U375  ( .A1(\sha1_round/N320 ), .A2(rnd_q[159]), .A3(\sha1_round/add_79_4/n336 ), .A4(\sha1_round/add_79_4/n72 ), .ZN(
        \sha1_round/add_79_4/n341 ) );
  NAND2_X2 \sha1_round/add_79_4/U374  ( .A1(\sha1_round/N322 ), .A2(rnd_q[129]), .ZN(\sha1_round/add_79_4/n70 ) );
  INV_X4 \sha1_round/add_79_4/U373  ( .A(\sha1_round/add_79_4/n70 ), .ZN(
        \sha1_round/add_79_4/n344 ) );
  INV_X4 \sha1_round/add_79_4/U372  ( .A(\sha1_round/add_79_4/n67 ), .ZN(
        \sha1_round/add_79_4/n345 ) );
  NAND2_X2 \sha1_round/add_79_4/U371  ( .A1(\sha1_round/add_79_4/n316 ), .A2(
        \sha1_round/add_79_4/n68 ), .ZN(\sha1_round/add_79_4/n280 ) );
  INV_X4 \sha1_round/add_79_4/U370  ( .A(\sha1_round/add_79_4/n280 ), .ZN(
        \sha1_round/add_79_4/n62 ) );
  INV_X4 \sha1_round/add_79_4/U369  ( .A(\sha1_round/add_79_4/n60 ), .ZN(
        \sha1_round/add_79_4/n318 ) );
  NAND2_X2 \sha1_round/add_79_4/U368  ( .A1(\sha1_round/add_79_4/n62 ), .A2(
        \sha1_round/add_79_4/n318 ), .ZN(\sha1_round/add_79_4/n329 ) );
  INV_X4 \sha1_round/add_79_4/U367  ( .A(\sha1_round/add_79_4/n75 ), .ZN(
        \sha1_round/add_79_4/n336 ) );
  INV_X4 \sha1_round/add_79_4/U366  ( .A(\sha1_round/add_79_4/n80 ), .ZN(
        \sha1_round/add_79_4/n337 ) );
  INV_X4 \sha1_round/add_79_4/U365  ( .A(\sha1_round/add_79_4/n72 ), .ZN(
        \sha1_round/add_79_4/n339 ) );
  INV_X4 \sha1_round/add_79_4/U364  ( .A(\sha1_round/add_79_4/n64 ), .ZN(
        \sha1_round/add_79_4/n314 ) );
  NAND2_X2 \sha1_round/add_79_4/U363  ( .A1(\sha1_round/N319 ), .A2(rnd_q[158]), .ZN(\sha1_round/add_79_4/n86 ) );
  INV_X4 \sha1_round/add_79_4/U362  ( .A(\sha1_round/add_79_4/n90 ), .ZN(
        \sha1_round/add_79_4/n335 ) );
  NAND2_X2 \sha1_round/add_79_4/U361  ( .A1(\sha1_round/add_79_4/n243 ), .A2(
        \sha1_round/add_79_4/n139 ), .ZN(\sha1_round/add_79_4/n333 ) );
  INV_X4 \sha1_round/add_79_4/U360  ( .A(\sha1_round/add_79_4/n85 ), .ZN(
        \sha1_round/add_79_4/n332 ) );
  NAND2_X2 \sha1_round/add_79_4/U359  ( .A1(\sha1_round/N318 ), .A2(rnd_q[157]), .ZN(\sha1_round/add_79_4/n87 ) );
  NAND2_X2 \sha1_round/add_79_4/U358  ( .A1(\sha1_round/add_79_4/n311 ), .A2(
        \sha1_round/add_79_4/n54 ), .ZN(\sha1_round/add_79_4/n328 ) );
  NAND2_X2 \sha1_round/add_79_4/U357  ( .A1(\sha1_round/N325 ), .A2(rnd_q[132]), .ZN(\sha1_round/add_79_4/n55 ) );
  NAND2_X2 \sha1_round/add_79_4/U356  ( .A1(\sha1_round/add_79_4/n328 ), .A2(
        \sha1_round/add_79_4/n55 ), .ZN(\sha1_round/add_79_4/n324 ) );
  INV_X4 \sha1_round/add_79_4/U355  ( .A(\sha1_round/N326 ), .ZN(
        \sha1_round/add_79_4/n326 ) );
  INV_X4 \sha1_round/add_79_4/U354  ( .A(rnd_q[133]), .ZN(
        \sha1_round/add_79_4/n327 ) );
  NAND2_X2 \sha1_round/add_79_4/U353  ( .A1(\sha1_round/N326 ), .A2(rnd_q[133]), .ZN(\sha1_round/add_79_4/n308 ) );
  NAND2_X2 \sha1_round/add_79_4/U352  ( .A1(\sha1_round/add_79_4/n313 ), .A2(
        \sha1_round/add_79_4/n308 ), .ZN(\sha1_round/add_79_4/n325 ) );
  XNOR2_X2 \sha1_round/add_79_4/U351  ( .A(\sha1_round/add_79_4/n324 ), .B(
        \sha1_round/add_79_4/n325 ), .ZN(sha1_round_wire[138]) );
  NAND2_X2 \sha1_round/add_79_4/U350  ( .A1(\sha1_round/add_79_4/n324 ), .A2(
        \sha1_round/add_79_4/n313 ), .ZN(\sha1_round/add_79_4/n323 ) );
  NAND2_X2 \sha1_round/add_79_4/U349  ( .A1(\sha1_round/add_79_4/n308 ), .A2(
        \sha1_round/add_79_4/n323 ), .ZN(\sha1_round/add_79_4/n319 ) );
  INV_X4 \sha1_round/add_79_4/U348  ( .A(rnd_q[134]), .ZN(
        \sha1_round/add_79_4/n322 ) );
  XNOR2_X2 \sha1_round/add_79_4/U347  ( .A(\sha1_round/add_79_4/n319 ), .B(
        \sha1_round/add_79_4/n320 ), .ZN(sha1_round_wire[139]) );
  NAND2_X2 \sha1_round/add_79_4/U346  ( .A1(\sha1_round/add_79_4/n312 ), .A2(
        \sha1_round/add_79_4/n55 ), .ZN(\sha1_round/add_79_4/n310 ) );
  INV_X4 \sha1_round/add_79_4/U345  ( .A(\sha1_round/add_79_4/n308 ), .ZN(
        \sha1_round/add_79_4/n306 ) );
  NAND2_X2 \sha1_round/add_79_4/U344  ( .A1(\sha1_round/N328 ), .A2(rnd_q[135]), .ZN(\sha1_round/add_79_4/n296 ) );
  INV_X4 \sha1_round/add_79_4/U343  ( .A(\sha1_round/add_79_4/n296 ), .ZN(
        \sha1_round/add_79_4/n275 ) );
  XNOR2_X2 \sha1_round/add_79_4/U342  ( .A(\sha1_round/add_79_4/n297 ), .B(
        \sha1_round/add_79_4/n301 ), .ZN(sha1_round_wire[140]) );
  NAND2_X2 \sha1_round/add_79_4/U341  ( .A1(\sha1_round/N329 ), .A2(rnd_q[136]), .ZN(\sha1_round/add_79_4/n271 ) );
  XNOR2_X2 \sha1_round/add_79_4/U340  ( .A(\sha1_round/add_79_4/n299 ), .B(
        \sha1_round/add_79_4/n45 ), .ZN(sha1_round_wire[141]) );
  INV_X4 \sha1_round/add_79_4/U339  ( .A(\sha1_round/add_79_4/n298 ), .ZN(
        \sha1_round/add_79_4/n278 ) );
  INV_X4 \sha1_round/add_79_4/U338  ( .A(rnd_q[138]), .ZN(
        \sha1_round/add_79_4/n289 ) );
  INV_X4 \sha1_round/add_79_4/U337  ( .A(\sha1_round/add_79_4/n233 ), .ZN(
        \sha1_round/add_79_4/n269 ) );
  XNOR2_X2 \sha1_round/add_79_4/U336  ( .A(\sha1_round/add_79_4/n286 ), .B(
        \sha1_round/add_79_4/n287 ), .ZN(sha1_round_wire[143]) );
  NOR2_X4 \sha1_round/add_79_4/U335  ( .A1(rnd_q[139]), .A2(\sha1_round/n509 ), 
        .ZN(\sha1_round/add_79_4/n254 ) );
  INV_X4 \sha1_round/add_79_4/U334  ( .A(\sha1_round/add_79_4/n86 ), .ZN(
        \sha1_round/add_79_4/n284 ) );
  INV_X4 \sha1_round/add_79_4/U333  ( .A(\sha1_round/add_79_4/n149 ), .ZN(
        \sha1_round/add_79_4/n272 ) );
  NOR2_X4 \sha1_round/add_79_4/U332  ( .A1(\sha1_round/add_79_4/n269 ), .A2(
        \sha1_round/add_79_4/n49 ), .ZN(\sha1_round/add_79_4/n277 ) );
  INV_X4 \sha1_round/add_79_4/U331  ( .A(\sha1_round/N333 ), .ZN(
        \sha1_round/add_79_4/n263 ) );
  INV_X4 \sha1_round/add_79_4/U330  ( .A(rnd_q[140]), .ZN(
        \sha1_round/add_79_4/n264 ) );
  XNOR2_X2 \sha1_round/add_79_4/U329  ( .A(\sha1_round/add_79_4/n262 ), .B(
        \sha1_round/add_79_4/n39 ), .ZN(sha1_round_wire[145]) );
  INV_X4 \sha1_round/add_79_4/U328  ( .A(\sha1_round/add_79_4/n247 ), .ZN(
        \sha1_round/add_79_4/n257 ) );
  XNOR2_X2 \sha1_round/add_79_4/U327  ( .A(\sha1_round/add_79_4/n255 ), .B(
        \sha1_round/add_79_4/n256 ), .ZN(sha1_round_wire[146]) );
  XNOR2_X2 \sha1_round/add_79_4/U326  ( .A(\sha1_round/add_79_4/n244 ), .B(
        \sha1_round/add_79_4/n38 ), .ZN(sha1_round_wire[147]) );
  NAND2_X2 \sha1_round/add_79_4/U325  ( .A1(\sha1_round/N317 ), .A2(rnd_q[156]), .ZN(\sha1_round/add_79_4/n139 ) );
  INV_X4 \sha1_round/add_79_4/U324  ( .A(\sha1_round/add_79_4/n139 ), .ZN(
        \sha1_round/add_79_4/n242 ) );
  XNOR2_X2 \sha1_round/add_79_4/U323  ( .A(\sha1_round/add_79_4/n243 ), .B(
        \sha1_round/add_79_4/n241 ), .ZN(sha1_round_wire[129]) );
  NOR2_X4 \sha1_round/add_79_4/U322  ( .A1(\sha1_round/add_79_4/n231 ), .A2(
        \sha1_round/add_79_4/n232 ), .ZN(\sha1_round/add_79_4/n216 ) );
  INV_X4 \sha1_round/add_79_4/U321  ( .A(\sha1_round/N337 ), .ZN(
        \sha1_round/add_79_4/n227 ) );
  INV_X4 \sha1_round/add_79_4/U320  ( .A(rnd_q[144]), .ZN(
        \sha1_round/add_79_4/n228 ) );
  XNOR2_X2 \sha1_round/add_79_4/U319  ( .A(\sha1_round/add_79_4/n226 ), .B(
        \sha1_round/add_79_4/n40 ), .ZN(sha1_round_wire[149]) );
  NAND2_X2 \sha1_round/add_79_4/U318  ( .A1(rnd_q[143]), .A2(\sha1_round/N336 ), .ZN(\sha1_round/add_79_4/n224 ) );
  NAND2_X2 \sha1_round/add_79_4/U317  ( .A1(\sha1_round/add_79_4/n220 ), .A2(
        \sha1_round/add_79_4/n204 ), .ZN(\sha1_round/add_79_4/n223 ) );
  NAND2_X2 \sha1_round/add_79_4/U316  ( .A1(\sha1_round/N338 ), .A2(rnd_q[145]), .ZN(\sha1_round/add_79_4/n201 ) );
  XNOR2_X2 \sha1_round/add_79_4/U315  ( .A(\sha1_round/add_79_4/n221 ), .B(
        \sha1_round/add_79_4/n46 ), .ZN(sha1_round_wire[150]) );
  NAND2_X2 \sha1_round/add_79_4/U314  ( .A1(\sha1_round/add_79_4/n223 ), .A2(
        \sha1_round/add_79_4/n203 ), .ZN(\sha1_round/add_79_4/n215 ) );
  NAND2_X2 \sha1_round/add_79_4/U313  ( .A1(\sha1_round/add_79_4/n217 ), .A2(
        \sha1_round/add_79_4/n203 ), .ZN(\sha1_round/add_79_4/n212 ) );
  NAND2_X2 \sha1_round/add_79_4/U312  ( .A1(\sha1_round/N339 ), .A2(rnd_q[146]), .ZN(\sha1_round/add_79_4/n155 ) );
  NAND2_X2 \sha1_round/add_79_4/U311  ( .A1(\sha1_round/add_79_4/n155 ), .A2(
        \sha1_round/add_79_4/n154 ), .ZN(\sha1_round/add_79_4/n214 ) );
  INV_X4 \sha1_round/add_79_4/U310  ( .A(\sha1_round/add_79_4/n212 ), .ZN(
        \sha1_round/add_79_4/n211 ) );
  NAND3_X2 \sha1_round/add_79_4/U309  ( .A1(\sha1_round/add_79_4/n209 ), .A2(
        \sha1_round/add_79_4/n210 ), .A3(\sha1_round/add_79_4/n136 ), .ZN(
        \sha1_round/add_79_4/n206 ) );
  NAND2_X2 \sha1_round/add_79_4/U308  ( .A1(\sha1_round/add_79_4/n220 ), .A2(
        \sha1_round/add_79_4/n204 ), .ZN(\sha1_round/add_79_4/n202 ) );
  NAND2_X2 \sha1_round/add_79_4/U307  ( .A1(\sha1_round/add_79_4/n202 ), .A2(
        \sha1_round/add_79_4/n203 ), .ZN(\sha1_round/add_79_4/n200 ) );
  NAND2_X2 \sha1_round/add_79_4/U306  ( .A1(\sha1_round/add_79_4/n199 ), .A2(
        \sha1_round/add_79_4/n155 ), .ZN(\sha1_round/add_79_4/n198 ) );
  NAND2_X2 \sha1_round/add_79_4/U305  ( .A1(\sha1_round/add_79_4/n149 ), .A2(
        \sha1_round/add_79_4/n196 ), .ZN(\sha1_round/add_79_4/n195 ) );
  NAND2_X2 \sha1_round/add_79_4/U304  ( .A1(\sha1_round/N340 ), .A2(rnd_q[147]), .ZN(\sha1_round/add_79_4/n185 ) );
  INV_X4 \sha1_round/add_79_4/U303  ( .A(rnd_q[147]), .ZN(
        \sha1_round/add_79_4/n193 ) );
  NAND2_X2 \sha1_round/add_79_4/U302  ( .A1(\sha1_round/add_79_4/n185 ), .A2(
        \sha1_round/add_79_4/n178 ), .ZN(\sha1_round/add_79_4/n191 ) );
  NAND2_X2 \sha1_round/add_79_4/U301  ( .A1(\sha1_round/add_79_4/n190 ), .A2(
        \sha1_round/add_79_4/n185 ), .ZN(\sha1_round/add_79_4/n186 ) );
  INV_X4 \sha1_round/add_79_4/U300  ( .A(\sha1_round/N341 ), .ZN(
        \sha1_round/add_79_4/n188 ) );
  INV_X4 \sha1_round/add_79_4/U299  ( .A(rnd_q[148]), .ZN(
        \sha1_round/add_79_4/n189 ) );
  XNOR2_X2 \sha1_round/add_79_4/U298  ( .A(\sha1_round/add_79_4/n186 ), .B(
        \sha1_round/add_79_4/n187 ), .ZN(sha1_round_wire[153]) );
  NAND2_X2 \sha1_round/add_79_4/U297  ( .A1(\sha1_round/add_79_4/n184 ), .A2(
        \sha1_round/add_79_4/n185 ), .ZN(\sha1_round/add_79_4/n183 ) );
  NAND2_X2 \sha1_round/add_79_4/U296  ( .A1(\sha1_round/add_79_4/n174 ), .A2(
        \sha1_round/add_79_4/n172 ), .ZN(\sha1_round/add_79_4/n181 ) );
  XNOR2_X2 \sha1_round/add_79_4/U295  ( .A(\sha1_round/add_79_4/n180 ), .B(
        \sha1_round/add_79_4/n181 ), .ZN(sha1_round_wire[154]) );
  INV_X4 \sha1_round/add_79_4/U294  ( .A(\sha1_round/add_79_4/n179 ), .ZN(
        \sha1_round/add_79_4/n175 ) );
  INV_X4 \sha1_round/add_79_4/U293  ( .A(\sha1_round/add_79_4/n178 ), .ZN(
        \sha1_round/add_79_4/n177 ) );
  NOR3_X4 \sha1_round/add_79_4/U292  ( .A1(\sha1_round/add_79_4/n175 ), .A2(
        \sha1_round/add_79_4/n176 ), .A3(\sha1_round/add_79_4/n177 ), .ZN(
        \sha1_round/add_79_4/n156 ) );
  NAND2_X2 \sha1_round/add_79_4/U291  ( .A1(\sha1_round/add_79_4/n173 ), .A2(
        \sha1_round/add_79_4/n174 ), .ZN(\sha1_round/add_79_4/n171 ) );
  INV_X4 \sha1_round/add_79_4/U290  ( .A(rnd_q[150]), .ZN(
        \sha1_round/add_79_4/n169 ) );
  XNOR2_X2 \sha1_round/add_79_4/U289  ( .A(\sha1_round/add_79_4/n166 ), .B(
        \sha1_round/add_79_4/n167 ), .ZN(sha1_round_wire[155]) );
  XNOR2_X2 \sha1_round/add_79_4/U288  ( .A(\sha1_round/add_79_4/n159 ), .B(
        \sha1_round/add_79_4/n160 ), .ZN(sha1_round_wire[156]) );
  NOR3_X4 \sha1_round/add_79_4/U287  ( .A1(\sha1_round/add_79_4/n272 ), .A2(
        \sha1_round/add_79_4/n147 ), .A3(\sha1_round/add_79_4/n148 ), .ZN(
        \sha1_round/add_79_4/n99 ) );
  NAND2_X2 \sha1_round/add_79_4/U286  ( .A1(\sha1_round/add_79_4/n42 ), .A2(
        \sha1_round/add_79_4/n139 ), .ZN(\sha1_round/add_79_4/n89 ) );
  NAND2_X2 \sha1_round/add_79_4/U285  ( .A1(\sha1_round/add_79_4/n90 ), .A2(
        \sha1_round/add_79_4/n87 ), .ZN(\sha1_round/add_79_4/n138 ) );
  XNOR2_X2 \sha1_round/add_79_4/U284  ( .A(\sha1_round/add_79_4/n89 ), .B(
        \sha1_round/add_79_4/n138 ), .ZN(sha1_round_wire[130]) );
  INV_X4 \sha1_round/add_79_4/U283  ( .A(\sha1_round/add_79_4/n131 ), .ZN(
        \sha1_round/add_79_4/n129 ) );
  INV_X4 \sha1_round/add_79_4/U282  ( .A(\sha1_round/add_79_4/n106 ), .ZN(
        \sha1_round/add_79_4/n128 ) );
  INV_X4 \sha1_round/add_79_4/U281  ( .A(\sha1_round/add_79_4/n105 ), .ZN(
        \sha1_round/add_79_4/n126 ) );
  NAND3_X2 \sha1_round/add_79_4/U280  ( .A1(\sha1_round/add_79_4/n123 ), .A2(
        \sha1_round/add_79_4/n124 ), .A3(\sha1_round/add_79_4/n125 ), .ZN(
        \sha1_round/add_79_4/n122 ) );
  INV_X4 \sha1_round/add_79_4/U279  ( .A(\sha1_round/add_79_4/n116 ), .ZN(
        \sha1_round/add_79_4/n120 ) );
  XNOR2_X2 \sha1_round/add_79_4/U278  ( .A(\sha1_round/add_79_4/n118 ), .B(
        \sha1_round/add_79_4/n119 ), .ZN(sha1_round_wire[158]) );
  NAND2_X2 \sha1_round/add_79_4/U277  ( .A1(\sha1_round/add_79_4/n116 ), .A2(
        \sha1_round/add_79_4/n117 ), .ZN(\sha1_round/add_79_4/n114 ) );
  NAND2_X2 \sha1_round/add_79_4/U276  ( .A1(\sha1_round/add_79_4/n108 ), .A2(
        \sha1_round/add_79_4/n109 ), .ZN(\sha1_round/add_79_4/n102 ) );
  INV_X4 \sha1_round/add_79_4/U275  ( .A(\sha1_round/add_79_4/n99 ), .ZN(
        \sha1_round/add_79_4/n98 ) );
  XNOR2_X2 \sha1_round/add_79_4/U274  ( .A(rnd_q[154]), .B(\sha1_round/N347 ), 
        .ZN(\sha1_round/add_79_4/n92 ) );
  NAND2_X2 \sha1_round/add_79_4/U273  ( .A1(\sha1_round/add_79_4/n89 ), .A2(
        \sha1_round/add_79_4/n90 ), .ZN(\sha1_round/add_79_4/n88 ) );
  NAND2_X2 \sha1_round/add_79_4/U272  ( .A1(\sha1_round/add_79_4/n87 ), .A2(
        \sha1_round/add_79_4/n88 ), .ZN(\sha1_round/add_79_4/n83 ) );
  NAND2_X2 \sha1_round/add_79_4/U271  ( .A1(\sha1_round/add_79_4/n85 ), .A2(
        \sha1_round/add_79_4/n86 ), .ZN(\sha1_round/add_79_4/n84 ) );
  XNOR2_X2 \sha1_round/add_79_4/U270  ( .A(\sha1_round/add_79_4/n83 ), .B(
        \sha1_round/add_79_4/n84 ), .ZN(sha1_round_wire[131]) );
  NAND2_X2 \sha1_round/add_79_4/U269  ( .A1(\sha1_round/N320 ), .A2(rnd_q[159]), .ZN(\sha1_round/add_79_4/n79 ) );
  NAND2_X2 \sha1_round/add_79_4/U268  ( .A1(\sha1_round/add_79_4/n337 ), .A2(
        \sha1_round/add_79_4/n79 ), .ZN(\sha1_round/add_79_4/n82 ) );
  XNOR2_X2 \sha1_round/add_79_4/U267  ( .A(\sha1_round/add_79_4/n82 ), .B(
        \sha1_round/add_79_4/n81 ), .ZN(sha1_round_wire[132]) );
  INV_X4 \sha1_round/add_79_4/U266  ( .A(\sha1_round/add_79_4/n81 ), .ZN(
        \sha1_round/add_79_4/n63 ) );
  NAND2_X2 \sha1_round/add_79_4/U265  ( .A1(\sha1_round/N321 ), .A2(rnd_q[128]), .ZN(\sha1_round/add_79_4/n74 ) );
  INV_X4 \sha1_round/add_79_4/U264  ( .A(\sha1_round/add_79_4/n74 ), .ZN(
        \sha1_round/add_79_4/n78 ) );
  XNOR2_X2 \sha1_round/add_79_4/U263  ( .A(\sha1_round/add_79_4/n76 ), .B(
        \sha1_round/add_79_4/n77 ), .ZN(sha1_round_wire[133]) );
  NAND2_X2 \sha1_round/add_79_4/U262  ( .A1(\sha1_round/add_79_4/n72 ), .A2(
        \sha1_round/add_79_4/n70 ), .ZN(\sha1_round/add_79_4/n73 ) );
  NAND2_X2 \sha1_round/add_79_4/U261  ( .A1(\sha1_round/add_79_4/n41 ), .A2(
        \sha1_round/add_79_4/n74 ), .ZN(\sha1_round/add_79_4/n71 ) );
  XNOR2_X2 \sha1_round/add_79_4/U260  ( .A(\sha1_round/add_79_4/n73 ), .B(
        \sha1_round/add_79_4/n71 ), .ZN(sha1_round_wire[134]) );
  NAND2_X2 \sha1_round/add_79_4/U259  ( .A1(\sha1_round/add_79_4/n71 ), .A2(
        \sha1_round/add_79_4/n72 ), .ZN(\sha1_round/add_79_4/n69 ) );
  NAND2_X2 \sha1_round/add_79_4/U258  ( .A1(\sha1_round/add_79_4/n69 ), .A2(
        \sha1_round/add_79_4/n70 ), .ZN(\sha1_round/add_79_4/n65 ) );
  NAND2_X2 \sha1_round/add_79_4/U257  ( .A1(\sha1_round/add_79_4/n67 ), .A2(
        \sha1_round/add_79_4/n68 ), .ZN(\sha1_round/add_79_4/n66 ) );
  XNOR2_X2 \sha1_round/add_79_4/U256  ( .A(\sha1_round/add_79_4/n65 ), .B(
        \sha1_round/add_79_4/n66 ), .ZN(sha1_round_wire[135]) );
  INV_X4 \sha1_round/add_79_4/U255  ( .A(\sha1_round/add_79_4/n312 ), .ZN(
        \sha1_round/add_79_4/n59 ) );
  XNOR2_X2 \sha1_round/add_79_4/U254  ( .A(\sha1_round/add_79_4/n57 ), .B(
        \sha1_round/add_79_4/n58 ), .ZN(sha1_round_wire[136]) );
  NAND2_X2 \sha1_round/add_79_4/U253  ( .A1(\sha1_round/add_79_4/n55 ), .A2(
        \sha1_round/add_79_4/n311 ), .ZN(\sha1_round/add_79_4/n53 ) );
  XNOR2_X2 \sha1_round/add_79_4/U252  ( .A(\sha1_round/add_79_4/n53 ), .B(
        \sha1_round/add_79_4/n54 ), .ZN(sha1_round_wire[137]) );
  NAND2_X4 \sha1_round/add_79_4/U251  ( .A1(\sha1_round/add_79_4/n251 ), .A2(
        \sha1_round/add_79_4/n252 ), .ZN(\sha1_round/add_79_4/n236 ) );
  NAND2_X1 \sha1_round/add_79_4/U250  ( .A1(\sha1_round/N333 ), .A2(rnd_q[140]), .ZN(\sha1_round/add_79_4/n260 ) );
  NOR2_X1 \sha1_round/add_79_4/U249  ( .A1(\sha1_round/add_79_4/n250 ), .A2(
        \sha1_round/add_79_4/n236 ), .ZN(\sha1_round/add_79_4/n245 ) );
  NAND2_X4 \sha1_round/add_79_4/U248  ( .A1(\sha1_round/add_79_4/n263 ), .A2(
        \sha1_round/add_79_4/n264 ), .ZN(\sha1_round/add_79_4/n252 ) );
  NAND2_X4 \sha1_round/add_79_4/U247  ( .A1(\sha1_round/add_79_4/n163 ), .A2(
        \sha1_round/add_79_4/n164 ), .ZN(\sha1_round/add_79_4/n111 ) );
  NAND3_X4 \sha1_round/add_79_4/U246  ( .A1(\sha1_round/add_79_4/n252 ), .A2(
        \sha1_round/n509 ), .A3(rnd_q[139]), .ZN(\sha1_round/add_79_4/n259 )
         );
  NOR3_X2 \sha1_round/add_79_4/U245  ( .A1(\sha1_round/add_79_4/n147 ), .A2(
        \sha1_round/add_79_4/n148 ), .A3(\sha1_round/add_79_4/n100 ), .ZN(
        \sha1_round/add_79_4/n196 ) );
  NOR3_X2 \sha1_round/add_79_4/U244  ( .A1(\sha1_round/add_79_4/n272 ), .A2(
        \sha1_round/add_79_4/n240 ), .A3(\sha1_round/add_79_4/n148 ), .ZN(
        \sha1_round/add_79_4/n267 ) );
  NAND2_X1 \sha1_round/add_79_4/U243  ( .A1(\sha1_round/add_79_4/n307 ), .A2(
        \sha1_round/add_79_4/n303 ), .ZN(\sha1_round/add_79_4/n320 ) );
  NAND2_X4 \sha1_round/add_79_4/U242  ( .A1(\sha1_round/add_79_4/n194 ), .A2(
        \sha1_round/add_79_4/n195 ), .ZN(\sha1_round/add_79_4/n165 ) );
  NAND2_X1 \sha1_round/add_79_4/U241  ( .A1(\sha1_round/N343 ), .A2(rnd_q[150]), .ZN(\sha1_round/add_79_4/n164 ) );
  NAND2_X4 \sha1_round/add_79_4/U240  ( .A1(\sha1_round/add_79_4/n168 ), .A2(
        \sha1_round/add_79_4/n169 ), .ZN(\sha1_round/add_79_4/n157 ) );
  NAND2_X1 \sha1_round/add_79_4/U239  ( .A1(\sha1_round/add_79_4/n164 ), .A2(
        \sha1_round/add_79_4/n157 ), .ZN(\sha1_round/add_79_4/n167 ) );
  NAND2_X1 \sha1_round/add_79_4/U238  ( .A1(\sha1_round/N346 ), .A2(rnd_q[153]), .ZN(\sha1_round/add_79_4/n116 ) );
  NAND2_X1 \sha1_round/add_79_4/U237  ( .A1(\sha1_round/N344 ), .A2(rnd_q[151]), .ZN(\sha1_round/add_79_4/n131 ) );
  NAND2_X1 \sha1_round/add_79_4/U236  ( .A1(rnd_q[144]), .A2(\sha1_round/N337 ), .ZN(\sha1_round/add_79_4/n204 ) );
  INV_X1 \sha1_round/add_79_4/U235  ( .A(\sha1_round/add_79_4/n252 ), .ZN(
        \sha1_round/add_79_4/n261 ) );
  NAND2_X1 \sha1_round/add_79_4/U234  ( .A1(\sha1_round/add_79_4/n117 ), .A2(
        \sha1_round/add_79_4/n127 ), .ZN(\sha1_round/add_79_4/n142 ) );
  NAND2_X1 \sha1_round/add_79_4/U233  ( .A1(\sha1_round/add_79_4/n136 ), .A2(
        \sha1_round/add_79_4/n127 ), .ZN(\sha1_round/add_79_4/n135 ) );
  NAND2_X1 \sha1_round/add_79_4/U232  ( .A1(\sha1_round/N334 ), .A2(rnd_q[141]), .ZN(\sha1_round/add_79_4/n247 ) );
  NAND2_X1 \sha1_round/add_79_4/U231  ( .A1(\sha1_round/add_79_4/n131 ), .A2(
        \sha1_round/add_79_4/n158 ), .ZN(\sha1_round/add_79_4/n160 ) );
  NAND2_X4 \sha1_round/add_79_4/U230  ( .A1(\sha1_round/add_79_4/n188 ), .A2(
        \sha1_round/add_79_4/n189 ), .ZN(\sha1_round/add_79_4/n179 ) );
  NAND2_X1 \sha1_round/add_79_4/U229  ( .A1(\sha1_round/add_79_4/n179 ), .A2(
        \sha1_round/add_79_4/n184 ), .ZN(\sha1_round/add_79_4/n187 ) );
  NOR2_X1 \sha1_round/add_79_4/U228  ( .A1(\sha1_round/add_79_4/n254 ), .A2(
        \sha1_round/add_79_4/n52 ), .ZN(\sha1_round/add_79_4/n266 ) );
  NOR2_X1 \sha1_round/add_79_4/U227  ( .A1(\sha1_round/add_79_4/n254 ), .A2(
        \sha1_round/add_79_4/n250 ), .ZN(\sha1_round/add_79_4/n265 ) );
  NOR3_X1 \sha1_round/add_79_4/U226  ( .A1(\sha1_round/add_79_4/n250 ), .A2(
        \sha1_round/add_79_4/n261 ), .A3(\sha1_round/add_79_4/n254 ), .ZN(
        \sha1_round/add_79_4/n258 ) );
  NAND3_X2 \sha1_round/add_79_4/U225  ( .A1(\sha1_round/add_79_4/n95 ), .A2(
        \sha1_round/add_79_4/n146 ), .A3(\sha1_round/add_79_4/n145 ), .ZN(
        \sha1_round/add_79_4/n94 ) );
  INV_X4 \sha1_round/add_79_4/U224  ( .A(\sha1_round/add_79_4/n273 ), .ZN(
        \sha1_round/add_79_4/n281 ) );
  NAND2_X2 \sha1_round/add_79_4/U223  ( .A1(\sha1_round/add_79_4/n86 ), .A2(
        \sha1_round/add_79_4/n331 ), .ZN(\sha1_round/add_79_4/n81 ) );
  AND2_X2 \sha1_round/add_79_4/U222  ( .A1(\sha1_round/n509 ), .A2(rnd_q[139]), 
        .ZN(\sha1_round/add_79_4/n52 ) );
  AND2_X2 \sha1_round/add_79_4/U221  ( .A1(\sha1_round/N336 ), .A2(rnd_q[143]), 
        .ZN(\sha1_round/add_79_4/n51 ) );
  NOR2_X2 \sha1_round/add_79_4/U220  ( .A1(\sha1_round/add_79_4/n344 ), .A2(
        \sha1_round/add_79_4/n345 ), .ZN(\sha1_round/add_79_4/n343 ) );
  NAND3_X1 \sha1_round/add_79_4/U219  ( .A1(rnd_q[128]), .A2(\sha1_round/N321 ), .A3(\sha1_round/add_79_4/n72 ), .ZN(\sha1_round/add_79_4/n342 ) );
  NAND3_X2 \sha1_round/add_79_4/U218  ( .A1(\sha1_round/add_79_4/n341 ), .A2(
        \sha1_round/add_79_4/n342 ), .A3(\sha1_round/add_79_4/n343 ), .ZN(
        \sha1_round/add_79_4/n316 ) );
  OR2_X2 \sha1_round/add_79_4/U217  ( .A1(rnd_q[155]), .A2(\sha1_round/N316 ), 
        .ZN(\sha1_round/add_79_4/n50 ) );
  OR2_X2 \sha1_round/add_79_4/U216  ( .A1(\sha1_round/N318 ), .A2(rnd_q[157]), 
        .ZN(\sha1_round/add_79_4/n90 ) );
  NOR2_X2 \sha1_round/add_79_4/U215  ( .A1(rnd_q[159]), .A2(\sha1_round/N320 ), 
        .ZN(\sha1_round/add_79_4/n80 ) );
  NOR2_X2 \sha1_round/add_79_4/U214  ( .A1(rnd_q[156]), .A2(\sha1_round/N317 ), 
        .ZN(\sha1_round/add_79_4/n140 ) );
  NOR2_X2 \sha1_round/add_79_4/U213  ( .A1(rnd_q[128]), .A2(\sha1_round/N321 ), 
        .ZN(\sha1_round/add_79_4/n75 ) );
  OR2_X2 \sha1_round/add_79_4/U212  ( .A1(\sha1_round/N319 ), .A2(rnd_q[158]), 
        .ZN(\sha1_round/add_79_4/n85 ) );
  AND2_X2 \sha1_round/add_79_4/U211  ( .A1(\sha1_round/add_79_4/n203 ), .A2(
        \sha1_round/add_79_4/n201 ), .ZN(\sha1_round/add_79_4/n46 ) );
  AND2_X2 \sha1_round/add_79_4/U210  ( .A1(\sha1_round/add_79_4/n271 ), .A2(
        \sha1_round/add_79_4/n298 ), .ZN(\sha1_round/add_79_4/n45 ) );
  NOR2_X1 \sha1_round/add_79_4/U209  ( .A1(\sha1_round/add_79_4/n112 ), .A2(
        \sha1_round/add_79_4/n120 ), .ZN(\sha1_round/add_79_4/n119 ) );
  NOR2_X1 \sha1_round/add_79_4/U208  ( .A1(\sha1_round/add_79_4/n269 ), .A2(
        \sha1_round/add_79_4/n5 ), .ZN(\sha1_round/add_79_4/n287 ) );
  NOR2_X1 \sha1_round/add_79_4/U207  ( .A1(\sha1_round/add_79_4/n3 ), .A2(
        \sha1_round/add_79_4/n49 ), .ZN(\sha1_round/add_79_4/n292 ) );
  NOR2_X1 \sha1_round/add_79_4/U206  ( .A1(\sha1_round/add_79_4/n48 ), .A2(
        \sha1_round/add_79_4/n297 ), .ZN(\sha1_round/add_79_4/n300 ) );
  NOR2_X2 \sha1_round/add_79_4/U205  ( .A1(\sha1_round/add_79_4/n275 ), .A2(
        \sha1_round/add_79_4/n300 ), .ZN(\sha1_round/add_79_4/n299 ) );
  NOR2_X1 \sha1_round/add_79_4/U204  ( .A1(\sha1_round/add_79_4/n275 ), .A2(
        \sha1_round/add_79_4/n48 ), .ZN(\sha1_round/add_79_4/n301 ) );
  NOR2_X2 \sha1_round/add_79_4/U203  ( .A1(\sha1_round/add_79_4/n59 ), .A2(
        \sha1_round/add_79_4/n60 ), .ZN(\sha1_round/add_79_4/n58 ) );
  NOR2_X2 \sha1_round/add_79_4/U202  ( .A1(\sha1_round/add_79_4/n265 ), .A2(
        \sha1_round/add_79_4/n52 ), .ZN(\sha1_round/add_79_4/n262 ) );
  NOR2_X1 \sha1_round/add_79_4/U201  ( .A1(\sha1_round/add_79_4/n218 ), .A2(
        \sha1_round/add_79_4/n51 ), .ZN(\sha1_round/add_79_4/n230 ) );
  NOR2_X2 \sha1_round/add_79_4/U200  ( .A1(\sha1_round/add_79_4/n242 ), .A2(
        \sha1_round/add_79_4/n140 ), .ZN(\sha1_round/add_79_4/n241 ) );
  NOR2_X2 \sha1_round/add_79_4/U199  ( .A1(\sha1_round/add_79_4/n335 ), .A2(
        \sha1_round/add_79_4/n140 ), .ZN(\sha1_round/add_79_4/n334 ) );
  NAND3_X1 \sha1_round/add_79_4/U198  ( .A1(\sha1_round/add_79_4/n318 ), .A2(
        \sha1_round/add_79_4/n314 ), .A3(\sha1_round/add_79_4/n81 ), .ZN(
        \sha1_round/add_79_4/n330 ) );
  NAND3_X2 \sha1_round/add_79_4/U197  ( .A1(\sha1_round/add_79_4/n312 ), .A2(
        \sha1_round/add_79_4/n329 ), .A3(\sha1_round/add_79_4/n330 ), .ZN(
        \sha1_round/add_79_4/n54 ) );
  NOR2_X1 \sha1_round/add_79_4/U196  ( .A1(\sha1_round/add_79_4/n253 ), .A2(
        \sha1_round/add_79_4/n257 ), .ZN(\sha1_round/add_79_4/n256 ) );
  NOR3_X2 \sha1_round/add_79_4/U195  ( .A1(\sha1_round/add_79_4/n7 ), .A2(
        \sha1_round/add_79_4/n284 ), .A3(\sha1_round/add_79_4/n285 ), .ZN(
        \sha1_round/add_79_4/n283 ) );
  AND2_X2 \sha1_round/add_79_4/U194  ( .A1(\sha1_round/add_79_4/n43 ), .A2(
        \sha1_round/add_79_4/n79 ), .ZN(\sha1_round/add_79_4/n76 ) );
  OR2_X2 \sha1_round/add_79_4/U193  ( .A1(\sha1_round/add_79_4/n140 ), .A2(
        \sha1_round/add_79_4/n243 ), .ZN(\sha1_round/add_79_4/n42 ) );
  NOR2_X2 \sha1_round/add_79_4/U192  ( .A1(\sha1_round/add_79_4/n332 ), .A2(
        \sha1_round/add_79_4/n87 ), .ZN(\sha1_round/add_79_4/n285 ) );
  NOR2_X1 \sha1_round/add_79_4/U191  ( .A1(\sha1_round/add_79_4/n278 ), .A2(
        \sha1_round/add_79_4/n296 ), .ZN(\sha1_round/add_79_4/n295 ) );
  AND2_X2 \sha1_round/add_79_4/U190  ( .A1(\sha1_round/add_79_4/n204 ), .A2(
        \sha1_round/add_79_4/n225 ), .ZN(\sha1_round/add_79_4/n40 ) );
  AND2_X2 \sha1_round/add_79_4/U189  ( .A1(\sha1_round/add_79_4/n260 ), .A2(
        \sha1_round/add_79_4/n252 ), .ZN(\sha1_round/add_79_4/n39 ) );
  AND2_X2 \sha1_round/add_79_4/U188  ( .A1(\sha1_round/add_79_4/n150 ), .A2(
        \sha1_round/add_79_4/n210 ), .ZN(\sha1_round/add_79_4/n38 ) );
  NOR2_X2 \sha1_round/add_79_4/U187  ( .A1(\sha1_round/add_79_4/n49 ), .A2(
        \sha1_round/add_79_4/n271 ), .ZN(\sha1_round/add_79_4/n270 ) );
  NOR2_X2 \sha1_round/add_79_4/U186  ( .A1(\sha1_round/add_79_4/n7 ), .A2(
        \sha1_round/add_79_4/n285 ), .ZN(\sha1_round/add_79_4/n331 ) );
  NOR2_X1 \sha1_round/add_79_4/U185  ( .A1(\sha1_round/add_79_4/n61 ), .A2(
        \sha1_round/add_79_4/n62 ), .ZN(\sha1_round/add_79_4/n57 ) );
  NOR2_X2 \sha1_round/add_79_4/U184  ( .A1(\sha1_round/add_79_4/n27 ), .A2(
        \sha1_round/add_79_4/n151 ), .ZN(\sha1_round/add_79_4/n143 ) );
  NOR2_X1 \sha1_round/add_79_4/U183  ( .A1(\sha1_round/add_79_4/n269 ), .A2(
        \sha1_round/add_79_4/n235 ), .ZN(\sha1_round/add_79_4/n268 ) );
  OR2_X4 \sha1_round/add_79_4/U182  ( .A1(\sha1_round/N329 ), .A2(rnd_q[136]), 
        .ZN(\sha1_round/add_79_4/n298 ) );
  OR2_X4 \sha1_round/add_79_4/U181  ( .A1(\sha1_round/N345 ), .A2(rnd_q[152]), 
        .ZN(\sha1_round/add_79_4/n127 ) );
  OR2_X4 \sha1_round/add_79_4/U180  ( .A1(\sha1_round/N322 ), .A2(rnd_q[129]), 
        .ZN(\sha1_round/add_79_4/n72 ) );
  OR2_X1 \sha1_round/add_79_4/U179  ( .A1(\sha1_round/add_79_4/n63 ), .A2(
        \sha1_round/add_79_4/n80 ), .ZN(\sha1_round/add_79_4/n43 ) );
  NOR2_X1 \sha1_round/add_79_4/U178  ( .A1(\sha1_round/add_79_4/n78 ), .A2(
        \sha1_round/add_79_4/n75 ), .ZN(\sha1_round/add_79_4/n77 ) );
  OR2_X4 \sha1_round/add_79_4/U177  ( .A1(\sha1_round/add_79_4/n75 ), .A2(
        \sha1_round/add_79_4/n76 ), .ZN(\sha1_round/add_79_4/n41 ) );
  AND2_X2 \sha1_round/add_79_4/U176  ( .A1(\sha1_round/add_79_4/n302 ), .A2(
        \sha1_round/add_79_4/n281 ), .ZN(\sha1_round/add_79_4/n37 ) );
  NAND3_X4 \sha1_round/add_79_4/U175  ( .A1(\sha1_round/add_79_4/n279 ), .A2(
        \sha1_round/add_79_4/n280 ), .A3(\sha1_round/add_79_4/n281 ), .ZN(
        \sha1_round/add_79_4/n149 ) );
  NOR2_X1 \sha1_round/add_79_4/U174  ( .A1(\sha1_round/add_79_4/n63 ), .A2(
        \sha1_round/add_79_4/n64 ), .ZN(\sha1_round/add_79_4/n61 ) );
  OR2_X4 \sha1_round/add_79_4/U173  ( .A1(\sha1_round/N338 ), .A2(rnd_q[145]), 
        .ZN(\sha1_round/add_79_4/n203 ) );
  OR2_X4 \sha1_round/add_79_4/U172  ( .A1(\sha1_round/N339 ), .A2(rnd_q[146]), 
        .ZN(\sha1_round/add_79_4/n154 ) );
  NOR2_X2 \sha1_round/add_79_4/U171  ( .A1(\sha1_round/add_79_4/n245 ), .A2(
        \sha1_round/add_79_4/n209 ), .ZN(\sha1_round/add_79_4/n244 ) );
  AND2_X4 \sha1_round/add_79_4/U170  ( .A1(\sha1_round/add_79_4/n21 ), .A2(
        \sha1_round/add_79_4/n150 ), .ZN(\sha1_round/add_79_4/n44 ) );
  NOR2_X2 \sha1_round/add_79_4/U169  ( .A1(\sha1_round/add_79_4/n134 ), .A2(
        \sha1_round/add_79_4/n9 ), .ZN(\sha1_round/add_79_4/n121 ) );
  NOR2_X2 \sha1_round/add_79_4/U168  ( .A1(rnd_q[131]), .A2(\sha1_round/N324 ), 
        .ZN(\sha1_round/add_79_4/n60 ) );
  NAND2_X2 \sha1_round/add_79_4/U167  ( .A1(\sha1_round/add_79_4/n21 ), .A2(
        \sha1_round/add_79_4/n150 ), .ZN(\sha1_round/add_79_4/n208 ) );
  NOR2_X1 \sha1_round/add_79_4/U166  ( .A1(\sha1_round/add_79_4/n99 ), .A2(
        \sha1_round/add_79_4/n137 ), .ZN(\sha1_round/add_79_4/n134 ) );
  NAND2_X2 \sha1_round/add_79_4/U165  ( .A1(\sha1_round/add_79_4/n208 ), .A2(
        \sha1_round/add_79_4/n136 ), .ZN(\sha1_round/add_79_4/n207 ) );
  XNOR2_X1 \sha1_round/add_79_4/U164  ( .A(\sha1_round/add_79_4/n291 ), .B(
        \sha1_round/add_79_4/n292 ), .ZN(sha1_round_wire[142]) );
  INV_X1 \sha1_round/add_79_4/U163  ( .A(\sha1_round/add_79_4/n271 ), .ZN(
        \sha1_round/add_79_4/n294 ) );
  NOR2_X4 \sha1_round/add_79_4/U162  ( .A1(\sha1_round/add_79_4/n273 ), .A2(
        \sha1_round/add_79_4/n11 ), .ZN(\sha1_round/add_79_4/n148 ) );
  NAND2_X4 \sha1_round/add_79_4/U161  ( .A1(\sha1_round/add_79_4/n156 ), .A2(
        \sha1_round/add_79_4/n110 ), .ZN(\sha1_round/add_79_4/n96 ) );
  NOR2_X4 \sha1_round/add_79_4/U160  ( .A1(\sha1_round/add_79_4/n129 ), .A2(
        \sha1_round/add_79_4/n130 ), .ZN(\sha1_round/add_79_4/n106 ) );
  NOR2_X2 \sha1_round/add_79_4/U159  ( .A1(\sha1_round/add_79_4/n106 ), .A2(
        \sha1_round/add_79_4/n107 ), .ZN(\sha1_round/add_79_4/n103 ) );
  NAND2_X4 \sha1_round/add_79_4/U158  ( .A1(\sha1_round/add_79_4/n158 ), .A2(
        \sha1_round/add_79_4/n157 ), .ZN(\sha1_round/add_79_4/n36 ) );
  INV_X4 \sha1_round/add_79_4/U157  ( .A(\sha1_round/add_79_4/n96 ), .ZN(
        \sha1_round/add_79_4/n145 ) );
  NAND2_X2 \sha1_round/add_79_4/U156  ( .A1(\sha1_round/add_79_4/n2 ), .A2(
        \sha1_round/add_79_4/n146 ), .ZN(\sha1_round/add_79_4/n144 ) );
  INV_X4 \sha1_round/add_79_4/U155  ( .A(\sha1_round/add_79_4/n92 ), .ZN(
        \sha1_round/add_79_4/n33 ) );
  NAND2_X2 \sha1_round/add_79_4/U154  ( .A1(\sha1_round/add_79_4/n91 ), .A2(
        \sha1_round/add_79_4/n92 ), .ZN(\sha1_round/add_79_4/n34 ) );
  NAND2_X2 \sha1_round/add_79_4/U153  ( .A1(\sha1_round/add_79_4/n17 ), .A2(
        \sha1_round/add_79_4/n165 ), .ZN(\sha1_round/add_79_4/n182 ) );
  NAND2_X2 \sha1_round/add_79_4/U152  ( .A1(\sha1_round/add_79_4/n156 ), .A2(
        \sha1_round/add_79_4/n165 ), .ZN(\sha1_round/add_79_4/n170 ) );
  NAND2_X2 \sha1_round/add_79_4/U151  ( .A1(\sha1_round/add_79_4/n178 ), .A2(
        \sha1_round/add_79_4/n165 ), .ZN(\sha1_round/add_79_4/n190 ) );
  NAND3_X4 \sha1_round/add_79_4/U150  ( .A1(\sha1_round/add_79_4/n215 ), .A2(
        \sha1_round/add_79_4/n201 ), .A3(\sha1_round/add_79_4/n6 ), .ZN(
        \sha1_round/add_79_4/n213 ) );
  NAND2_X2 \sha1_round/add_79_4/U149  ( .A1(\sha1_round/add_79_4/n1 ), .A2(
        \sha1_round/add_79_4/n165 ), .ZN(\sha1_round/add_79_4/n161 ) );
  NAND3_X1 \sha1_round/add_79_4/U148  ( .A1(\sha1_round/add_79_4/n68 ), .A2(
        \sha1_round/add_79_4/n316 ), .A3(\sha1_round/add_79_4/n274 ), .ZN(
        \sha1_round/add_79_4/n315 ) );
  NAND3_X1 \sha1_round/add_79_4/U147  ( .A1(\sha1_round/add_79_4/n314 ), .A2(
        \sha1_round/add_79_4/n274 ), .A3(\sha1_round/add_79_4/n81 ), .ZN(
        \sha1_round/add_79_4/n302 ) );
  NAND3_X4 \sha1_round/add_79_4/U146  ( .A1(\sha1_round/add_79_4/n153 ), .A2(
        \sha1_round/add_79_4/n145 ), .A3(\sha1_round/add_79_4/n154 ), .ZN(
        \sha1_round/add_79_4/n105 ) );
  NAND2_X2 \sha1_round/add_79_4/U145  ( .A1(\sha1_round/add_79_4/n183 ), .A2(
        \sha1_round/add_79_4/n179 ), .ZN(\sha1_round/add_79_4/n173 ) );
  INV_X1 \sha1_round/add_79_4/U144  ( .A(\sha1_round/add_79_4/n176 ), .ZN(
        \sha1_round/add_79_4/n172 ) );
  NOR2_X4 \sha1_round/add_79_4/U143  ( .A1(\sha1_round/add_79_4/n112 ), .A2(
        \sha1_round/add_79_4/n113 ), .ZN(\sha1_round/add_79_4/n101 ) );
  NAND3_X2 \sha1_round/add_79_4/U142  ( .A1(\sha1_round/add_79_4/n152 ), .A2(
        \sha1_round/add_79_4/n105 ), .A3(\sha1_round/add_79_4/n131 ), .ZN(
        \sha1_round/add_79_4/n151 ) );
  NAND2_X2 \sha1_round/add_79_4/U141  ( .A1(\sha1_round/add_79_4/n182 ), .A2(
        \sha1_round/add_79_4/n173 ), .ZN(\sha1_round/add_79_4/n180 ) );
  INV_X2 \sha1_round/add_79_4/U140  ( .A(\sha1_round/add_79_4/n253 ), .ZN(
        \sha1_round/add_79_4/n249 ) );
  NAND2_X4 \sha1_round/add_79_4/U139  ( .A1(\sha1_round/add_79_4/n128 ), .A2(
        \sha1_round/add_79_4/n127 ), .ZN(\sha1_round/add_79_4/n124 ) );
  NOR2_X4 \sha1_round/add_79_4/U138  ( .A1(rnd_q[141]), .A2(\sha1_round/N334 ), 
        .ZN(\sha1_round/add_79_4/n253 ) );
  NAND2_X4 \sha1_round/add_79_4/U137  ( .A1(\sha1_round/add_79_4/n93 ), .A2(
        \sha1_round/add_79_4/n94 ), .ZN(\sha1_round/add_79_4/n91 ) );
  NOR2_X2 \sha1_round/add_79_4/U136  ( .A1(\sha1_round/add_79_4/n107 ), .A2(
        \sha1_round/add_79_4/n100 ), .ZN(\sha1_round/add_79_4/n95 ) );
  NAND2_X2 \sha1_round/add_79_4/U135  ( .A1(\sha1_round/add_79_4/n126 ), .A2(
        \sha1_round/add_79_4/n127 ), .ZN(\sha1_round/add_79_4/n125 ) );
  AND2_X4 \sha1_round/add_79_4/U134  ( .A1(\sha1_round/add_79_4/n132 ), .A2(
        \sha1_round/add_79_4/n117 ), .ZN(\sha1_round/add_79_4/n123 ) );
  NOR2_X1 \sha1_round/add_79_4/U133  ( .A1(\sha1_round/add_79_4/n218 ), .A2(
        \sha1_round/add_79_4/n216 ), .ZN(\sha1_round/add_79_4/n229 ) );
  NAND2_X4 \sha1_round/add_79_4/U132  ( .A1(\sha1_round/add_79_4/n15 ), .A2(
        \sha1_round/add_79_4/n238 ), .ZN(\sha1_round/add_79_4/n147 ) );
  NOR2_X1 \sha1_round/add_79_4/U131  ( .A1(\sha1_round/add_79_4/n216 ), .A2(
        \sha1_round/add_79_4/n14 ), .ZN(\sha1_round/add_79_4/n222 ) );
  INV_X4 \sha1_round/add_79_4/U130  ( .A(\sha1_round/add_79_4/n214 ), .ZN(
        \sha1_round/add_79_4/n29 ) );
  NAND2_X2 \sha1_round/add_79_4/U129  ( .A1(\sha1_round/add_79_4/n213 ), .A2(
        \sha1_round/add_79_4/n214 ), .ZN(\sha1_round/add_79_4/n30 ) );
  OR2_X4 \sha1_round/add_79_4/U128  ( .A1(\sha1_round/N323 ), .A2(rnd_q[130]), 
        .ZN(\sha1_round/add_79_4/n68 ) );
  AND2_X4 \sha1_round/add_79_4/U127  ( .A1(\sha1_round/add_79_4/n315 ), .A2(
        \sha1_round/add_79_4/n37 ), .ZN(\sha1_round/add_79_4/n297 ) );
  NAND2_X2 \sha1_round/add_79_4/U126  ( .A1(\sha1_round/add_79_4/n27 ), .A2(
        \sha1_round/add_79_4/n101 ), .ZN(\sha1_round/add_79_4/n109 ) );
  NAND2_X2 \sha1_round/add_79_4/U125  ( .A1(\sha1_round/add_79_4/n111 ), .A2(
        \sha1_round/add_79_4/n20 ), .ZN(\sha1_round/add_79_4/n26 ) );
  INV_X2 \sha1_round/add_79_4/U124  ( .A(\sha1_round/add_79_4/n142 ), .ZN(
        \sha1_round/add_79_4/n23 ) );
  INV_X4 \sha1_round/add_79_4/U123  ( .A(\sha1_round/add_79_4/n141 ), .ZN(
        \sha1_round/add_79_4/n22 ) );
  NAND2_X4 \sha1_round/add_79_4/U122  ( .A1(\sha1_round/add_79_4/n276 ), .A2(
        \sha1_round/add_79_4/n277 ), .ZN(\sha1_round/add_79_4/n240 ) );
  NAND2_X2 \sha1_round/add_79_4/U121  ( .A1(\sha1_round/add_79_4/n133 ), .A2(
        \sha1_round/add_79_4/n111 ), .ZN(\sha1_round/add_79_4/n132 ) );
  NOR2_X4 \sha1_round/add_79_4/U120  ( .A1(\sha1_round/add_79_4/n235 ), .A2(
        \sha1_round/add_79_4/n236 ), .ZN(\sha1_round/add_79_4/n234 ) );
  NAND2_X4 \sha1_round/add_79_4/U119  ( .A1(\sha1_round/add_79_4/n4 ), .A2(
        \sha1_round/add_79_4/n234 ), .ZN(\sha1_round/add_79_4/n21 ) );
  NOR3_X4 \sha1_round/add_79_4/U118  ( .A1(\sha1_round/add_79_4/n270 ), .A2(
        \sha1_round/add_79_4/n3 ), .A3(\sha1_round/add_79_4/n5 ), .ZN(
        \sha1_round/add_79_4/n235 ) );
  NAND2_X2 \sha1_round/add_79_4/U117  ( .A1(\sha1_round/add_79_4/n306 ), .A2(
        \sha1_round/add_79_4/n307 ), .ZN(\sha1_round/add_79_4/n305 ) );
  NOR2_X2 \sha1_round/add_79_4/U116  ( .A1(\sha1_round/add_79_4/n258 ), .A2(
        \sha1_round/add_79_4/n248 ), .ZN(\sha1_round/add_79_4/n255 ) );
  INV_X2 \sha1_round/add_79_4/U115  ( .A(\sha1_round/add_79_4/n149 ), .ZN(
        \sha1_round/add_79_4/n237 ) );
  NAND2_X1 \sha1_round/add_79_4/U114  ( .A1(\sha1_round/N327 ), .A2(rnd_q[134]), .ZN(\sha1_round/add_79_4/n303 ) );
  NAND3_X2 \sha1_round/add_79_4/U113  ( .A1(\sha1_round/add_79_4/n44 ), .A2(
        \sha1_round/add_79_4/n97 ), .A3(\sha1_round/add_79_4/n98 ), .ZN(
        \sha1_round/add_79_4/n146 ) );
  INV_X2 \sha1_round/add_79_4/U112  ( .A(\sha1_round/add_79_4/n19 ), .ZN(
        \sha1_round/add_79_4/n20 ) );
  INV_X1 \sha1_round/add_79_4/U111  ( .A(\sha1_round/add_79_4/n110 ), .ZN(
        \sha1_round/add_79_4/n19 ) );
  XNOR2_X1 \sha1_round/add_79_4/U110  ( .A(\sha1_round/add_79_4/n216 ), .B(
        \sha1_round/add_79_4/n230 ), .ZN(sha1_round_wire[148]) );
  NOR2_X2 \sha1_round/add_79_4/U109  ( .A1(\sha1_round/add_79_4/n283 ), .A2(
        \sha1_round/add_79_4/n64 ), .ZN(\sha1_round/add_79_4/n282 ) );
  NOR2_X4 \sha1_round/add_79_4/U108  ( .A1(\sha1_round/add_79_4/n282 ), .A2(
        \sha1_round/add_79_4/n275 ), .ZN(\sha1_round/add_79_4/n279 ) );
  INV_X4 \sha1_round/add_79_4/U107  ( .A(\sha1_round/add_79_4/n236 ), .ZN(
        \sha1_round/add_79_4/n239 ) );
  NAND2_X1 \sha1_round/add_79_4/U106  ( .A1(\sha1_round/add_79_4/n114 ), .A2(
        \sha1_round/add_79_4/n115 ), .ZN(\sha1_round/add_79_4/n108 ) );
  INV_X2 \sha1_round/add_79_4/U105  ( .A(\sha1_round/add_79_4/n47 ), .ZN(
        \sha1_round/add_79_4/n210 ) );
  INV_X2 \sha1_round/add_79_4/U104  ( .A(\sha1_round/add_79_4/n26 ), .ZN(
        \sha1_round/add_79_4/n27 ) );
  OR2_X2 \sha1_round/add_79_4/U103  ( .A1(\sha1_round/N346 ), .A2(rnd_q[153]), 
        .ZN(\sha1_round/add_79_4/n115 ) );
  INV_X4 \sha1_round/add_79_4/U102  ( .A(\sha1_round/add_79_4/n115 ), .ZN(
        \sha1_round/add_79_4/n112 ) );
  NOR2_X4 \sha1_round/add_79_4/U101  ( .A1(rnd_q[149]), .A2(\sha1_round/N342 ), 
        .ZN(\sha1_round/add_79_4/n176 ) );
  NAND2_X2 \sha1_round/add_79_4/U100  ( .A1(\sha1_round/N323 ), .A2(rnd_q[130]), .ZN(\sha1_round/add_79_4/n67 ) );
  NOR2_X2 \sha1_round/add_79_4/U99  ( .A1(\sha1_round/add_79_4/n229 ), .A2(
        \sha1_round/add_79_4/n51 ), .ZN(\sha1_round/add_79_4/n226 ) );
  NOR2_X2 \sha1_round/add_79_4/U98  ( .A1(\sha1_round/add_79_4/n197 ), .A2(
        \sha1_round/add_79_4/n198 ), .ZN(\sha1_round/add_79_4/n194 ) );
  AND2_X4 \sha1_round/add_79_4/U97  ( .A1(\sha1_round/add_79_4/n318 ), .A2(
        \sha1_round/add_79_4/n313 ), .ZN(\sha1_round/add_79_4/n18 ) );
  INV_X4 \sha1_round/add_79_4/U96  ( .A(\sha1_round/add_79_4/n205 ), .ZN(
        \sha1_round/add_79_4/n220 ) );
  AND2_X4 \sha1_round/add_79_4/U95  ( .A1(\sha1_round/add_79_4/n178 ), .A2(
        \sha1_round/add_79_4/n179 ), .ZN(\sha1_round/add_79_4/n17 ) );
  AND2_X4 \sha1_round/add_79_4/U94  ( .A1(\sha1_round/add_79_4/n243 ), .A2(
        \sha1_round/add_79_4/n50 ), .ZN(sha1_round_wire[128]) );
  NOR2_X2 \sha1_round/add_79_4/U93  ( .A1(rnd_q[132]), .A2(\sha1_round/N325 ), 
        .ZN(\sha1_round/add_79_4/n56 ) );
  AND2_X2 \sha1_round/add_79_4/U92  ( .A1(\sha1_round/add_79_4/n239 ), .A2(
        \sha1_round/add_79_4/n210 ), .ZN(\sha1_round/add_79_4/n15 ) );
  OR2_X4 \sha1_round/add_79_4/U91  ( .A1(\sha1_round/add_79_4/n219 ), .A2(
        \sha1_round/add_79_4/n218 ), .ZN(\sha1_round/add_79_4/n14 ) );
  AND2_X4 \sha1_round/add_79_4/U90  ( .A1(\sha1_round/add_79_4/n150 ), .A2(
        \sha1_round/add_79_4/n21 ), .ZN(\sha1_round/add_79_4/n13 ) );
  AND2_X4 \sha1_round/add_79_4/U89  ( .A1(\sha1_round/add_79_4/n303 ), .A2(
        \sha1_round/add_79_4/n305 ), .ZN(\sha1_round/add_79_4/n12 ) );
  OR2_X4 \sha1_round/add_79_4/U88  ( .A1(\sha1_round/add_79_4/n274 ), .A2(
        \sha1_round/add_79_4/n275 ), .ZN(\sha1_round/add_79_4/n11 ) );
  OR2_X4 \sha1_round/add_79_4/U87  ( .A1(\sha1_round/add_79_4/n295 ), .A2(
        \sha1_round/add_79_4/n294 ), .ZN(\sha1_round/add_79_4/n10 ) );
  OR2_X1 \sha1_round/add_79_4/U86  ( .A1(\sha1_round/add_79_4/n135 ), .A2(
        \sha1_round/add_79_4/n96 ), .ZN(\sha1_round/add_79_4/n9 ) );
  OR2_X4 \sha1_round/add_79_4/U85  ( .A1(\sha1_round/add_79_4/n278 ), .A2(
        \sha1_round/add_79_4/n48 ), .ZN(\sha1_round/add_79_4/n8 ) );
  AND3_X4 \sha1_round/add_79_4/U84  ( .A1(\sha1_round/add_79_4/n85 ), .A2(
        \sha1_round/add_79_4/n333 ), .A3(\sha1_round/add_79_4/n334 ), .ZN(
        \sha1_round/add_79_4/n7 ) );
  OR2_X4 \sha1_round/add_79_4/U83  ( .A1(\sha1_round/add_79_4/n216 ), .A2(
        \sha1_round/add_79_4/n212 ), .ZN(\sha1_round/add_79_4/n6 ) );
  AND2_X4 \sha1_round/add_79_4/U82  ( .A1(\sha1_round/add_79_4/n233 ), .A2(
        \sha1_round/add_79_4/n210 ), .ZN(\sha1_round/add_79_4/n4 ) );
  AND2_X4 \sha1_round/add_79_4/U81  ( .A1(\sha1_round/N330 ), .A2(rnd_q[137]), 
        .ZN(\sha1_round/add_79_4/n3 ) );
  NOR3_X4 \sha1_round/add_79_4/U80  ( .A1(\sha1_round/add_79_4/n102 ), .A2(
        \sha1_round/add_79_4/n103 ), .A3(\sha1_round/add_79_4/n104 ), .ZN(
        \sha1_round/add_79_4/n93 ) );
  NAND2_X1 \sha1_round/add_79_4/U79  ( .A1(\sha1_round/N345 ), .A2(rnd_q[152]), 
        .ZN(\sha1_round/add_79_4/n117 ) );
  INV_X2 \sha1_round/add_79_4/U78  ( .A(\sha1_round/N340 ), .ZN(
        \sha1_round/add_79_4/n192 ) );
  NAND2_X1 \sha1_round/add_79_4/U77  ( .A1(\sha1_round/add_79_4/n111 ), .A2(
        \sha1_round/add_79_4/n157 ), .ZN(\sha1_round/add_79_4/n162 ) );
  INV_X4 \sha1_round/add_79_4/U76  ( .A(\sha1_round/add_79_4/n101 ), .ZN(
        \sha1_round/add_79_4/n107 ) );
  NAND2_X1 \sha1_round/add_79_4/U75  ( .A1(\sha1_round/N335 ), .A2(rnd_q[142]), 
        .ZN(\sha1_round/add_79_4/n150 ) );
  AND2_X2 \sha1_round/add_79_4/U74  ( .A1(\sha1_round/N331 ), .A2(rnd_q[138]), 
        .ZN(\sha1_round/add_79_4/n5 ) );
  INV_X4 \sha1_round/add_79_4/U73  ( .A(\sha1_round/add_79_4/n91 ), .ZN(
        \sha1_round/add_79_4/n32 ) );
  NAND2_X2 \sha1_round/add_79_4/U72  ( .A1(\sha1_round/add_79_4/n24 ), .A2(
        \sha1_round/add_79_4/n25 ), .ZN(sha1_round_wire[157]) );
  NOR3_X2 \sha1_round/add_79_4/U71  ( .A1(\sha1_round/add_79_4/n237 ), .A2(
        \sha1_round/add_79_4/n147 ), .A3(\sha1_round/add_79_4/n148 ), .ZN(
        \sha1_round/add_79_4/n231 ) );
  NOR2_X2 \sha1_round/add_79_4/U70  ( .A1(\sha1_round/add_79_4/n49 ), .A2(
        \sha1_round/add_79_4/n291 ), .ZN(\sha1_round/add_79_4/n290 ) );
  NOR2_X2 \sha1_round/add_79_4/U69  ( .A1(\sha1_round/add_79_4/n3 ), .A2(
        \sha1_round/add_79_4/n290 ), .ZN(\sha1_round/add_79_4/n286 ) );
  INV_X4 \sha1_round/add_79_4/U68  ( .A(\sha1_round/add_79_4/n213 ), .ZN(
        \sha1_round/add_79_4/n28 ) );
  NAND2_X2 \sha1_round/add_79_4/U67  ( .A1(\sha1_round/add_79_4/n32 ), .A2(
        \sha1_round/add_79_4/n33 ), .ZN(\sha1_round/add_79_4/n35 ) );
  NAND2_X2 \sha1_round/add_79_4/U66  ( .A1(\sha1_round/add_79_4/n206 ), .A2(
        \sha1_round/add_79_4/n207 ), .ZN(\sha1_round/add_79_4/n197 ) );
  NAND2_X2 \sha1_round/add_79_4/U65  ( .A1(\sha1_round/add_79_4/n227 ), .A2(
        \sha1_round/add_79_4/n228 ), .ZN(\sha1_round/add_79_4/n225 ) );
  NOR2_X2 \sha1_round/add_79_4/U64  ( .A1(\sha1_round/N330 ), .A2(rnd_q[137]), 
        .ZN(\sha1_round/add_79_4/n49 ) );
  NOR2_X2 \sha1_round/add_79_4/U63  ( .A1(\sha1_round/add_79_4/n56 ), .A2(
        \sha1_round/add_79_4/n317 ), .ZN(\sha1_round/add_79_4/n274 ) );
  INV_X4 \sha1_round/add_79_4/U62  ( .A(\sha1_round/add_79_4/n68 ), .ZN(
        \sha1_round/add_79_4/n340 ) );
  NAND2_X2 \sha1_round/add_79_4/U61  ( .A1(\sha1_round/N341 ), .A2(rnd_q[148]), 
        .ZN(\sha1_round/add_79_4/n184 ) );
  NOR2_X2 \sha1_round/add_79_4/U60  ( .A1(\sha1_round/add_79_4/n219 ), .A2(
        \sha1_round/add_79_4/n224 ), .ZN(\sha1_round/add_79_4/n205 ) );
  NOR2_X2 \sha1_round/add_79_4/U59  ( .A1(\sha1_round/add_79_4/n218 ), .A2(
        \sha1_round/add_79_4/n219 ), .ZN(\sha1_round/add_79_4/n217 ) );
  NOR2_X2 \sha1_round/add_79_4/U58  ( .A1(\sha1_round/add_79_4/n107 ), .A2(
        \sha1_round/add_79_4/n105 ), .ZN(\sha1_round/add_79_4/n104 ) );
  INV_X4 \sha1_round/add_79_4/U57  ( .A(\sha1_round/add_79_4/n127 ), .ZN(
        \sha1_round/add_79_4/n113 ) );
  NOR2_X2 \sha1_round/add_79_4/U56  ( .A1(\sha1_round/add_79_4/n222 ), .A2(
        \sha1_round/add_79_4/n223 ), .ZN(\sha1_round/add_79_4/n221 ) );
  NAND2_X2 \sha1_round/add_79_4/U55  ( .A1(\sha1_round/add_79_4/n22 ), .A2(
        \sha1_round/add_79_4/n23 ), .ZN(\sha1_round/add_79_4/n25 ) );
  INV_X4 \sha1_round/add_79_4/U54  ( .A(\sha1_round/add_79_4/n240 ), .ZN(
        \sha1_round/add_79_4/n238 ) );
  NOR2_X2 \sha1_round/add_79_4/U53  ( .A1(\sha1_round/N328 ), .A2(rnd_q[135]), 
        .ZN(\sha1_round/add_79_4/n48 ) );
  NAND2_X2 \sha1_round/add_79_4/U52  ( .A1(\sha1_round/add_79_4/n288 ), .A2(
        \sha1_round/add_79_4/n289 ), .ZN(\sha1_round/add_79_4/n233 ) );
  INV_X4 \sha1_round/add_79_4/U51  ( .A(\sha1_round/add_79_4/n225 ), .ZN(
        \sha1_round/add_79_4/n219 ) );
  XNOR2_X1 \sha1_round/add_79_4/U50  ( .A(\sha1_round/add_79_4/n266 ), .B(
        \sha1_round/add_79_4/n250 ), .ZN(sha1_round_wire[144]) );
  NAND2_X1 \sha1_round/add_79_4/U49  ( .A1(\sha1_round/N324 ), .A2(rnd_q[131]), 
        .ZN(\sha1_round/add_79_4/n312 ) );
  OR2_X4 \sha1_round/add_79_4/U48  ( .A1(\sha1_round/N344 ), .A2(rnd_q[151]), 
        .ZN(\sha1_round/add_79_4/n158 ) );
  NAND3_X4 \sha1_round/add_79_4/U47  ( .A1(\sha1_round/add_79_4/n309 ), .A2(
        \sha1_round/add_79_4/n310 ), .A3(\sha1_round/add_79_4/n311 ), .ZN(
        \sha1_round/add_79_4/n304 ) );
  NAND2_X4 \sha1_round/add_79_4/U46  ( .A1(\sha1_round/add_79_4/n12 ), .A2(
        \sha1_round/add_79_4/n304 ), .ZN(\sha1_round/add_79_4/n273 ) );
  NAND2_X4 \sha1_round/add_79_4/U45  ( .A1(\sha1_round/add_79_4/n259 ), .A2(
        \sha1_round/add_79_4/n260 ), .ZN(\sha1_round/add_79_4/n248 ) );
  INV_X2 \sha1_round/add_79_4/U44  ( .A(\sha1_round/N331 ), .ZN(
        \sha1_round/add_79_4/n288 ) );
  AND2_X4 \sha1_round/add_79_4/U43  ( .A1(\sha1_round/add_79_4/n136 ), .A2(
        \sha1_round/add_79_4/n145 ), .ZN(\sha1_round/add_79_4/n2 ) );
  NOR2_X2 \sha1_round/add_79_4/U42  ( .A1(\sha1_round/add_79_4/n297 ), .A2(
        \sha1_round/add_79_4/n8 ), .ZN(\sha1_round/add_79_4/n293 ) );
  NOR2_X2 \sha1_round/add_79_4/U41  ( .A1(\sha1_round/add_79_4/n293 ), .A2(
        \sha1_round/add_79_4/n10 ), .ZN(\sha1_round/add_79_4/n291 ) );
  NAND2_X2 \sha1_round/add_79_4/U40  ( .A1(\sha1_round/add_79_4/n141 ), .A2(
        \sha1_round/add_79_4/n142 ), .ZN(\sha1_round/add_79_4/n24 ) );
  NAND2_X2 \sha1_round/add_79_4/U39  ( .A1(\sha1_round/add_79_4/n192 ), .A2(
        \sha1_round/add_79_4/n193 ), .ZN(\sha1_round/add_79_4/n178 ) );
  NOR2_X2 \sha1_round/add_79_4/U38  ( .A1(rnd_q[143]), .A2(\sha1_round/N336 ), 
        .ZN(\sha1_round/add_79_4/n218 ) );
  NAND2_X2 \sha1_round/add_79_4/U37  ( .A1(\sha1_round/add_79_4/n209 ), .A2(
        \sha1_round/add_79_4/n210 ), .ZN(\sha1_round/add_79_4/n97 ) );
  NOR2_X2 \sha1_round/add_79_4/U36  ( .A1(\sha1_round/N335 ), .A2(rnd_q[142]), 
        .ZN(\sha1_round/add_79_4/n47 ) );
  INV_X4 \sha1_round/add_79_4/U35  ( .A(\sha1_round/N327 ), .ZN(
        \sha1_round/add_79_4/n321 ) );
  NAND2_X2 \sha1_round/add_79_4/U34  ( .A1(\sha1_round/add_79_4/n321 ), .A2(
        \sha1_round/add_79_4/n322 ), .ZN(\sha1_round/add_79_4/n307 ) );
  NAND2_X2 \sha1_round/add_79_4/U33  ( .A1(\sha1_round/add_79_4/n326 ), .A2(
        \sha1_round/add_79_4/n327 ), .ZN(\sha1_round/add_79_4/n313 ) );
  NOR2_X2 \sha1_round/add_79_4/U32  ( .A1(\sha1_round/add_79_4/n339 ), .A2(
        \sha1_round/add_79_4/n340 ), .ZN(\sha1_round/add_79_4/n338 ) );
  NAND2_X2 \sha1_round/add_79_4/U31  ( .A1(\sha1_round/add_79_4/n143 ), .A2(
        \sha1_round/add_79_4/n144 ), .ZN(\sha1_round/add_79_4/n141 ) );
  NOR2_X2 \sha1_round/add_79_4/U30  ( .A1(\sha1_round/add_79_4/n278 ), .A2(
        \sha1_round/add_79_4/n48 ), .ZN(\sha1_round/add_79_4/n276 ) );
  NOR2_X4 \sha1_round/add_79_4/U29  ( .A1(\sha1_round/add_79_4/n96 ), .A2(
        \sha1_round/add_79_4/n155 ), .ZN(\sha1_round/add_79_4/n130 ) );
  NAND2_X4 \sha1_round/add_79_4/U28  ( .A1(\sha1_round/add_79_4/n248 ), .A2(
        \sha1_round/add_79_4/n249 ), .ZN(\sha1_round/add_79_4/n246 ) );
  NAND2_X4 \sha1_round/add_79_4/U27  ( .A1(\sha1_round/add_79_4/n246 ), .A2(
        \sha1_round/add_79_4/n247 ), .ZN(\sha1_round/add_79_4/n209 ) );
  NAND2_X4 \sha1_round/add_79_4/U26  ( .A1(\sha1_round/add_79_4/n200 ), .A2(
        \sha1_round/add_79_4/n201 ), .ZN(\sha1_round/add_79_4/n153 ) );
  NAND2_X4 \sha1_round/add_79_4/U25  ( .A1(\sha1_round/add_79_4/n153 ), .A2(
        \sha1_round/add_79_4/n154 ), .ZN(\sha1_round/add_79_4/n199 ) );
  NOR2_X4 \sha1_round/add_79_4/U24  ( .A1(\sha1_round/add_79_4/n267 ), .A2(
        \sha1_round/add_79_4/n268 ), .ZN(\sha1_round/add_79_4/n250 ) );
  XNOR2_X1 \sha1_round/add_79_4/U23  ( .A(\sha1_round/add_79_4/n165 ), .B(
        \sha1_round/add_79_4/n191 ), .ZN(sha1_round_wire[152]) );
  NOR2_X4 \sha1_round/add_79_4/U22  ( .A1(\sha1_round/add_79_4/n122 ), .A2(
        \sha1_round/add_79_4/n121 ), .ZN(\sha1_round/add_79_4/n118 ) );
  NAND2_X4 \sha1_round/add_79_4/U21  ( .A1(\sha1_round/add_79_4/n161 ), .A2(
        \sha1_round/add_79_4/n162 ), .ZN(\sha1_round/add_79_4/n159 ) );
  NAND2_X4 \sha1_round/add_79_4/U20  ( .A1(\sha1_round/add_79_4/n171 ), .A2(
        \sha1_round/add_79_4/n172 ), .ZN(\sha1_round/add_79_4/n163 ) );
  NAND2_X4 \sha1_round/add_79_4/U19  ( .A1(\sha1_round/add_79_4/n170 ), .A2(
        \sha1_round/add_79_4/n163 ), .ZN(\sha1_round/add_79_4/n166 ) );
  NAND2_X4 \sha1_round/add_79_4/U18  ( .A1(\sha1_round/add_79_4/n211 ), .A2(
        \sha1_round/add_79_4/n154 ), .ZN(\sha1_round/add_79_4/n100 ) );
  INV_X8 \sha1_round/add_79_4/U17  ( .A(\sha1_round/add_79_4/n100 ), .ZN(
        \sha1_round/add_79_4/n136 ) );
  NAND2_X4 \sha1_round/add_79_4/U16  ( .A1(\sha1_round/add_79_4/n13 ), .A2(
        \sha1_round/add_79_4/n97 ), .ZN(\sha1_round/add_79_4/n232 ) );
  NAND2_X1 \sha1_round/add_79_4/U15  ( .A1(\sha1_round/add_79_4/n44 ), .A2(
        \sha1_round/add_79_4/n97 ), .ZN(\sha1_round/add_79_4/n137 ) );
  NAND2_X1 \sha1_round/add_79_4/U14  ( .A1(\sha1_round/N342 ), .A2(rnd_q[149]), 
        .ZN(\sha1_round/add_79_4/n174 ) );
  NAND3_X4 \sha1_round/add_79_4/U13  ( .A1(\sha1_round/add_79_4/n336 ), .A2(
        \sha1_round/add_79_4/n337 ), .A3(\sha1_round/add_79_4/n338 ), .ZN(
        \sha1_round/add_79_4/n64 ) );
  AND2_X2 \sha1_round/add_79_4/U12  ( .A1(\sha1_round/add_79_4/n157 ), .A2(
        \sha1_round/add_79_4/n156 ), .ZN(\sha1_round/add_79_4/n1 ) );
  INV_X1 \sha1_round/add_79_4/U11  ( .A(\sha1_round/add_79_4/n130 ), .ZN(
        \sha1_round/add_79_4/n152 ) );
  AND2_X4 \sha1_round/add_79_4/U10  ( .A1(\sha1_round/add_79_4/n307 ), .A2(
        \sha1_round/add_79_4/n313 ), .ZN(\sha1_round/add_79_4/n309 ) );
  INV_X4 \sha1_round/add_79_4/U9  ( .A(\sha1_round/add_79_4/n36 ), .ZN(
        \sha1_round/add_79_4/n110 ) );
  NOR2_X1 \sha1_round/add_79_4/U8  ( .A1(\sha1_round/add_79_4/n113 ), .A2(
        \sha1_round/add_79_4/n36 ), .ZN(\sha1_round/add_79_4/n133 ) );
  NAND2_X4 \sha1_round/add_79_4/U7  ( .A1(\sha1_round/add_79_4/n34 ), .A2(
        \sha1_round/add_79_4/n35 ), .ZN(sha1_round_wire[159]) );
  NOR2_X4 \sha1_round/add_79_4/U6  ( .A1(\sha1_round/add_79_4/n253 ), .A2(
        \sha1_round/add_79_4/n254 ), .ZN(\sha1_round/add_79_4/n251 ) );
  NAND2_X1 \sha1_round/add_79_4/U5  ( .A1(\sha1_round/add_79_4/n18 ), .A2(
        \sha1_round/add_79_4/n307 ), .ZN(\sha1_round/add_79_4/n317 ) );
  INV_X4 \sha1_round/add_79_4/U4  ( .A(\sha1_round/N343 ), .ZN(
        \sha1_round/add_79_4/n168 ) );
  NAND2_X4 \sha1_round/add_79_4/U3  ( .A1(\sha1_round/add_79_4/n30 ), .A2(
        \sha1_round/add_79_4/n31 ), .ZN(sha1_round_wire[151]) );
  NAND2_X4 \sha1_round/add_79_4/U2  ( .A1(\sha1_round/add_79_4/n28 ), .A2(
        \sha1_round/add_79_4/n29 ), .ZN(\sha1_round/add_79_4/n31 ) );
  INV_X4 \sha1_round/add_79_3/U418  ( .A(\sha1_round/N256 ), .ZN(
        \sha1_round/add_79_3/n386 ) );
  INV_X4 \sha1_round/add_79_3/U417  ( .A(\sha1_round/N288 ), .ZN(
        \sha1_round/add_79_3/n387 ) );
  NAND3_X4 \sha1_round/add_79_3/U416  ( .A1(\sha1_round/add_79_3/n383 ), .A2(
        \sha1_round/add_79_3/n378 ), .A3(\sha1_round/add_79_3/n384 ), .ZN(
        \sha1_round/add_79_3/n239 ) );
  NOR2_X4 \sha1_round/add_79_3/U415  ( .A1(\sha1_round/N259 ), .A2(
        \sha1_round/N291 ), .ZN(\sha1_round/add_79_3/n88 ) );
  NAND3_X4 \sha1_round/add_79_3/U414  ( .A1(\sha1_round/add_79_3/n239 ), .A2(
        \sha1_round/add_79_3/n16 ), .A3(\sha1_round/add_79_3/n380 ), .ZN(
        \sha1_round/add_79_3/n81 ) );
  NAND2_X2 \sha1_round/add_79_3/U413  ( .A1(\sha1_round/N284 ), .A2(
        \sha1_round/N252 ), .ZN(\sha1_round/add_79_3/n375 ) );
  NAND2_X2 \sha1_round/add_79_3/U412  ( .A1(\sha1_round/N285 ), .A2(
        \sha1_round/N253 ), .ZN(\sha1_round/add_79_3/n376 ) );
  NAND2_X2 \sha1_round/add_79_3/U411  ( .A1(\sha1_round/add_79_3/n375 ), .A2(
        \sha1_round/add_79_3/n376 ), .ZN(\sha1_round/add_79_3/n372 ) );
  INV_X4 \sha1_round/add_79_3/U410  ( .A(\sha1_round/add_79_3/n146 ), .ZN(
        \sha1_round/add_79_3/n373 ) );
  INV_X4 \sha1_round/add_79_3/U409  ( .A(\sha1_round/add_79_3/n111 ), .ZN(
        \sha1_round/add_79_3/n374 ) );
  NAND4_X2 \sha1_round/add_79_3/U408  ( .A1(\sha1_round/add_79_3/n372 ), .A2(
        \sha1_round/add_79_3/n314 ), .A3(\sha1_round/add_79_3/n373 ), .A4(
        \sha1_round/add_79_3/n374 ), .ZN(\sha1_round/add_79_3/n371 ) );
  NAND2_X2 \sha1_round/add_79_3/U407  ( .A1(\sha1_round/N287 ), .A2(
        \sha1_round/N255 ), .ZN(\sha1_round/add_79_3/n309 ) );
  INV_X4 \sha1_round/add_79_3/U406  ( .A(\sha1_round/N293 ), .ZN(
        \sha1_round/add_79_3/n367 ) );
  INV_X4 \sha1_round/add_79_3/U405  ( .A(\sha1_round/N261 ), .ZN(
        \sha1_round/add_79_3/n368 ) );
  INV_X4 \sha1_round/add_79_3/U404  ( .A(\sha1_round/add_79_3/n74 ), .ZN(
        \sha1_round/add_79_3/n365 ) );
  NOR2_X4 \sha1_round/add_79_3/U403  ( .A1(\sha1_round/add_79_3/n364 ), .A2(
        \sha1_round/add_79_3/n365 ), .ZN(\sha1_round/add_79_3/n360 ) );
  INV_X4 \sha1_round/add_79_3/U402  ( .A(\sha1_round/add_79_3/n348 ), .ZN(
        \sha1_round/add_79_3/n359 ) );
  INV_X4 \sha1_round/add_79_3/U401  ( .A(\sha1_round/N294 ), .ZN(
        \sha1_round/add_79_3/n362 ) );
  XNOR2_X2 \sha1_round/add_79_3/U400  ( .A(\sha1_round/add_79_3/n360 ), .B(
        \sha1_round/add_79_3/n361 ), .ZN(\sha1_round/N326 ) );
  INV_X4 \sha1_round/add_79_3/U399  ( .A(\sha1_round/N295 ), .ZN(
        \sha1_round/add_79_3/n356 ) );
  NAND2_X2 \sha1_round/add_79_3/U398  ( .A1(\sha1_round/add_79_3/n76 ), .A2(
        \sha1_round/add_79_3/n74 ), .ZN(\sha1_round/add_79_3/n346 ) );
  NOR2_X4 \sha1_round/add_79_3/U397  ( .A1(\sha1_round/add_79_3/n321 ), .A2(
        \sha1_round/add_79_3/n322 ), .ZN(\sha1_round/add_79_3/n347 ) );
  NAND3_X4 \sha1_round/add_79_3/U396  ( .A1(\sha1_round/add_79_3/n347 ), .A2(
        \sha1_round/add_79_3/n346 ), .A3(\sha1_round/add_79_3/n73 ), .ZN(
        \sha1_round/add_79_3/n245 ) );
  INV_X4 \sha1_round/add_79_3/U395  ( .A(\sha1_round/add_79_3/n84 ), .ZN(
        \sha1_round/add_79_3/n342 ) );
  INV_X4 \sha1_round/add_79_3/U394  ( .A(\sha1_round/N297 ), .ZN(
        \sha1_round/add_79_3/n336 ) );
  NAND2_X2 \sha1_round/add_79_3/U393  ( .A1(\sha1_round/add_79_3/n336 ), .A2(
        \sha1_round/add_79_3/n337 ), .ZN(\sha1_round/add_79_3/n298 ) );
  NAND2_X2 \sha1_round/add_79_3/U392  ( .A1(\sha1_round/N297 ), .A2(
        \sha1_round/N265 ), .ZN(\sha1_round/add_79_3/n294 ) );
  NAND2_X2 \sha1_round/add_79_3/U391  ( .A1(\sha1_round/add_79_3/n52 ), .A2(
        \sha1_round/add_79_3/n294 ), .ZN(\sha1_round/add_79_3/n335 ) );
  INV_X4 \sha1_round/add_79_3/U390  ( .A(\sha1_round/N298 ), .ZN(
        \sha1_round/add_79_3/n331 ) );
  XNOR2_X2 \sha1_round/add_79_3/U389  ( .A(\sha1_round/add_79_3/n329 ), .B(
        \sha1_round/add_79_3/n330 ), .ZN(\sha1_round/N330 ) );
  INV_X4 \sha1_round/add_79_3/U388  ( .A(\sha1_round/N299 ), .ZN(
        \sha1_round/add_79_3/n326 ) );
  INV_X4 \sha1_round/add_79_3/U387  ( .A(\sha1_round/N267 ), .ZN(
        \sha1_round/add_79_3/n327 ) );
  XNOR2_X2 \sha1_round/add_79_3/U386  ( .A(\sha1_round/add_79_3/n324 ), .B(
        \sha1_round/add_79_3/n325 ), .ZN(\sha1_round/N331 ) );
  INV_X4 \sha1_round/add_79_3/U385  ( .A(\sha1_round/add_79_3/n323 ), .ZN(
        \sha1_round/add_79_3/n246 ) );
  INV_X4 \sha1_round/add_79_3/U384  ( .A(\sha1_round/add_79_3/n314 ), .ZN(
        \sha1_round/add_79_3/n107 ) );
  NAND2_X2 \sha1_round/add_79_3/U383  ( .A1(\sha1_round/N284 ), .A2(
        \sha1_round/N252 ), .ZN(\sha1_round/add_79_3/n313 ) );
  NAND2_X2 \sha1_round/add_79_3/U382  ( .A1(\sha1_round/N254 ), .A2(
        \sha1_round/N286 ), .ZN(\sha1_round/add_79_3/n312 ) );
  INV_X4 \sha1_round/add_79_3/U381  ( .A(\sha1_round/add_79_3/n309 ), .ZN(
        \sha1_round/add_79_3/n106 ) );
  NAND2_X2 \sha1_round/add_79_3/U380  ( .A1(\sha1_round/add_79_3/n306 ), .A2(
        \sha1_round/add_79_3/n307 ), .ZN(\sha1_round/add_79_3/n240 ) );
  INV_X4 \sha1_round/add_79_3/U379  ( .A(\sha1_round/add_79_3/n235 ), .ZN(
        \sha1_round/add_79_3/n296 ) );
  NOR2_X4 \sha1_round/add_79_3/U378  ( .A1(\sha1_round/add_79_3/n58 ), .A2(
        \sha1_round/add_79_3/n295 ), .ZN(\sha1_round/add_79_3/n277 ) );
  NOR2_X4 \sha1_round/add_79_3/U377  ( .A1(\sha1_round/N268 ), .A2(
        \sha1_round/N300 ), .ZN(\sha1_round/add_79_3/n276 ) );
  XNOR2_X2 \sha1_round/add_79_3/U376  ( .A(\sha1_round/add_79_3/n288 ), .B(
        \sha1_round/add_79_3/n289 ), .ZN(\sha1_round/N332 ) );
  INV_X4 \sha1_round/add_79_3/U375  ( .A(\sha1_round/N301 ), .ZN(
        \sha1_round/add_79_3/n285 ) );
  XNOR2_X2 \sha1_round/add_79_3/U374  ( .A(\sha1_round/add_79_3/n284 ), .B(
        \sha1_round/add_79_3/n8 ), .ZN(\sha1_round/N333 ) );
  NAND2_X2 \sha1_round/add_79_3/U373  ( .A1(\sha1_round/add_79_3/n269 ), .A2(
        \sha1_round/add_79_3/n259 ), .ZN(\sha1_round/add_79_3/n268 ) );
  INV_X4 \sha1_round/add_79_3/U372  ( .A(\sha1_round/N303 ), .ZN(
        \sha1_round/add_79_3/n265 ) );
  INV_X4 \sha1_round/add_79_3/U371  ( .A(\sha1_round/N271 ), .ZN(
        \sha1_round/add_79_3/n266 ) );
  XNOR2_X2 \sha1_round/add_79_3/U370  ( .A(\sha1_round/add_79_3/n262 ), .B(
        \sha1_round/add_79_3/n263 ), .ZN(\sha1_round/N335 ) );
  INV_X4 \sha1_round/add_79_3/U369  ( .A(\sha1_round/add_79_3/n376 ), .ZN(
        \sha1_round/add_79_3/n261 ) );
  XNOR2_X2 \sha1_round/add_79_3/U368  ( .A(\sha1_round/add_79_3/n313 ), .B(
        \sha1_round/add_79_3/n260 ), .ZN(\sha1_round/N317 ) );
  NAND2_X2 \sha1_round/add_79_3/U367  ( .A1(\sha1_round/N304 ), .A2(
        \sha1_round/N272 ), .ZN(\sha1_round/add_79_3/n226 ) );
  NAND2_X2 \sha1_round/add_79_3/U366  ( .A1(\sha1_round/add_79_3/n226 ), .A2(
        \sha1_round/add_79_3/n228 ), .ZN(\sha1_round/add_79_3/n229 ) );
  INV_X4 \sha1_round/add_79_3/U365  ( .A(\sha1_round/add_79_3/n257 ), .ZN(
        \sha1_round/add_79_3/n256 ) );
  NOR2_X4 \sha1_round/add_79_3/U364  ( .A1(\sha1_round/add_79_3/n253 ), .A2(
        \sha1_round/add_79_3/n252 ), .ZN(\sha1_round/add_79_3/n230 ) );
  INV_X4 \sha1_round/add_79_3/U363  ( .A(\sha1_round/add_79_3/n250 ), .ZN(
        \sha1_round/add_79_3/n249 ) );
  NAND3_X4 \sha1_round/add_79_3/U362  ( .A1(\sha1_round/add_79_3/n232 ), .A2(
        \sha1_round/add_79_3/n230 ), .A3(\sha1_round/add_79_3/n231 ), .ZN(
        \sha1_round/add_79_3/n148 ) );
  INV_X4 \sha1_round/add_79_3/U361  ( .A(\sha1_round/add_79_3/n218 ), .ZN(
        \sha1_round/add_79_3/n228 ) );
  INV_X4 \sha1_round/add_79_3/U360  ( .A(\sha1_round/N305 ), .ZN(
        \sha1_round/add_79_3/n224 ) );
  INV_X4 \sha1_round/add_79_3/U359  ( .A(\sha1_round/N273 ), .ZN(
        \sha1_round/add_79_3/n225 ) );
  XNOR2_X2 \sha1_round/add_79_3/U358  ( .A(\sha1_round/add_79_3/n222 ), .B(
        \sha1_round/add_79_3/n223 ), .ZN(\sha1_round/N337 ) );
  INV_X4 \sha1_round/add_79_3/U357  ( .A(\sha1_round/add_79_3/n208 ), .ZN(
        \sha1_round/add_79_3/n220 ) );
  NAND2_X2 \sha1_round/add_79_3/U356  ( .A1(\sha1_round/add_79_3/n215 ), .A2(
        \sha1_round/add_79_3/n216 ), .ZN(\sha1_round/add_79_3/n211 ) );
  INV_X4 \sha1_round/add_79_3/U355  ( .A(\sha1_round/N306 ), .ZN(
        \sha1_round/add_79_3/n213 ) );
  INV_X4 \sha1_round/add_79_3/U354  ( .A(\sha1_round/N274 ), .ZN(
        \sha1_round/add_79_3/n214 ) );
  NAND2_X2 \sha1_round/add_79_3/U353  ( .A1(\sha1_round/N306 ), .A2(
        \sha1_round/N274 ), .ZN(\sha1_round/add_79_3/n209 ) );
  NAND2_X2 \sha1_round/add_79_3/U352  ( .A1(\sha1_round/add_79_3/n200 ), .A2(
        \sha1_round/add_79_3/n209 ), .ZN(\sha1_round/add_79_3/n212 ) );
  XNOR2_X2 \sha1_round/add_79_3/U351  ( .A(\sha1_round/add_79_3/n211 ), .B(
        \sha1_round/add_79_3/n212 ), .ZN(\sha1_round/N338 ) );
  INV_X4 \sha1_round/add_79_3/U350  ( .A(\sha1_round/add_79_3/n198 ), .ZN(
        \sha1_round/add_79_3/n206 ) );
  NAND2_X2 \sha1_round/add_79_3/U349  ( .A1(\sha1_round/add_79_3/n204 ), .A2(
        \sha1_round/add_79_3/n205 ), .ZN(\sha1_round/add_79_3/n202 ) );
  NAND2_X2 \sha1_round/add_79_3/U348  ( .A1(\sha1_round/N307 ), .A2(
        \sha1_round/N275 ), .ZN(\sha1_round/add_79_3/n150 ) );
  NAND2_X2 \sha1_round/add_79_3/U347  ( .A1(\sha1_round/add_79_3/n197 ), .A2(
        \sha1_round/add_79_3/n150 ), .ZN(\sha1_round/add_79_3/n203 ) );
  NAND2_X2 \sha1_round/add_79_3/U346  ( .A1(\sha1_round/N308 ), .A2(
        \sha1_round/N276 ), .ZN(\sha1_round/add_79_3/n174 ) );
  INV_X4 \sha1_round/add_79_3/U345  ( .A(\sha1_round/N308 ), .ZN(
        \sha1_round/add_79_3/n195 ) );
  INV_X4 \sha1_round/add_79_3/U344  ( .A(\sha1_round/N276 ), .ZN(
        \sha1_round/add_79_3/n196 ) );
  XNOR2_X2 \sha1_round/add_79_3/U343  ( .A(\sha1_round/add_79_3/n186 ), .B(
        \sha1_round/add_79_3/n194 ), .ZN(\sha1_round/N340 ) );
  NAND2_X2 \sha1_round/add_79_3/U342  ( .A1(\sha1_round/add_79_3/n178 ), .A2(
        \sha1_round/add_79_3/n186 ), .ZN(\sha1_round/add_79_3/n193 ) );
  INV_X4 \sha1_round/add_79_3/U341  ( .A(\sha1_round/N309 ), .ZN(
        \sha1_round/add_79_3/n191 ) );
  INV_X4 \sha1_round/add_79_3/U340  ( .A(\sha1_round/N277 ), .ZN(
        \sha1_round/add_79_3/n192 ) );
  NAND2_X2 \sha1_round/add_79_3/U339  ( .A1(\sha1_round/add_79_3/n172 ), .A2(
        \sha1_round/add_79_3/n179 ), .ZN(\sha1_round/add_79_3/n183 ) );
  INV_X4 \sha1_round/add_79_3/U338  ( .A(\sha1_round/add_79_3/n179 ), .ZN(
        \sha1_round/add_79_3/n176 ) );
  NAND2_X2 \sha1_round/add_79_3/U337  ( .A1(\sha1_round/add_79_3/n185 ), .A2(
        \sha1_round/add_79_3/n186 ), .ZN(\sha1_round/add_79_3/n184 ) );
  NAND2_X2 \sha1_round/add_79_3/U336  ( .A1(\sha1_round/add_79_3/n183 ), .A2(
        \sha1_round/add_79_3/n184 ), .ZN(\sha1_round/add_79_3/n181 ) );
  NAND2_X2 \sha1_round/add_79_3/U335  ( .A1(\sha1_round/N311 ), .A2(
        \sha1_round/N279 ), .ZN(\sha1_round/add_79_3/n157 ) );
  INV_X4 \sha1_round/add_79_3/U334  ( .A(\sha1_round/N311 ), .ZN(
        \sha1_round/add_79_3/n166 ) );
  INV_X4 \sha1_round/add_79_3/U333  ( .A(\sha1_round/N279 ), .ZN(
        \sha1_round/add_79_3/n167 ) );
  NAND2_X2 \sha1_round/add_79_3/U332  ( .A1(\sha1_round/add_79_3/n166 ), .A2(
        \sha1_round/add_79_3/n167 ), .ZN(\sha1_round/add_79_3/n158 ) );
  NOR2_X4 \sha1_round/add_79_3/U331  ( .A1(\sha1_round/add_79_3/n164 ), .A2(
        \sha1_round/add_79_3/n165 ), .ZN(\sha1_round/add_79_3/n161 ) );
  NAND2_X2 \sha1_round/add_79_3/U330  ( .A1(\sha1_round/N312 ), .A2(
        \sha1_round/N280 ), .ZN(\sha1_round/add_79_3/n136 ) );
  INV_X4 \sha1_round/add_79_3/U329  ( .A(\sha1_round/add_79_3/n153 ), .ZN(
        \sha1_round/add_79_3/n151 ) );
  NAND2_X2 \sha1_round/add_79_3/U328  ( .A1(\sha1_round/add_79_3/n64 ), .A2(
        \sha1_round/add_79_3/n65 ), .ZN(\sha1_round/add_79_3/n127 ) );
  INV_X4 \sha1_round/add_79_3/U327  ( .A(\sha1_round/add_79_3/n150 ), .ZN(
        \sha1_round/add_79_3/n149 ) );
  NAND4_X2 \sha1_round/add_79_3/U326  ( .A1(\sha1_round/add_79_3/n129 ), .A2(
        \sha1_round/add_79_3/n136 ), .A3(\sha1_round/add_79_3/n127 ), .A4(
        \sha1_round/add_79_3/n126 ), .ZN(\sha1_round/add_79_3/n147 ) );
  NAND2_X2 \sha1_round/add_79_3/U325  ( .A1(\sha1_round/N313 ), .A2(
        \sha1_round/N281 ), .ZN(\sha1_round/add_79_3/n134 ) );
  NAND2_X2 \sha1_round/add_79_3/U324  ( .A1(\sha1_round/N286 ), .A2(
        \sha1_round/N254 ), .ZN(\sha1_round/add_79_3/n110 ) );
  NAND2_X2 \sha1_round/add_79_3/U323  ( .A1(\sha1_round/add_79_3/n374 ), .A2(
        \sha1_round/add_79_3/n110 ), .ZN(\sha1_round/add_79_3/n145 ) );
  NAND2_X2 \sha1_round/add_79_3/U322  ( .A1(\sha1_round/add_79_3/n62 ), .A2(
        \sha1_round/add_79_3/n376 ), .ZN(\sha1_round/add_79_3/n113 ) );
  XNOR2_X2 \sha1_round/add_79_3/U321  ( .A(\sha1_round/add_79_3/n145 ), .B(
        \sha1_round/add_79_3/n113 ), .ZN(\sha1_round/N318 ) );
  NAND2_X2 \sha1_round/add_79_3/U320  ( .A1(\sha1_round/N314 ), .A2(
        \sha1_round/N282 ), .ZN(\sha1_round/add_79_3/n135 ) );
  NAND2_X2 \sha1_round/add_79_3/U319  ( .A1(\sha1_round/add_79_3/n135 ), .A2(
        \sha1_round/add_79_3/n139 ), .ZN(\sha1_round/add_79_3/n141 ) );
  XNOR2_X2 \sha1_round/add_79_3/U318  ( .A(\sha1_round/add_79_3/n140 ), .B(
        \sha1_round/add_79_3/n141 ), .ZN(\sha1_round/N346 ) );
  INV_X4 \sha1_round/add_79_3/U317  ( .A(\sha1_round/add_79_3/n139 ), .ZN(
        \sha1_round/add_79_3/n133 ) );
  INV_X4 \sha1_round/add_79_3/U316  ( .A(\sha1_round/add_79_3/n138 ), .ZN(
        \sha1_round/add_79_3/n137 ) );
  INV_X4 \sha1_round/add_79_3/U315  ( .A(\sha1_round/add_79_3/n135 ), .ZN(
        \sha1_round/add_79_3/n131 ) );
  NAND2_X2 \sha1_round/add_79_3/U314  ( .A1(\sha1_round/add_79_3/n128 ), .A2(
        \sha1_round/add_79_3/n121 ), .ZN(\sha1_round/add_79_3/n117 ) );
  INV_X4 \sha1_round/add_79_3/U313  ( .A(\sha1_round/add_79_3/n121 ), .ZN(
        \sha1_round/add_79_3/n125 ) );
  NAND2_X2 \sha1_round/add_79_3/U312  ( .A1(\sha1_round/add_79_3/n120 ), .A2(
        \sha1_round/add_79_3/n121 ), .ZN(\sha1_round/add_79_3/n119 ) );
  NAND4_X2 \sha1_round/add_79_3/U311  ( .A1(\sha1_round/add_79_3/n116 ), .A2(
        \sha1_round/add_79_3/n117 ), .A3(\sha1_round/add_79_3/n118 ), .A4(
        \sha1_round/add_79_3/n119 ), .ZN(\sha1_round/add_79_3/n114 ) );
  XNOR2_X2 \sha1_round/add_79_3/U310  ( .A(\sha1_round/N315 ), .B(
        \sha1_round/N283 ), .ZN(\sha1_round/add_79_3/n115 ) );
  XNOR2_X2 \sha1_round/add_79_3/U309  ( .A(\sha1_round/add_79_3/n114 ), .B(
        \sha1_round/add_79_3/n115 ), .ZN(\sha1_round/N347 ) );
  INV_X4 \sha1_round/add_79_3/U308  ( .A(\sha1_round/add_79_3/n113 ), .ZN(
        \sha1_round/add_79_3/n112 ) );
  INV_X4 \sha1_round/add_79_3/U307  ( .A(\sha1_round/add_79_3/n110 ), .ZN(
        \sha1_round/add_79_3/n109 ) );
  XNOR2_X2 \sha1_round/add_79_3/U306  ( .A(\sha1_round/add_79_3/n104 ), .B(
        \sha1_round/add_79_3/n105 ), .ZN(\sha1_round/N319 ) );
  NAND2_X2 \sha1_round/add_79_3/U305  ( .A1(\sha1_round/N288 ), .A2(
        \sha1_round/N256 ), .ZN(\sha1_round/add_79_3/n98 ) );
  NAND2_X2 \sha1_round/add_79_3/U304  ( .A1(\sha1_round/add_79_3/n98 ), .A2(
        \sha1_round/add_79_3/n100 ), .ZN(\sha1_round/add_79_3/n103 ) );
  NAND2_X2 \sha1_round/add_79_3/U303  ( .A1(\sha1_round/add_79_3/n93 ), .A2(
        \sha1_round/add_79_3/n95 ), .ZN(\sha1_round/add_79_3/n97 ) );
  INV_X4 \sha1_round/add_79_3/U302  ( .A(\sha1_round/add_79_3/n102 ), .ZN(
        \sha1_round/add_79_3/n100 ) );
  XNOR2_X2 \sha1_round/add_79_3/U301  ( .A(\sha1_round/add_79_3/n97 ), .B(
        \sha1_round/add_79_3/n94 ), .ZN(\sha1_round/N321 ) );
  NAND2_X2 \sha1_round/add_79_3/U300  ( .A1(\sha1_round/add_79_3/n94 ), .A2(
        \sha1_round/add_79_3/n95 ), .ZN(\sha1_round/add_79_3/n92 ) );
  XNOR2_X2 \sha1_round/add_79_3/U299  ( .A(\sha1_round/add_79_3/n63 ), .B(
        \sha1_round/add_79_3/n91 ), .ZN(\sha1_round/N322 ) );
  NAND2_X2 \sha1_round/add_79_3/U298  ( .A1(\sha1_round/add_79_3/n76 ), .A2(
        \sha1_round/add_79_3/n77 ), .ZN(\sha1_round/add_79_3/n82 ) );
  INV_X4 \sha1_round/add_79_3/U297  ( .A(\sha1_round/add_79_3/n81 ), .ZN(
        \sha1_round/add_79_3/n79 ) );
  NAND2_X2 \sha1_round/add_79_3/U296  ( .A1(\sha1_round/add_79_3/n77 ), .A2(
        \sha1_round/add_79_3/n78 ), .ZN(\sha1_round/add_79_3/n75 ) );
  NAND2_X2 \sha1_round/add_79_3/U295  ( .A1(\sha1_round/add_79_3/n75 ), .A2(
        \sha1_round/add_79_3/n76 ), .ZN(\sha1_round/add_79_3/n71 ) );
  XNOR2_X2 \sha1_round/add_79_3/U294  ( .A(\sha1_round/add_79_3/n71 ), .B(
        \sha1_round/add_79_3/n72 ), .ZN(\sha1_round/N325 ) );
  NAND2_X4 \sha1_round/add_79_3/U293  ( .A1(\sha1_round/add_79_3/n234 ), .A2(
        \sha1_round/add_79_3/n233 ), .ZN(\sha1_round/add_79_3/n232 ) );
  NAND3_X2 \sha1_round/add_79_3/U292  ( .A1(\sha1_round/add_79_3/n19 ), .A2(
        \sha1_round/add_79_3/n350 ), .A3(\sha1_round/add_79_3/n351 ), .ZN(
        \sha1_round/add_79_3/n303 ) );
  NAND2_X4 \sha1_round/add_79_3/U291  ( .A1(\sha1_round/add_79_3/n66 ), .A2(
        \sha1_round/add_79_3/n148 ), .ZN(\sha1_round/add_79_3/n180 ) );
  NAND2_X1 \sha1_round/add_79_3/U290  ( .A1(\sha1_round/add_79_3/n148 ), .A2(
        \sha1_round/add_79_3/n207 ), .ZN(\sha1_round/add_79_3/n216 ) );
  NAND2_X1 \sha1_round/add_79_3/U289  ( .A1(\sha1_round/add_79_3/n206 ), .A2(
        \sha1_round/add_79_3/n148 ), .ZN(\sha1_round/add_79_3/n205 ) );
  NAND2_X1 \sha1_round/add_79_3/U288  ( .A1(\sha1_round/N299 ), .A2(
        \sha1_round/N267 ), .ZN(\sha1_round/add_79_3/n291 ) );
  NAND2_X1 \sha1_round/add_79_3/U287  ( .A1(\sha1_round/add_79_3/n291 ), .A2(
        \sha1_round/add_79_3/n247 ), .ZN(\sha1_round/add_79_3/n325 ) );
  NAND3_X2 \sha1_round/add_79_3/U286  ( .A1(\sha1_round/add_79_3/n249 ), .A2(
        \sha1_round/add_79_3/n248 ), .A3(\sha1_round/add_79_3/n247 ), .ZN(
        \sha1_round/add_79_3/n231 ) );
  NAND2_X4 \sha1_round/add_79_3/U285  ( .A1(\sha1_round/add_79_3/n286 ), .A2(
        \sha1_round/add_79_3/n285 ), .ZN(\sha1_round/add_79_3/n274 ) );
  NOR2_X1 \sha1_round/add_79_3/U284  ( .A1(\sha1_round/add_79_3/n87 ), .A2(
        \sha1_round/add_79_3/n385 ), .ZN(\sha1_round/add_79_3/n86 ) );
  NAND3_X2 \sha1_round/add_79_3/U283  ( .A1(\sha1_round/add_79_3/n50 ), .A2(
        \sha1_round/add_79_3/n302 ), .A3(\sha1_round/add_79_3/n245 ), .ZN(
        \sha1_round/add_79_3/n341 ) );
  NAND2_X1 \sha1_round/add_79_3/U282  ( .A1(\sha1_round/add_79_3/n302 ), .A2(
        \sha1_round/add_79_3/n20 ), .ZN(\sha1_round/add_79_3/n355 ) );
  NAND2_X2 \sha1_round/add_79_3/U281  ( .A1(\sha1_round/add_79_3/n148 ), .A2(
        \sha1_round/add_79_3/n228 ), .ZN(\sha1_round/add_79_3/n227 ) );
  NAND2_X4 \sha1_round/add_79_3/U280  ( .A1(\sha1_round/add_79_3/n327 ), .A2(
        \sha1_round/add_79_3/n326 ), .ZN(\sha1_round/add_79_3/n247 ) );
  NOR2_X2 \sha1_round/add_79_3/U279  ( .A1(\sha1_round/add_79_3/n276 ), .A2(
        \sha1_round/add_79_3/n69 ), .ZN(\sha1_round/add_79_3/n289 ) );
  NAND2_X1 \sha1_round/add_79_3/U278  ( .A1(\sha1_round/add_79_3/n208 ), .A2(
        \sha1_round/add_79_3/n219 ), .ZN(\sha1_round/add_79_3/n223 ) );
  NAND3_X2 \sha1_round/add_79_3/U277  ( .A1(\sha1_round/N272 ), .A2(
        \sha1_round/N304 ), .A3(\sha1_round/add_79_3/n219 ), .ZN(
        \sha1_round/add_79_3/n210 ) );
  NAND2_X1 \sha1_round/add_79_3/U276  ( .A1(\sha1_round/N309 ), .A2(
        \sha1_round/N277 ), .ZN(\sha1_round/add_79_3/n173 ) );
  NAND2_X1 \sha1_round/add_79_3/U275  ( .A1(\sha1_round/N258 ), .A2(
        \sha1_round/N290 ), .ZN(\sha1_round/add_79_3/n381 ) );
  NAND2_X1 \sha1_round/add_79_3/U274  ( .A1(\sha1_round/add_79_3/n73 ), .A2(
        \sha1_round/add_79_3/n74 ), .ZN(\sha1_round/add_79_3/n72 ) );
  NAND2_X4 \sha1_round/add_79_3/U273  ( .A1(\sha1_round/add_79_3/n266 ), .A2(
        \sha1_round/add_79_3/n265 ), .ZN(\sha1_round/add_79_3/n251 ) );
  NAND2_X1 \sha1_round/add_79_3/U272  ( .A1(\sha1_round/N310 ), .A2(
        \sha1_round/N278 ), .ZN(\sha1_round/add_79_3/n160 ) );
  NOR3_X2 \sha1_round/add_79_3/U271  ( .A1(\sha1_round/add_79_3/n13 ), .A2(
        \sha1_round/add_79_3/n146 ), .A3(\sha1_round/add_79_3/n111 ), .ZN(
        \sha1_round/add_79_3/n310 ) );
  OR2_X4 \sha1_round/add_79_3/U270  ( .A1(\sha1_round/N252 ), .A2(
        \sha1_round/N284 ), .ZN(\sha1_round/add_79_3/n70 ) );
  AND2_X2 \sha1_round/add_79_3/U269  ( .A1(\sha1_round/add_79_3/n313 ), .A2(
        \sha1_round/add_79_3/n70 ), .ZN(\sha1_round/N316 ) );
  AND2_X2 \sha1_round/add_79_3/U268  ( .A1(\sha1_round/N300 ), .A2(
        \sha1_round/N268 ), .ZN(\sha1_round/add_79_3/n69 ) );
  AND2_X2 \sha1_round/add_79_3/U267  ( .A1(\sha1_round/N290 ), .A2(
        \sha1_round/N258 ), .ZN(\sha1_round/add_79_3/n68 ) );
  NOR2_X2 \sha1_round/add_79_3/U266  ( .A1(\sha1_round/add_79_3/n275 ), .A2(
        \sha1_round/add_79_3/n276 ), .ZN(\sha1_round/add_79_3/n273 ) );
  NOR2_X2 \sha1_round/add_79_3/U265  ( .A1(\sha1_round/add_79_3/n310 ), .A2(
        \sha1_round/add_79_3/n311 ), .ZN(\sha1_round/add_79_3/n306 ) );
  NOR2_X2 \sha1_round/add_79_3/U264  ( .A1(\sha1_round/add_79_3/n106 ), .A2(
        \sha1_round/add_79_3/n308 ), .ZN(\sha1_round/add_79_3/n307 ) );
  NAND2_X1 \sha1_round/add_79_3/U263  ( .A1(\sha1_round/N302 ), .A2(
        \sha1_round/N270 ), .ZN(\sha1_round/add_79_3/n259 ) );
  NOR2_X2 \sha1_round/add_79_3/U262  ( .A1(\sha1_round/add_79_3/n88 ), .A2(
        \sha1_round/add_79_3/n381 ), .ZN(\sha1_round/add_79_3/n323 ) );
  OR2_X2 \sha1_round/add_79_3/U261  ( .A1(\sha1_round/N314 ), .A2(
        \sha1_round/N282 ), .ZN(\sha1_round/add_79_3/n139 ) );
  OR2_X2 \sha1_round/add_79_3/U260  ( .A1(\sha1_round/N312 ), .A2(
        \sha1_round/N280 ), .ZN(\sha1_round/add_79_3/n152 ) );
  OR2_X2 \sha1_round/add_79_3/U259  ( .A1(\sha1_round/N313 ), .A2(
        \sha1_round/N281 ), .ZN(\sha1_round/add_79_3/n138 ) );
  NOR2_X2 \sha1_round/add_79_3/U258  ( .A1(\sha1_round/N253 ), .A2(
        \sha1_round/N285 ), .ZN(\sha1_round/add_79_3/n146 ) );
  NOR2_X1 \sha1_round/add_79_3/U257  ( .A1(\sha1_round/add_79_3/n111 ), .A2(
        \sha1_round/add_79_3/n112 ), .ZN(\sha1_round/add_79_3/n108 ) );
  INV_X4 \sha1_round/add_79_3/U256  ( .A(\sha1_round/add_79_3/n244 ), .ZN(
        \sha1_round/add_79_3/n87 ) );
  NOR2_X1 \sha1_round/add_79_3/U255  ( .A1(\sha1_round/add_79_3/n102 ), .A2(
        \sha1_round/add_79_3/n96 ), .ZN(\sha1_round/add_79_3/n318 ) );
  AND2_X2 \sha1_round/add_79_3/U254  ( .A1(\sha1_round/add_79_3/n92 ), .A2(
        \sha1_round/add_79_3/n93 ), .ZN(\sha1_round/add_79_3/n63 ) );
  NOR2_X1 \sha1_round/add_79_3/U253  ( .A1(\sha1_round/add_79_3/n176 ), .A2(
        \sha1_round/add_79_3/n188 ), .ZN(\sha1_round/add_79_3/n185 ) );
  NOR2_X2 \sha1_round/add_79_3/U252  ( .A1(\sha1_round/add_79_3/n258 ), .A2(
        \sha1_round/add_79_3/n259 ), .ZN(\sha1_round/add_79_3/n252 ) );
  NOR3_X2 \sha1_round/add_79_3/U251  ( .A1(\sha1_round/add_79_3/n241 ), .A2(
        \sha1_round/add_79_3/n4 ), .A3(\sha1_round/add_79_3/n243 ), .ZN(
        \sha1_round/add_79_3/n304 ) );
  AND2_X2 \sha1_round/add_79_3/U250  ( .A1(\sha1_round/add_79_3/n136 ), .A2(
        \sha1_round/add_79_3/n129 ), .ZN(\sha1_round/add_79_3/n144 ) );
  NOR2_X2 \sha1_round/add_79_3/U249  ( .A1(\sha1_round/add_79_3/n133 ), .A2(
        \sha1_round/add_79_3/n137 ), .ZN(\sha1_round/add_79_3/n121 ) );
  NAND2_X2 \sha1_round/add_79_3/U248  ( .A1(\sha1_round/add_79_3/n341 ), .A2(
        \sha1_round/add_79_3/n299 ), .ZN(\sha1_round/add_79_3/n340 ) );
  NOR2_X2 \sha1_round/add_79_3/U247  ( .A1(\sha1_round/add_79_3/n322 ), .A2(
        \sha1_round/add_79_3/n348 ), .ZN(\sha1_round/add_79_3/n242 ) );
  NOR2_X1 \sha1_round/add_79_3/U246  ( .A1(\sha1_round/add_79_3/n68 ), .A2(
        \sha1_round/add_79_3/n90 ), .ZN(\sha1_round/add_79_3/n91 ) );
  NOR2_X2 \sha1_round/add_79_3/U245  ( .A1(\sha1_round/add_79_3/n89 ), .A2(
        \sha1_round/add_79_3/n68 ), .ZN(\sha1_round/add_79_3/n85 ) );
  NOR2_X2 \sha1_round/add_79_3/U244  ( .A1(\sha1_round/add_79_3/n220 ), .A2(
        \sha1_round/add_79_3/n221 ), .ZN(\sha1_round/add_79_3/n215 ) );
  NOR2_X2 \sha1_round/add_79_3/U243  ( .A1(\sha1_round/add_79_3/n108 ), .A2(
        \sha1_round/add_79_3/n109 ), .ZN(\sha1_round/add_79_3/n104 ) );
  NOR2_X2 \sha1_round/add_79_3/U242  ( .A1(\sha1_round/add_79_3/n319 ), .A2(
        \sha1_round/add_79_3/n320 ), .ZN(\sha1_round/add_79_3/n351 ) );
  XNOR2_X2 \sha1_round/add_79_3/U241  ( .A(\sha1_round/add_79_3/n202 ), .B(
        \sha1_round/add_79_3/n203 ), .ZN(\sha1_round/N339 ) );
  NOR2_X1 \sha1_round/add_79_3/U240  ( .A1(\sha1_round/add_79_3/n125 ), .A2(
        \sha1_round/add_79_3/n126 ), .ZN(\sha1_round/add_79_3/n124 ) );
  NOR2_X1 \sha1_round/add_79_3/U239  ( .A1(\sha1_round/add_79_3/n125 ), .A2(
        \sha1_round/add_79_3/n127 ), .ZN(\sha1_round/add_79_3/n123 ) );
  NOR2_X2 \sha1_round/add_79_3/U238  ( .A1(\sha1_round/add_79_3/n123 ), .A2(
        \sha1_round/add_79_3/n124 ), .ZN(\sha1_round/add_79_3/n118 ) );
  NOR2_X1 \sha1_round/add_79_3/U237  ( .A1(\sha1_round/add_79_3/n352 ), .A2(
        \sha1_round/add_79_3/n81 ), .ZN(\sha1_round/add_79_3/n349 ) );
  AND4_X2 \sha1_round/add_79_3/U236  ( .A1(\sha1_round/add_79_3/n304 ), .A2(
        \sha1_round/add_79_3/n5 ), .A3(\sha1_round/add_79_3/n239 ), .A4(
        \sha1_round/add_79_3/n305 ), .ZN(\sha1_round/add_79_3/n58 ) );
  NOR2_X1 \sha1_round/add_79_3/U235  ( .A1(\sha1_round/add_79_3/n359 ), .A2(
        \sha1_round/add_79_3/n321 ), .ZN(\sha1_round/add_79_3/n361 ) );
  NOR2_X1 \sha1_round/add_79_3/U234  ( .A1(\sha1_round/add_79_3/n107 ), .A2(
        \sha1_round/add_79_3/n312 ), .ZN(\sha1_round/add_79_3/n311 ) );
  NOR3_X1 \sha1_round/add_79_3/U233  ( .A1(\sha1_round/add_79_3/n376 ), .A2(
        \sha1_round/add_79_3/n107 ), .A3(\sha1_round/add_79_3/n111 ), .ZN(
        \sha1_round/add_79_3/n308 ) );
  NAND3_X2 \sha1_round/add_79_3/U232  ( .A1(\sha1_round/N254 ), .A2(
        \sha1_round/N286 ), .A3(\sha1_round/add_79_3/n314 ), .ZN(
        \sha1_round/add_79_3/n370 ) );
  OR2_X4 \sha1_round/add_79_3/U231  ( .A1(\sha1_round/N296 ), .A2(
        \sha1_round/N264 ), .ZN(\sha1_round/add_79_3/n299 ) );
  NAND3_X2 \sha1_round/add_79_3/U230  ( .A1(\sha1_round/N257 ), .A2(
        \sha1_round/N289 ), .A3(\sha1_round/add_79_3/n378 ), .ZN(
        \sha1_round/add_79_3/n382 ) );
  OR2_X4 \sha1_round/add_79_3/U229  ( .A1(\sha1_round/N307 ), .A2(
        \sha1_round/N275 ), .ZN(\sha1_round/add_79_3/n197 ) );
  INV_X1 \sha1_round/add_79_3/U228  ( .A(\sha1_round/add_79_3/n96 ), .ZN(
        \sha1_round/add_79_3/n95 ) );
  AND2_X2 \sha1_round/add_79_3/U227  ( .A1(\sha1_round/add_79_3/n157 ), .A2(
        \sha1_round/add_79_3/n158 ), .ZN(\sha1_round/add_79_3/n60 ) );
  INV_X1 \sha1_round/add_79_3/U226  ( .A(\sha1_round/add_79_3/n251 ), .ZN(
        \sha1_round/add_79_3/n258 ) );
  INV_X4 \sha1_round/add_79_3/U225  ( .A(\sha1_round/add_79_3/n197 ), .ZN(
        \sha1_round/add_79_3/n67 ) );
  INV_X1 \sha1_round/add_79_3/U224  ( .A(\sha1_round/add_79_3/n177 ), .ZN(
        \sha1_round/add_79_3/n175 ) );
  AND2_X2 \sha1_round/add_79_3/U223  ( .A1(\sha1_round/add_79_3/n301 ), .A2(
        \sha1_round/add_79_3/n299 ), .ZN(\sha1_round/add_79_3/n57 ) );
  XNOR2_X2 \sha1_round/add_79_3/U222  ( .A(\sha1_round/add_79_3/n344 ), .B(
        \sha1_round/add_79_3/n57 ), .ZN(\sha1_round/N328 ) );
  NOR2_X1 \sha1_round/add_79_3/U221  ( .A1(\sha1_round/add_79_3/n133 ), .A2(
        \sha1_round/add_79_3/n134 ), .ZN(\sha1_round/add_79_3/n132 ) );
  NOR3_X1 \sha1_round/add_79_3/U220  ( .A1(\sha1_round/add_79_3/n130 ), .A2(
        \sha1_round/add_79_3/n131 ), .A3(\sha1_round/add_79_3/n132 ), .ZN(
        \sha1_round/add_79_3/n116 ) );
  NOR2_X1 \sha1_round/add_79_3/U219  ( .A1(\sha1_round/add_79_3/n125 ), .A2(
        \sha1_round/add_79_3/n136 ), .ZN(\sha1_round/add_79_3/n130 ) );
  OR2_X4 \sha1_round/add_79_3/U218  ( .A1(\sha1_round/add_79_3/n146 ), .A2(
        \sha1_round/add_79_3/n313 ), .ZN(\sha1_round/add_79_3/n62 ) );
  NOR2_X1 \sha1_round/add_79_3/U217  ( .A1(\sha1_round/add_79_3/n106 ), .A2(
        \sha1_round/add_79_3/n107 ), .ZN(\sha1_round/add_79_3/n105 ) );
  INV_X1 \sha1_round/add_79_3/U216  ( .A(\sha1_round/add_79_3/n259 ), .ZN(
        \sha1_round/add_79_3/n280 ) );
  INV_X1 \sha1_round/add_79_3/U215  ( .A(\sha1_round/add_79_3/n254 ), .ZN(
        \sha1_round/add_79_3/n264 ) );
  NOR2_X1 \sha1_round/add_79_3/U214  ( .A1(\sha1_round/add_79_3/n261 ), .A2(
        \sha1_round/add_79_3/n146 ), .ZN(\sha1_round/add_79_3/n260 ) );
  XOR2_X2 \sha1_round/add_79_3/U213  ( .A(\sha1_round/add_79_3/n349 ), .B(
        \sha1_round/add_79_3/n82 ), .Z(\sha1_round/N324 ) );
  NOR2_X1 \sha1_round/add_79_3/U212  ( .A1(\sha1_round/add_79_3/n83 ), .A2(
        \sha1_round/add_79_3/n84 ), .ZN(\sha1_round/add_79_3/n352 ) );
  NOR2_X1 \sha1_round/add_79_3/U211  ( .A1(\sha1_round/add_79_3/n264 ), .A2(
        \sha1_round/add_79_3/n258 ), .ZN(\sha1_round/add_79_3/n263 ) );
  AND3_X4 \sha1_round/add_79_3/U210  ( .A1(\sha1_round/add_79_3/n200 ), .A2(
        \sha1_round/add_79_3/n197 ), .A3(\sha1_round/add_79_3/n201 ), .ZN(
        \sha1_round/add_79_3/n64 ) );
  NAND2_X1 \sha1_round/add_79_3/U209  ( .A1(\sha1_round/N298 ), .A2(
        \sha1_round/N266 ), .ZN(\sha1_round/add_79_3/n292 ) );
  XNOR2_X2 \sha1_round/add_79_3/U208  ( .A(\sha1_round/add_79_3/n51 ), .B(
        \sha1_round/add_79_3/n1 ), .ZN(\sha1_round/N344 ) );
  INV_X1 \sha1_round/add_79_3/U207  ( .A(\sha1_round/add_79_3/n101 ), .ZN(
        \sha1_round/add_79_3/n83 ) );
  INV_X1 \sha1_round/add_79_3/U206  ( .A(\sha1_round/add_79_3/n122 ), .ZN(
        \sha1_round/add_79_3/n120 ) );
  NOR2_X2 \sha1_round/add_79_3/U205  ( .A1(\sha1_round/add_79_3/n272 ), .A2(
        \sha1_round/add_79_3/n18 ), .ZN(\sha1_round/add_79_3/n267 ) );
  NOR2_X2 \sha1_round/add_79_3/U204  ( .A1(\sha1_round/add_79_3/n276 ), .A2(
        \sha1_round/add_79_3/n272 ), .ZN(\sha1_round/add_79_3/n287 ) );
  NAND2_X2 \sha1_round/add_79_3/U203  ( .A1(\sha1_round/N291 ), .A2(
        \sha1_round/N259 ), .ZN(\sha1_round/add_79_3/n244 ) );
  NOR2_X2 \sha1_round/add_79_3/U202  ( .A1(\sha1_round/add_79_3/n250 ), .A2(
        \sha1_round/add_79_3/n290 ), .ZN(\sha1_round/add_79_3/n55 ) );
  INV_X4 \sha1_round/add_79_3/U201  ( .A(\sha1_round/add_79_3/n4 ), .ZN(
        \sha1_round/add_79_3/n50 ) );
  INV_X1 \sha1_round/add_79_3/U200  ( .A(\sha1_round/add_79_3/n274 ), .ZN(
        \sha1_round/add_79_3/n283 ) );
  NOR2_X2 \sha1_round/add_79_3/U199  ( .A1(\sha1_round/add_79_3/n161 ), .A2(
        \sha1_round/add_79_3/n163 ), .ZN(\sha1_round/add_79_3/n169 ) );
  NAND2_X4 \sha1_round/add_79_3/U198  ( .A1(\sha1_round/add_79_3/n331 ), .A2(
        \sha1_round/add_79_3/n332 ), .ZN(\sha1_round/add_79_3/n297 ) );
  NAND2_X1 \sha1_round/add_79_3/U197  ( .A1(\sha1_round/add_79_3/n297 ), .A2(
        \sha1_round/add_79_3/n292 ), .ZN(\sha1_round/add_79_3/n330 ) );
  NAND2_X1 \sha1_round/add_79_3/U196  ( .A1(\sha1_round/N305 ), .A2(
        \sha1_round/N273 ), .ZN(\sha1_round/add_79_3/n208 ) );
  NOR2_X4 \sha1_round/add_79_3/U195  ( .A1(\sha1_round/add_79_3/n277 ), .A2(
        \sha1_round/add_79_3/n55 ), .ZN(\sha1_round/add_79_3/n288 ) );
  NOR2_X4 \sha1_round/add_79_3/U194  ( .A1(\sha1_round/add_79_3/n277 ), .A2(
        \sha1_round/add_79_3/n55 ), .ZN(\sha1_round/add_79_3/n272 ) );
  NAND2_X1 \sha1_round/add_79_3/U193  ( .A1(\sha1_round/add_79_3/n201 ), .A2(
        \sha1_round/add_79_3/n200 ), .ZN(\sha1_round/add_79_3/n204 ) );
  INV_X4 \sha1_round/add_79_3/U192  ( .A(\sha1_round/add_79_3/n165 ), .ZN(
        \sha1_round/add_79_3/n187 ) );
  NOR2_X2 \sha1_round/add_79_3/U191  ( .A1(\sha1_round/add_79_3/n287 ), .A2(
        \sha1_round/add_79_3/n69 ), .ZN(\sha1_round/add_79_3/n284 ) );
  INV_X4 \sha1_round/add_79_3/U190  ( .A(\sha1_round/add_79_3/n180 ), .ZN(
        \sha1_round/add_79_3/n164 ) );
  INV_X4 \sha1_round/add_79_3/U189  ( .A(\sha1_round/add_79_3/n178 ), .ZN(
        \sha1_round/add_79_3/n188 ) );
  NAND2_X1 \sha1_round/add_79_3/U188  ( .A1(\sha1_round/add_79_3/n174 ), .A2(
        \sha1_round/add_79_3/n178 ), .ZN(\sha1_round/add_79_3/n194 ) );
  NAND2_X2 \sha1_round/add_79_3/U187  ( .A1(\sha1_round/add_79_3/n69 ), .A2(
        \sha1_round/add_79_3/n274 ), .ZN(\sha1_round/add_79_3/n270 ) );
  INV_X4 \sha1_round/add_79_3/U186  ( .A(\sha1_round/add_79_3/n279 ), .ZN(
        \sha1_round/add_79_3/n47 ) );
  NAND2_X4 \sha1_round/add_79_3/U185  ( .A1(\sha1_round/add_79_3/n48 ), .A2(
        \sha1_round/add_79_3/n49 ), .ZN(\sha1_round/N334 ) );
  NAND2_X4 \sha1_round/add_79_3/U184  ( .A1(\sha1_round/add_79_3/n46 ), .A2(
        \sha1_round/add_79_3/n47 ), .ZN(\sha1_round/add_79_3/n49 ) );
  NAND2_X2 \sha1_round/add_79_3/U183  ( .A1(\sha1_round/add_79_3/n278 ), .A2(
        \sha1_round/add_79_3/n279 ), .ZN(\sha1_round/add_79_3/n48 ) );
  NAND2_X4 \sha1_round/add_79_3/U182  ( .A1(\sha1_round/add_79_3/n10 ), .A2(
        \sha1_round/add_79_3/n178 ), .ZN(\sha1_round/add_79_3/n163 ) );
  NAND4_X2 \sha1_round/add_79_3/U181  ( .A1(\sha1_round/add_79_3/n126 ), .A2(
        \sha1_round/add_79_3/n144 ), .A3(\sha1_round/add_79_3/n127 ), .A4(
        \sha1_round/add_79_3/n122 ), .ZN(\sha1_round/add_79_3/n143 ) );
  NOR2_X2 \sha1_round/add_79_3/U180  ( .A1(\sha1_round/add_79_3/n198 ), .A2(
        \sha1_round/add_79_3/n67 ), .ZN(\sha1_round/add_79_3/n66 ) );
  AND2_X4 \sha1_round/add_79_3/U179  ( .A1(\sha1_round/add_79_3/n151 ), .A2(
        \sha1_round/add_79_3/n152 ), .ZN(\sha1_round/add_79_3/n65 ) );
  INV_X4 \sha1_round/add_79_3/U178  ( .A(\sha1_round/add_79_3/n60 ), .ZN(
        \sha1_round/add_79_3/n43 ) );
  INV_X4 \sha1_round/add_79_3/U177  ( .A(\sha1_round/add_79_3/n168 ), .ZN(
        \sha1_round/add_79_3/n42 ) );
  NAND2_X4 \sha1_round/add_79_3/U176  ( .A1(\sha1_round/add_79_3/n45 ), .A2(
        \sha1_round/add_79_3/n44 ), .ZN(\sha1_round/N343 ) );
  NAND2_X4 \sha1_round/add_79_3/U175  ( .A1(\sha1_round/add_79_3/n42 ), .A2(
        \sha1_round/add_79_3/n43 ), .ZN(\sha1_round/add_79_3/n45 ) );
  NAND2_X2 \sha1_round/add_79_3/U174  ( .A1(\sha1_round/add_79_3/n168 ), .A2(
        \sha1_round/add_79_3/n60 ), .ZN(\sha1_round/add_79_3/n44 ) );
  NAND2_X1 \sha1_round/add_79_3/U173  ( .A1(\sha1_round/add_79_3/n173 ), .A2(
        \sha1_round/add_79_3/n179 ), .ZN(\sha1_round/add_79_3/n190 ) );
  INV_X2 \sha1_round/add_79_3/U172  ( .A(\sha1_round/add_79_3/n190 ), .ZN(
        \sha1_round/add_79_3/n39 ) );
  INV_X4 \sha1_round/add_79_3/U171  ( .A(\sha1_round/add_79_3/n189 ), .ZN(
        \sha1_round/add_79_3/n38 ) );
  NAND2_X4 \sha1_round/add_79_3/U170  ( .A1(\sha1_round/add_79_3/n40 ), .A2(
        \sha1_round/add_79_3/n41 ), .ZN(\sha1_round/N341 ) );
  NAND2_X4 \sha1_round/add_79_3/U169  ( .A1(\sha1_round/add_79_3/n38 ), .A2(
        \sha1_round/add_79_3/n39 ), .ZN(\sha1_round/add_79_3/n41 ) );
  NAND2_X2 \sha1_round/add_79_3/U168  ( .A1(\sha1_round/add_79_3/n189 ), .A2(
        \sha1_round/add_79_3/n190 ), .ZN(\sha1_round/add_79_3/n40 ) );
  NAND3_X2 \sha1_round/add_79_3/U167  ( .A1(\sha1_round/add_79_3/n238 ), .A2(
        \sha1_round/add_79_3/n305 ), .A3(\sha1_round/add_79_3/n15 ), .ZN(
        \sha1_round/add_79_3/n233 ) );
  NAND2_X1 \sha1_round/add_79_3/U166  ( .A1(\sha1_round/add_79_3/n160 ), .A2(
        \sha1_round/add_79_3/n177 ), .ZN(\sha1_round/add_79_3/n182 ) );
  INV_X1 \sha1_round/add_79_3/U165  ( .A(\sha1_round/add_79_3/n182 ), .ZN(
        \sha1_round/add_79_3/n35 ) );
  INV_X4 \sha1_round/add_79_3/U164  ( .A(\sha1_round/add_79_3/n181 ), .ZN(
        \sha1_round/add_79_3/n34 ) );
  INV_X1 \sha1_round/add_79_3/U163  ( .A(\sha1_round/add_79_3/n86 ), .ZN(
        \sha1_round/add_79_3/n31 ) );
  INV_X4 \sha1_round/add_79_3/U162  ( .A(\sha1_round/add_79_3/n85 ), .ZN(
        \sha1_round/add_79_3/n30 ) );
  NAND2_X4 \sha1_round/add_79_3/U161  ( .A1(\sha1_round/add_79_3/n32 ), .A2(
        \sha1_round/add_79_3/n33 ), .ZN(\sha1_round/N323 ) );
  NAND2_X4 \sha1_round/add_79_3/U160  ( .A1(\sha1_round/add_79_3/n30 ), .A2(
        \sha1_round/add_79_3/n31 ), .ZN(\sha1_round/add_79_3/n33 ) );
  NAND2_X2 \sha1_round/add_79_3/U159  ( .A1(\sha1_round/add_79_3/n85 ), .A2(
        \sha1_round/add_79_3/n86 ), .ZN(\sha1_round/add_79_3/n32 ) );
  NAND3_X4 \sha1_round/add_79_3/U158  ( .A1(\sha1_round/add_79_3/n208 ), .A2(
        \sha1_round/add_79_3/n209 ), .A3(\sha1_round/add_79_3/n210 ), .ZN(
        \sha1_round/add_79_3/n201 ) );
  NAND2_X4 \sha1_round/add_79_3/U157  ( .A1(\sha1_round/add_79_3/n29 ), .A2(
        \sha1_round/add_79_3/n201 ), .ZN(\sha1_round/add_79_3/n199 ) );
  AND2_X2 \sha1_round/add_79_3/U156  ( .A1(\sha1_round/add_79_3/n200 ), .A2(
        \sha1_round/add_79_3/n197 ), .ZN(\sha1_round/add_79_3/n29 ) );
  NAND3_X2 \sha1_round/add_79_3/U155  ( .A1(\sha1_round/add_79_3/n245 ), .A2(
        \sha1_round/add_79_3/n303 ), .A3(\sha1_round/add_79_3/n12 ), .ZN(
        \sha1_round/add_79_3/n300 ) );
  NAND2_X4 \sha1_round/add_79_3/U154  ( .A1(\sha1_round/add_79_3/n328 ), .A2(
        \sha1_round/add_79_3/n292 ), .ZN(\sha1_round/add_79_3/n324 ) );
  INV_X4 \sha1_round/add_79_3/U153  ( .A(\sha1_round/N262 ), .ZN(
        \sha1_round/add_79_3/n363 ) );
  NAND2_X1 \sha1_round/add_79_3/U152  ( .A1(\sha1_round/N303 ), .A2(
        \sha1_round/N271 ), .ZN(\sha1_round/add_79_3/n254 ) );
  NAND2_X1 \sha1_round/add_79_3/U151  ( .A1(\sha1_round/add_79_3/n282 ), .A2(
        \sha1_round/add_79_3/n256 ), .ZN(\sha1_round/add_79_3/n269 ) );
  NOR2_X2 \sha1_round/add_79_3/U150  ( .A1(\sha1_round/add_79_3/n90 ), .A2(
        \sha1_round/add_79_3/n63 ), .ZN(\sha1_round/add_79_3/n89 ) );
  NOR2_X2 \sha1_round/add_79_3/U149  ( .A1(\sha1_round/add_79_3/n267 ), .A2(
        \sha1_round/add_79_3/n268 ), .ZN(\sha1_round/add_79_3/n262 ) );
  INV_X1 \sha1_round/add_79_3/U148  ( .A(\sha1_round/add_79_3/n88 ), .ZN(
        \sha1_round/add_79_3/n377 ) );
  NAND2_X2 \sha1_round/add_79_3/U147  ( .A1(\sha1_round/add_79_3/n76 ), .A2(
        \sha1_round/add_79_3/n80 ), .ZN(\sha1_round/add_79_3/n28 ) );
  NOR2_X2 \sha1_round/add_79_3/U146  ( .A1(\sha1_round/add_79_3/n319 ), .A2(
        \sha1_round/add_79_3/n320 ), .ZN(\sha1_round/add_79_3/n316 ) );
  NOR2_X2 \sha1_round/add_79_3/U145  ( .A1(\sha1_round/N291 ), .A2(
        \sha1_round/N259 ), .ZN(\sha1_round/add_79_3/n385 ) );
  NOR2_X2 \sha1_round/add_79_3/U144  ( .A1(\sha1_round/add_79_3/n321 ), .A2(
        \sha1_round/add_79_3/n322 ), .ZN(\sha1_round/add_79_3/n315 ) );
  AND2_X4 \sha1_round/add_79_3/U143  ( .A1(\sha1_round/add_79_3/n134 ), .A2(
        \sha1_round/add_79_3/n138 ), .ZN(\sha1_round/add_79_3/n27 ) );
  XNOR2_X2 \sha1_round/add_79_3/U142  ( .A(\sha1_round/add_79_3/n56 ), .B(
        \sha1_round/add_79_3/n27 ), .ZN(\sha1_round/N345 ) );
  NOR2_X2 \sha1_round/add_79_3/U141  ( .A1(\sha1_round/add_79_3/n28 ), .A2(
        \sha1_round/add_79_3/n81 ), .ZN(\sha1_round/add_79_3/n26 ) );
  OR2_X4 \sha1_round/add_79_3/U140  ( .A1(\sha1_round/N292 ), .A2(
        \sha1_round/N260 ), .ZN(\sha1_round/add_79_3/n77 ) );
  INV_X1 \sha1_round/add_79_3/U139  ( .A(\sha1_round/add_79_3/n129 ), .ZN(
        \sha1_round/add_79_3/n128 ) );
  NOR2_X2 \sha1_round/add_79_3/U138  ( .A1(\sha1_round/add_79_3/n26 ), .A2(
        \sha1_round/add_79_3/n366 ), .ZN(\sha1_round/add_79_3/n364 ) );
  NOR2_X1 \sha1_round/add_79_3/U137  ( .A1(\sha1_round/add_79_3/n345 ), .A2(
        \sha1_round/add_79_3/n341 ), .ZN(\sha1_round/add_79_3/n344 ) );
  NAND2_X2 \sha1_round/add_79_3/U136  ( .A1(\sha1_round/N294 ), .A2(
        \sha1_round/N262 ), .ZN(\sha1_round/add_79_3/n348 ) );
  NAND2_X1 \sha1_round/add_79_3/U135  ( .A1(\sha1_round/add_79_3/n336 ), .A2(
        \sha1_round/add_79_3/n337 ), .ZN(\sha1_round/add_79_3/n52 ) );
  OR2_X2 \sha1_round/add_79_3/U134  ( .A1(\sha1_round/add_79_3/n293 ), .A2(
        \sha1_round/add_79_3/n294 ), .ZN(\sha1_round/add_79_3/n61 ) );
  AND3_X4 \sha1_round/add_79_3/U133  ( .A1(\sha1_round/add_79_3/n61 ), .A2(
        \sha1_round/add_79_3/n292 ), .A3(\sha1_round/add_79_3/n291 ), .ZN(
        \sha1_round/add_79_3/n250 ) );
  OR2_X4 \sha1_round/add_79_3/U132  ( .A1(\sha1_round/N310 ), .A2(
        \sha1_round/N278 ), .ZN(\sha1_round/add_79_3/n177 ) );
  INV_X4 \sha1_round/add_79_3/U131  ( .A(\sha1_round/add_79_3/n353 ), .ZN(
        \sha1_round/add_79_3/n23 ) );
  NAND2_X4 \sha1_round/add_79_3/U130  ( .A1(\sha1_round/add_79_3/n24 ), .A2(
        \sha1_round/add_79_3/n25 ), .ZN(\sha1_round/N327 ) );
  NAND2_X4 \sha1_round/add_79_3/U129  ( .A1(\sha1_round/add_79_3/n23 ), .A2(
        \sha1_round/add_79_3/n355 ), .ZN(\sha1_round/add_79_3/n25 ) );
  NAND2_X2 \sha1_round/add_79_3/U128  ( .A1(\sha1_round/add_79_3/n353 ), .A2(
        \sha1_round/add_79_3/n354 ), .ZN(\sha1_round/add_79_3/n24 ) );
  NAND2_X2 \sha1_round/add_79_3/U127  ( .A1(\sha1_round/add_79_3/n14 ), .A2(
        \sha1_round/add_79_3/n377 ), .ZN(\sha1_round/add_79_3/n84 ) );
  INV_X4 \sha1_round/add_79_3/U126  ( .A(\sha1_round/N269 ), .ZN(
        \sha1_round/add_79_3/n286 ) );
  NAND2_X1 \sha1_round/add_79_3/U125  ( .A1(\sha1_round/N301 ), .A2(
        \sha1_round/N269 ), .ZN(\sha1_round/add_79_3/n271 ) );
  NAND2_X2 \sha1_round/add_79_3/U124  ( .A1(\sha1_round/add_79_3/n181 ), .A2(
        \sha1_round/add_79_3/n182 ), .ZN(\sha1_round/add_79_3/n36 ) );
  OR2_X4 \sha1_round/add_79_3/U123  ( .A1(\sha1_round/N287 ), .A2(
        \sha1_round/N255 ), .ZN(\sha1_round/add_79_3/n314 ) );
  INV_X4 \sha1_round/add_79_3/U122  ( .A(\sha1_round/add_79_3/n297 ), .ZN(
        \sha1_round/add_79_3/n293 ) );
  INV_X4 \sha1_round/add_79_3/U121  ( .A(\sha1_round/add_79_3/n21 ), .ZN(
        \sha1_round/add_79_3/n237 ) );
  NAND3_X2 \sha1_round/add_79_3/U120  ( .A1(\sha1_round/add_79_3/n22 ), .A2(
        \sha1_round/add_79_3/n247 ), .A3(\sha1_round/add_79_3/n297 ), .ZN(
        \sha1_round/add_79_3/n21 ) );
  NAND2_X2 \sha1_round/add_79_3/U119  ( .A1(\sha1_round/add_79_3/n164 ), .A2(
        \sha1_round/add_79_3/n65 ), .ZN(\sha1_round/add_79_3/n122 ) );
  NAND2_X1 \sha1_round/add_79_3/U118  ( .A1(\sha1_round/add_79_3/n79 ), .A2(
        \sha1_round/add_79_3/n80 ), .ZN(\sha1_round/add_79_3/n78 ) );
  NAND2_X1 \sha1_round/add_79_3/U117  ( .A1(\sha1_round/add_79_3/n17 ), .A2(
        \sha1_round/add_79_3/n356 ), .ZN(\sha1_round/add_79_3/n20 ) );
  INV_X1 \sha1_round/add_79_3/U116  ( .A(\sha1_round/add_79_3/n7 ), .ZN(
        \sha1_round/add_79_3/n18 ) );
  INV_X4 \sha1_round/add_79_3/U115  ( .A(\sha1_round/add_79_3/n219 ), .ZN(
        \sha1_round/add_79_3/n217 ) );
  INV_X1 \sha1_round/add_79_3/U114  ( .A(\sha1_round/N263 ), .ZN(
        \sha1_round/add_79_3/n17 ) );
  INV_X4 \sha1_round/add_79_3/U113  ( .A(\sha1_round/N266 ), .ZN(
        \sha1_round/add_79_3/n332 ) );
  AND2_X2 \sha1_round/add_79_3/U112  ( .A1(\sha1_round/add_79_3/n298 ), .A2(
        \sha1_round/add_79_3/n299 ), .ZN(\sha1_round/add_79_3/n22 ) );
  NAND2_X1 \sha1_round/add_79_3/U111  ( .A1(\sha1_round/N293 ), .A2(
        \sha1_round/N261 ), .ZN(\sha1_round/add_79_3/n74 ) );
  NAND2_X1 \sha1_round/add_79_3/U110  ( .A1(\sha1_round/add_79_3/n73 ), .A2(
        \sha1_round/add_79_3/n77 ), .ZN(\sha1_round/add_79_3/n366 ) );
  INV_X4 \sha1_round/add_79_3/U109  ( .A(\sha1_round/add_79_3/n163 ), .ZN(
        \sha1_round/add_79_3/n162 ) );
  NAND4_X1 \sha1_round/add_79_3/U108  ( .A1(\sha1_round/add_79_3/n342 ), .A2(
        \sha1_round/add_79_3/n343 ), .A3(\sha1_round/add_79_3/n299 ), .A4(
        \sha1_round/add_79_3/n101 ), .ZN(\sha1_round/add_79_3/n338 ) );
  NAND3_X1 \sha1_round/add_79_3/U107  ( .A1(\sha1_round/add_79_3/n81 ), .A2(
        \sha1_round/add_79_3/n343 ), .A3(\sha1_round/add_79_3/n299 ), .ZN(
        \sha1_round/add_79_3/n339 ) );
  INV_X1 \sha1_round/add_79_3/U106  ( .A(\sha1_round/add_79_3/n303 ), .ZN(
        \sha1_round/add_79_3/n343 ) );
  NOR2_X1 \sha1_round/add_79_3/U105  ( .A1(\sha1_round/add_79_3/n349 ), .A2(
        \sha1_round/add_79_3/n303 ), .ZN(\sha1_round/add_79_3/n345 ) );
  NAND2_X2 \sha1_round/add_79_3/U104  ( .A1(\sha1_round/add_79_3/n173 ), .A2(
        \sha1_round/add_79_3/n174 ), .ZN(\sha1_round/add_79_3/n172 ) );
  XNOR2_X1 \sha1_round/add_79_3/U103  ( .A(\sha1_round/add_79_3/n334 ), .B(
        \sha1_round/add_79_3/n335 ), .ZN(\sha1_round/N329 ) );
  NAND2_X2 \sha1_round/add_79_3/U102  ( .A1(\sha1_round/add_79_3/n142 ), .A2(
        \sha1_round/add_79_3/n134 ), .ZN(\sha1_round/add_79_3/n140 ) );
  INV_X4 \sha1_round/add_79_3/U101  ( .A(\sha1_round/N265 ), .ZN(
        \sha1_round/add_79_3/n337 ) );
  NAND2_X2 \sha1_round/add_79_3/U100  ( .A1(\sha1_round/N296 ), .A2(
        \sha1_round/N264 ), .ZN(\sha1_round/add_79_3/n301 ) );
  NOR2_X2 \sha1_round/add_79_3/U99  ( .A1(\sha1_round/add_79_3/n257 ), .A2(
        \sha1_round/add_79_3/n280 ), .ZN(\sha1_round/add_79_3/n279 ) );
  NOR2_X2 \sha1_round/add_79_3/U98  ( .A1(\sha1_round/N270 ), .A2(
        \sha1_round/N302 ), .ZN(\sha1_round/add_79_3/n257 ) );
  NOR2_X2 \sha1_round/add_79_3/U97  ( .A1(\sha1_round/N270 ), .A2(
        \sha1_round/N302 ), .ZN(\sha1_round/add_79_3/n275 ) );
  OR2_X4 \sha1_round/add_79_3/U96  ( .A1(\sha1_round/add_79_3/n382 ), .A2(
        \sha1_round/add_79_3/n88 ), .ZN(\sha1_round/add_79_3/n16 ) );
  NAND2_X2 \sha1_round/add_79_3/U95  ( .A1(\sha1_round/add_79_3/n296 ), .A2(
        \sha1_round/add_79_3/n237 ), .ZN(\sha1_round/add_79_3/n295 ) );
  AND2_X4 \sha1_round/add_79_3/U94  ( .A1(\sha1_round/add_79_3/n239 ), .A2(
        \sha1_round/add_79_3/n5 ), .ZN(\sha1_round/add_79_3/n15 ) );
  INV_X4 \sha1_round/add_79_3/U93  ( .A(\sha1_round/add_79_3/n355 ), .ZN(
        \sha1_round/add_79_3/n354 ) );
  AND2_X4 \sha1_round/add_79_3/U92  ( .A1(\sha1_round/add_79_3/n378 ), .A2(
        \sha1_round/add_79_3/n379 ), .ZN(\sha1_round/add_79_3/n14 ) );
  OR2_X4 \sha1_round/add_79_3/U91  ( .A1(\sha1_round/add_79_3/n107 ), .A2(
        \sha1_round/add_79_3/n313 ), .ZN(\sha1_round/add_79_3/n13 ) );
  AND2_X4 \sha1_round/add_79_3/U90  ( .A1(\sha1_round/add_79_3/n301 ), .A2(
        \sha1_round/add_79_3/n302 ), .ZN(\sha1_round/add_79_3/n12 ) );
  AND2_X4 \sha1_round/add_79_3/U89  ( .A1(\sha1_round/add_79_3/n256 ), .A2(
        \sha1_round/add_79_3/n251 ), .ZN(\sha1_round/add_79_3/n11 ) );
  AND2_X4 \sha1_round/add_79_3/U88  ( .A1(\sha1_round/add_79_3/n179 ), .A2(
        \sha1_round/add_79_3/n177 ), .ZN(\sha1_round/add_79_3/n10 ) );
  NOR2_X2 \sha1_round/add_79_3/U87  ( .A1(\sha1_round/N272 ), .A2(
        \sha1_round/N304 ), .ZN(\sha1_round/add_79_3/n218 ) );
  NAND2_X2 \sha1_round/add_79_3/U86  ( .A1(\sha1_round/add_79_3/n199 ), .A2(
        \sha1_round/add_79_3/n150 ), .ZN(\sha1_round/add_79_3/n165 ) );
  AND4_X4 \sha1_round/add_79_3/U85  ( .A1(\sha1_round/add_79_3/n315 ), .A2(
        \sha1_round/add_79_3/n316 ), .A3(\sha1_round/add_79_3/n317 ), .A4(
        \sha1_round/add_79_3/n318 ), .ZN(\sha1_round/add_79_3/n9 ) );
  NOR2_X2 \sha1_round/add_79_3/U84  ( .A1(\sha1_round/N256 ), .A2(
        \sha1_round/N288 ), .ZN(\sha1_round/add_79_3/n102 ) );
  NOR2_X2 \sha1_round/add_79_3/U83  ( .A1(\sha1_round/N254 ), .A2(
        \sha1_round/N286 ), .ZN(\sha1_round/add_79_3/n111 ) );
  INV_X4 \sha1_round/add_79_3/U82  ( .A(\sha1_round/N263 ), .ZN(
        \sha1_round/add_79_3/n357 ) );
  AND2_X4 \sha1_round/add_79_3/U81  ( .A1(\sha1_round/add_79_3/n271 ), .A2(
        \sha1_round/add_79_3/n274 ), .ZN(\sha1_round/add_79_3/n8 ) );
  AND2_X4 \sha1_round/add_79_3/U80  ( .A1(\sha1_round/add_79_3/n273 ), .A2(
        \sha1_round/add_79_3/n274 ), .ZN(\sha1_round/add_79_3/n7 ) );
  OR2_X4 \sha1_round/add_79_3/U79  ( .A1(\sha1_round/add_79_3/n283 ), .A2(
        \sha1_round/add_79_3/n276 ), .ZN(\sha1_round/add_79_3/n6 ) );
  AND2_X4 \sha1_round/add_79_3/U78  ( .A1(\sha1_round/add_79_3/n302 ), .A2(
        \sha1_round/add_79_3/n301 ), .ZN(\sha1_round/add_79_3/n5 ) );
  INV_X2 \sha1_round/add_79_3/U77  ( .A(\sha1_round/add_79_3/n247 ), .ZN(
        \sha1_round/add_79_3/n290 ) );
  NOR2_X2 \sha1_round/add_79_3/U76  ( .A1(\sha1_round/add_79_3/n102 ), .A2(
        \sha1_round/add_79_3/n96 ), .ZN(\sha1_round/add_79_3/n379 ) );
  NOR2_X2 \sha1_round/add_79_3/U75  ( .A1(\sha1_round/add_79_3/n96 ), .A2(
        \sha1_round/add_79_3/n385 ), .ZN(\sha1_round/add_79_3/n384 ) );
  NAND2_X2 \sha1_round/add_79_3/U74  ( .A1(\sha1_round/add_79_3/n143 ), .A2(
        \sha1_round/add_79_3/n138 ), .ZN(\sha1_round/add_79_3/n142 ) );
  NAND2_X2 \sha1_round/add_79_3/U73  ( .A1(\sha1_round/N263 ), .A2(
        \sha1_round/N295 ), .ZN(\sha1_round/add_79_3/n302 ) );
  NAND3_X4 \sha1_round/add_79_3/U72  ( .A1(\sha1_round/add_79_3/n244 ), .A2(
        \sha1_round/add_79_3/n245 ), .A3(\sha1_round/add_79_3/n246 ), .ZN(
        \sha1_round/add_79_3/n241 ) );
  NAND2_X4 \sha1_round/add_79_3/U71  ( .A1(\sha1_round/add_79_3/n329 ), .A2(
        \sha1_round/add_79_3/n297 ), .ZN(\sha1_round/add_79_3/n328 ) );
  NAND2_X2 \sha1_round/add_79_3/U70  ( .A1(\sha1_round/add_79_3/n149 ), .A2(
        \sha1_round/add_79_3/n65 ), .ZN(\sha1_round/add_79_3/n126 ) );
  NAND2_X2 \sha1_round/add_79_3/U69  ( .A1(\sha1_round/add_79_3/n195 ), .A2(
        \sha1_round/add_79_3/n196 ), .ZN(\sha1_round/add_79_3/n178 ) );
  NAND2_X2 \sha1_round/add_79_3/U68  ( .A1(\sha1_round/add_79_3/n213 ), .A2(
        \sha1_round/add_79_3/n214 ), .ZN(\sha1_round/add_79_3/n200 ) );
  INV_X4 \sha1_round/add_79_3/U67  ( .A(\sha1_round/add_79_3/n278 ), .ZN(
        \sha1_round/add_79_3/n46 ) );
  NAND2_X2 \sha1_round/add_79_3/U66  ( .A1(\sha1_round/add_79_3/n98 ), .A2(
        \sha1_round/add_79_3/n99 ), .ZN(\sha1_round/add_79_3/n94 ) );
  NAND2_X2 \sha1_round/add_79_3/U65  ( .A1(\sha1_round/N292 ), .A2(
        \sha1_round/N260 ), .ZN(\sha1_round/add_79_3/n76 ) );
  NOR2_X2 \sha1_round/add_79_3/U64  ( .A1(\sha1_round/add_79_3/n147 ), .A2(
        \sha1_round/add_79_3/n120 ), .ZN(\sha1_round/add_79_3/n56 ) );
  NOR3_X2 \sha1_round/add_79_3/U63  ( .A1(\sha1_round/add_79_3/n241 ), .A2(
        \sha1_round/add_79_3/n4 ), .A3(\sha1_round/add_79_3/n243 ), .ZN(
        \sha1_round/add_79_3/n238 ) );
  INV_X4 \sha1_round/add_79_3/U62  ( .A(\sha1_round/add_79_3/n53 ), .ZN(
        \sha1_round/add_79_3/n54 ) );
  NOR2_X2 \sha1_round/add_79_3/U61  ( .A1(\sha1_round/add_79_3/n235 ), .A2(
        \sha1_round/add_79_3/n54 ), .ZN(\sha1_round/add_79_3/n234 ) );
  NAND2_X2 \sha1_round/add_79_3/U60  ( .A1(\sha1_round/add_79_3/n11 ), .A2(
        \sha1_round/add_79_3/n282 ), .ZN(\sha1_round/add_79_3/n255 ) );
  NAND2_X2 \sha1_round/add_79_3/U59  ( .A1(\sha1_round/add_79_3/n255 ), .A2(
        \sha1_round/add_79_3/n254 ), .ZN(\sha1_round/add_79_3/n253 ) );
  INV_X4 \sha1_round/add_79_3/U58  ( .A(\sha1_round/add_79_3/n77 ), .ZN(
        \sha1_round/add_79_3/n319 ) );
  NOR2_X2 \sha1_round/add_79_3/U57  ( .A1(\sha1_round/add_79_3/n217 ), .A2(
        \sha1_round/add_79_3/n218 ), .ZN(\sha1_round/add_79_3/n207 ) );
  NOR2_X2 \sha1_round/add_79_3/U56  ( .A1(\sha1_round/add_79_3/n175 ), .A2(
        \sha1_round/add_79_3/n176 ), .ZN(\sha1_round/add_79_3/n171 ) );
  NAND2_X2 \sha1_round/add_79_3/U55  ( .A1(\sha1_round/add_79_3/n171 ), .A2(
        \sha1_round/add_79_3/n172 ), .ZN(\sha1_round/add_79_3/n159 ) );
  NAND2_X2 \sha1_round/add_79_3/U54  ( .A1(\sha1_round/add_79_3/n162 ), .A2(
        \sha1_round/add_79_3/n158 ), .ZN(\sha1_round/add_79_3/n153 ) );
  NOR2_X2 \sha1_round/add_79_3/U53  ( .A1(\sha1_round/add_79_3/n4 ), .A2(
        \sha1_round/add_79_3/n300 ), .ZN(\sha1_round/add_79_3/n235 ) );
  INV_X4 \sha1_round/add_79_3/U52  ( .A(\sha1_round/add_79_3/n19 ), .ZN(
        \sha1_round/add_79_3/n322 ) );
  NAND2_X2 \sha1_round/add_79_3/U51  ( .A1(\sha1_round/add_79_3/n207 ), .A2(
        \sha1_round/add_79_3/n200 ), .ZN(\sha1_round/add_79_3/n198 ) );
  NOR2_X2 \sha1_round/add_79_3/U50  ( .A1(\sha1_round/add_79_3/n386 ), .A2(
        \sha1_round/add_79_3/n387 ), .ZN(\sha1_round/add_79_3/n383 ) );
  INV_X4 \sha1_round/add_79_3/U49  ( .A(\sha1_round/add_79_3/n16 ), .ZN(
        \sha1_round/add_79_3/n243 ) );
  AND2_X4 \sha1_round/add_79_3/U48  ( .A1(\sha1_round/add_79_3/n371 ), .A2(
        \sha1_round/add_79_3/n370 ), .ZN(\sha1_round/add_79_3/n369 ) );
  NAND2_X4 \sha1_round/add_79_3/U47  ( .A1(\sha1_round/add_79_3/n226 ), .A2(
        \sha1_round/add_79_3/n227 ), .ZN(\sha1_round/add_79_3/n222 ) );
  NOR2_X4 \sha1_round/add_79_3/U46  ( .A1(\sha1_round/add_79_3/n87 ), .A2(
        \sha1_round/add_79_3/n323 ), .ZN(\sha1_round/add_79_3/n380 ) );
  NOR2_X4 \sha1_round/add_79_3/U45  ( .A1(\sha1_round/add_79_3/n288 ), .A2(
        \sha1_round/add_79_3/n6 ), .ZN(\sha1_round/add_79_3/n281 ) );
  NOR2_X4 \sha1_round/add_79_3/U44  ( .A1(\sha1_round/add_79_3/n281 ), .A2(
        \sha1_round/add_79_3/n282 ), .ZN(\sha1_round/add_79_3/n278 ) );
  NAND2_X4 \sha1_round/add_79_3/U43  ( .A1(\sha1_round/add_79_3/n7 ), .A2(
        \sha1_round/add_79_3/n251 ), .ZN(\sha1_round/add_79_3/n236 ) );
  INV_X4 \sha1_round/add_79_3/U42  ( .A(\sha1_round/add_79_3/n236 ), .ZN(
        \sha1_round/add_79_3/n248 ) );
  INV_X1 \sha1_round/add_79_3/U41  ( .A(\sha1_round/add_79_3/n210 ), .ZN(
        \sha1_round/add_79_3/n221 ) );
  NAND2_X4 \sha1_round/add_79_3/U40  ( .A1(\sha1_round/add_79_3/n357 ), .A2(
        \sha1_round/add_79_3/n356 ), .ZN(\sha1_round/add_79_3/n19 ) );
  NAND2_X2 \sha1_round/add_79_3/U39  ( .A1(\sha1_round/add_79_3/n34 ), .A2(
        \sha1_round/add_79_3/n35 ), .ZN(\sha1_round/add_79_3/n37 ) );
  NAND2_X2 \sha1_round/add_79_3/U38  ( .A1(\sha1_round/add_79_3/n294 ), .A2(
        \sha1_round/add_79_3/n333 ), .ZN(\sha1_round/add_79_3/n329 ) );
  NOR2_X2 \sha1_round/add_79_3/U37  ( .A1(\sha1_round/add_79_3/n360 ), .A2(
        \sha1_round/add_79_3/n321 ), .ZN(\sha1_round/add_79_3/n358 ) );
  INV_X4 \sha1_round/add_79_3/U36  ( .A(\sha1_round/add_79_3/n350 ), .ZN(
        \sha1_round/add_79_3/n321 ) );
  NAND2_X2 \sha1_round/add_79_3/U35  ( .A1(\sha1_round/add_79_3/n170 ), .A2(
        \sha1_round/add_79_3/n158 ), .ZN(\sha1_round/add_79_3/n156 ) );
  NAND2_X2 \sha1_round/add_79_3/U34  ( .A1(\sha1_round/add_79_3/n156 ), .A2(
        \sha1_round/add_79_3/n157 ), .ZN(\sha1_round/add_79_3/n154 ) );
  NOR2_X2 \sha1_round/add_79_3/U33  ( .A1(\sha1_round/add_79_3/n161 ), .A2(
        \sha1_round/add_79_3/n153 ), .ZN(\sha1_round/add_79_3/n155 ) );
  NAND2_X2 \sha1_round/add_79_3/U32  ( .A1(\sha1_round/add_79_3/n191 ), .A2(
        \sha1_round/add_79_3/n192 ), .ZN(\sha1_round/add_79_3/n179 ) );
  NAND2_X2 \sha1_round/add_79_3/U31  ( .A1(\sha1_round/add_79_3/n9 ), .A2(
        \sha1_round/add_79_3/n240 ), .ZN(\sha1_round/add_79_3/n305 ) );
  NOR2_X4 \sha1_round/add_79_3/U30  ( .A1(\sha1_round/N258 ), .A2(
        \sha1_round/N290 ), .ZN(\sha1_round/add_79_3/n90 ) );
  NOR2_X1 \sha1_round/add_79_3/U29  ( .A1(\sha1_round/add_79_3/n90 ), .A2(
        \sha1_round/add_79_3/n88 ), .ZN(\sha1_round/add_79_3/n317 ) );
  INV_X8 \sha1_round/add_79_3/U28  ( .A(\sha1_round/add_79_3/n90 ), .ZN(
        \sha1_round/add_79_3/n378 ) );
  NAND2_X4 \sha1_round/add_79_3/U27  ( .A1(\sha1_round/add_79_3/n369 ), .A2(
        \sha1_round/add_79_3/n309 ), .ZN(\sha1_round/add_79_3/n101 ) );
  NAND2_X4 \sha1_round/add_79_3/U26  ( .A1(\sha1_round/add_79_3/n100 ), .A2(
        \sha1_round/add_79_3/n101 ), .ZN(\sha1_round/add_79_3/n99 ) );
  XNOR2_X1 \sha1_round/add_79_3/U25  ( .A(\sha1_round/add_79_3/n103 ), .B(
        \sha1_round/add_79_3/n101 ), .ZN(\sha1_round/N320 ) );
  NAND2_X4 \sha1_round/add_79_3/U24  ( .A1(\sha1_round/add_79_3/n342 ), .A2(
        \sha1_round/add_79_3/n101 ), .ZN(\sha1_round/add_79_3/n80 ) );
  NAND2_X4 \sha1_round/add_79_3/U23  ( .A1(\sha1_round/add_79_3/n367 ), .A2(
        \sha1_round/add_79_3/n368 ), .ZN(\sha1_round/add_79_3/n73 ) );
  INV_X8 \sha1_round/add_79_3/U22  ( .A(\sha1_round/add_79_3/n73 ), .ZN(
        \sha1_round/add_79_3/n320 ) );
  NOR2_X4 \sha1_round/add_79_3/U21  ( .A1(\sha1_round/N257 ), .A2(
        \sha1_round/N289 ), .ZN(\sha1_round/add_79_3/n96 ) );
  NAND2_X1 \sha1_round/add_79_3/U20  ( .A1(\sha1_round/N289 ), .A2(
        \sha1_round/N257 ), .ZN(\sha1_round/add_79_3/n93 ) );
  NAND2_X4 \sha1_round/add_79_3/U19  ( .A1(\sha1_round/add_79_3/n187 ), .A2(
        \sha1_round/add_79_3/n180 ), .ZN(\sha1_round/add_79_3/n186 ) );
  NOR2_X2 \sha1_round/add_79_3/U18  ( .A1(\sha1_round/add_79_3/n155 ), .A2(
        \sha1_round/add_79_3/n154 ), .ZN(\sha1_round/add_79_3/n51 ) );
  NOR2_X4 \sha1_round/add_79_3/U17  ( .A1(\sha1_round/add_79_3/n358 ), .A2(
        \sha1_round/add_79_3/n359 ), .ZN(\sha1_round/add_79_3/n353 ) );
  INV_X8 \sha1_round/add_79_3/U16  ( .A(\sha1_round/add_79_3/n3 ), .ZN(
        \sha1_round/add_79_3/n4 ) );
  INV_X4 \sha1_round/add_79_3/U15  ( .A(\sha1_round/add_79_3/n242 ), .ZN(
        \sha1_round/add_79_3/n3 ) );
  NAND4_X4 \sha1_round/add_79_3/U14  ( .A1(\sha1_round/add_79_3/n338 ), .A2(
        \sha1_round/add_79_3/n339 ), .A3(\sha1_round/add_79_3/n301 ), .A4(
        \sha1_round/add_79_3/n340 ), .ZN(\sha1_round/add_79_3/n334 ) );
  NAND2_X4 \sha1_round/add_79_3/U13  ( .A1(\sha1_round/add_79_3/n334 ), .A2(
        \sha1_round/add_79_3/n52 ), .ZN(\sha1_round/add_79_3/n333 ) );
  NAND2_X4 \sha1_round/add_79_3/U12  ( .A1(\sha1_round/add_79_3/n193 ), .A2(
        \sha1_round/add_79_3/n174 ), .ZN(\sha1_round/add_79_3/n189 ) );
  NAND2_X4 \sha1_round/add_79_3/U11  ( .A1(\sha1_round/add_79_3/n36 ), .A2(
        \sha1_round/add_79_3/n37 ), .ZN(\sha1_round/N342 ) );
  NOR2_X4 \sha1_round/add_79_3/U10  ( .A1(\sha1_round/add_79_3/n236 ), .A2(
        \sha1_round/add_79_3/n21 ), .ZN(\sha1_round/add_79_3/n53 ) );
  NAND2_X4 \sha1_round/add_79_3/U9  ( .A1(\sha1_round/add_79_3/n363 ), .A2(
        \sha1_round/add_79_3/n362 ), .ZN(\sha1_round/add_79_3/n350 ) );
  NAND2_X4 \sha1_round/add_79_3/U8  ( .A1(\sha1_round/add_79_3/n224 ), .A2(
        \sha1_round/add_79_3/n225 ), .ZN(\sha1_round/add_79_3/n219 ) );
  NAND2_X4 \sha1_round/add_79_3/U7  ( .A1(\sha1_round/add_79_3/n154 ), .A2(
        \sha1_round/add_79_3/n152 ), .ZN(\sha1_round/add_79_3/n129 ) );
  NAND2_X4 \sha1_round/add_79_3/U6  ( .A1(\sha1_round/add_79_3/n159 ), .A2(
        \sha1_round/add_79_3/n160 ), .ZN(\sha1_round/add_79_3/n170 ) );
  XNOR2_X1 \sha1_round/add_79_3/U5  ( .A(\sha1_round/add_79_3/n229 ), .B(
        \sha1_round/add_79_3/n148 ), .ZN(\sha1_round/N336 ) );
  AND2_X4 \sha1_round/add_79_3/U4  ( .A1(\sha1_round/add_79_3/n136 ), .A2(
        \sha1_round/add_79_3/n152 ), .ZN(\sha1_round/add_79_3/n1 ) );
  NAND2_X2 \sha1_round/add_79_3/U3  ( .A1(\sha1_round/add_79_3/n270 ), .A2(
        \sha1_round/add_79_3/n271 ), .ZN(\sha1_round/add_79_3/n282 ) );
  NOR2_X4 \sha1_round/add_79_3/U2  ( .A1(\sha1_round/add_79_3/n169 ), .A2(
        \sha1_round/add_79_3/n170 ), .ZN(\sha1_round/add_79_3/n168 ) );
  NAND2_X2 \sha1_round/add_79/U405  ( .A1(\sha1_round/k_23 ), .A2(
        \sha1_round/f [0]), .ZN(\sha1_round/add_79/n270 ) );
  NOR2_X4 \sha1_round/add_79/U404  ( .A1(\sha1_round/add_79/n377 ), .A2(
        \sha1_round/add_79/n83 ), .ZN(\sha1_round/add_79/n376 ) );
  NAND3_X4 \sha1_round/add_79/U403  ( .A1(\sha1_round/add_79/n374 ), .A2(
        \sha1_round/add_79/n375 ), .A3(\sha1_round/add_79/n376 ), .ZN(
        \sha1_round/add_79/n109 ) );
  INV_X4 \sha1_round/add_79/U402  ( .A(\sha1_round/add_79/n380 ), .ZN(
        \sha1_round/add_79/n121 ) );
  INV_X4 \sha1_round/add_79/U401  ( .A(\sha1_round/add_79/n306 ), .ZN(
        \sha1_round/add_79/n129 ) );
  INV_X4 \sha1_round/add_79/U400  ( .A(\sha1_round/k[13] ), .ZN(
        \sha1_round/add_79/n354 ) );
  INV_X4 \sha1_round/add_79/U399  ( .A(\sha1_round/f [11]), .ZN(
        \sha1_round/add_79/n355 ) );
  INV_X4 \sha1_round/add_79/U398  ( .A(\sha1_round/add_79/n343 ), .ZN(
        \sha1_round/add_79/n345 ) );
  XNOR2_X2 \sha1_round/add_79/U397  ( .A(\sha1_round/add_79/n352 ), .B(
        \sha1_round/add_79/n353 ), .ZN(\sha1_round/add_79/n351 ) );
  INV_X4 \sha1_round/add_79/U396  ( .A(\sha1_round/f [12]), .ZN(
        \sha1_round/add_79/n350 ) );
  NAND2_X2 \sha1_round/add_79/U395  ( .A1(\sha1_round/add_79/n92 ), .A2(
        \sha1_round/add_79/n350 ), .ZN(\sha1_round/add_79/n313 ) );
  NAND2_X2 \sha1_round/add_79/U394  ( .A1(\sha1_round/add_79/n313 ), .A2(
        \sha1_round/add_79/n302 ), .ZN(\sha1_round/add_79/n337 ) );
  NAND2_X2 \sha1_round/add_79/U393  ( .A1(\sha1_round/k_30 ), .A2(
        \sha1_round/f [8]), .ZN(\sha1_round/add_79/n341 ) );
  NAND4_X2 \sha1_round/add_79/U392  ( .A1(\sha1_round/add_79/n341 ), .A2(
        \sha1_round/add_79/n342 ), .A3(\sha1_round/add_79/n343 ), .A4(
        \sha1_round/add_79/n344 ), .ZN(\sha1_round/add_79/n339 ) );
  XNOR2_X2 \sha1_round/add_79/U391  ( .A(\sha1_round/add_79/n336 ), .B(
        \sha1_round/add_79/n337 ), .ZN(\sha1_round/N264 ) );
  INV_X4 \sha1_round/add_79/U390  ( .A(\sha1_round/add_79/n323 ), .ZN(
        \sha1_round/add_79/n334 ) );
  XNOR2_X2 \sha1_round/add_79/U389  ( .A(\sha1_round/add_79/n333 ), .B(
        \sha1_round/add_79/n20 ), .ZN(\sha1_round/N265 ) );
  INV_X4 \sha1_round/add_79/U388  ( .A(\sha1_round/add_79/n313 ), .ZN(
        \sha1_round/add_79/n330 ) );
  NAND2_X2 \sha1_round/add_79/U387  ( .A1(\sha1_round/add_79/n294 ), .A2(
        \sha1_round/add_79/n327 ), .ZN(\sha1_round/add_79/n326 ) );
  NAND2_X2 \sha1_round/add_79/U386  ( .A1(\sha1_round/k[15] ), .A2(
        \sha1_round/f [15]), .ZN(\sha1_round/add_79/n295 ) );
  INV_X4 \sha1_round/add_79/U385  ( .A(\sha1_round/add_79/n318 ), .ZN(
        \sha1_round/add_79/n314 ) );
  INV_X4 \sha1_round/add_79/U384  ( .A(\sha1_round/add_79/n289 ), .ZN(
        \sha1_round/add_79/n316 ) );
  INV_X4 \sha1_round/add_79/U383  ( .A(\sha1_round/add_79/n238 ), .ZN(
        \sha1_round/add_79/n297 ) );
  NAND3_X2 \sha1_round/add_79/U382  ( .A1(\sha1_round/add_79/n70 ), .A2(
        \sha1_round/add_79/n306 ), .A3(\sha1_round/add_79/n307 ), .ZN(
        \sha1_round/add_79/n305 ) );
  NAND2_X2 \sha1_round/add_79/U381  ( .A1(\sha1_round/add_79/n304 ), .A2(
        \sha1_round/add_79/n305 ), .ZN(\sha1_round/add_79/n298 ) );
  INV_X4 \sha1_round/add_79/U380  ( .A(\sha1_round/add_79/n303 ), .ZN(
        \sha1_round/add_79/n300 ) );
  INV_X4 \sha1_round/add_79/U379  ( .A(\sha1_round/add_79/n302 ), .ZN(
        \sha1_round/add_79/n301 ) );
  NAND2_X2 \sha1_round/add_79/U378  ( .A1(\sha1_round/k[13] ), .A2(
        \sha1_round/f [13]), .ZN(\sha1_round/add_79/n296 ) );
  INV_X4 \sha1_round/add_79/U377  ( .A(\sha1_round/k_26 ), .ZN(
        \sha1_round/add_79/n201 ) );
  INV_X4 \sha1_round/add_79/U376  ( .A(\sha1_round/f [16]), .ZN(
        \sha1_round/add_79/n292 ) );
  NAND2_X2 \sha1_round/add_79/U375  ( .A1(\sha1_round/add_79/n201 ), .A2(
        \sha1_round/add_79/n292 ), .ZN(\sha1_round/add_79/n280 ) );
  NAND2_X2 \sha1_round/add_79/U374  ( .A1(\sha1_round/add_79/n293 ), .A2(
        \sha1_round/add_79/n233 ), .ZN(\sha1_round/add_79/n279 ) );
  NAND2_X2 \sha1_round/add_79/U373  ( .A1(\sha1_round/add_79/n279 ), .A2(
        \sha1_round/add_79/n280 ), .ZN(\sha1_round/add_79/n284 ) );
  INV_X4 \sha1_round/add_79/U372  ( .A(\sha1_round/add_79/n275 ), .ZN(
        \sha1_round/add_79/n239 ) );
  INV_X4 \sha1_round/add_79/U371  ( .A(\sha1_round/add_79/n280 ), .ZN(
        \sha1_round/add_79/n278 ) );
  NAND2_X2 \sha1_round/add_79/U370  ( .A1(\sha1_round/add_79/n231 ), .A2(
        \sha1_round/add_79/n279 ), .ZN(\sha1_round/add_79/n274 ) );
  XNOR2_X2 \sha1_round/add_79/U369  ( .A(\sha1_round/add_79/n250 ), .B(
        \sha1_round/add_79/n262 ), .ZN(\sha1_round/N270 ) );
  INV_X4 \sha1_round/add_79/U368  ( .A(\sha1_round/add_79/n266 ), .ZN(
        \sha1_round/add_79/n272 ) );
  XNOR2_X2 \sha1_round/add_79/U367  ( .A(\sha1_round/add_79/n270 ), .B(
        \sha1_round/add_79/n268 ), .ZN(\sha1_round/N253 ) );
  INV_X4 \sha1_round/add_79/U366  ( .A(\sha1_round/f [20]), .ZN(
        \sha1_round/add_79/n265 ) );
  NAND2_X2 \sha1_round/add_79/U365  ( .A1(\sha1_round/add_79/n201 ), .A2(
        \sha1_round/add_79/n265 ), .ZN(\sha1_round/add_79/n259 ) );
  NAND2_X2 \sha1_round/add_79/U364  ( .A1(\sha1_round/add_79/n258 ), .A2(
        \sha1_round/add_79/n259 ), .ZN(\sha1_round/add_79/n264 ) );
  NAND2_X2 \sha1_round/add_79/U363  ( .A1(\sha1_round/f [19]), .A2(
        \sha1_round/k_26 ), .ZN(\sha1_round/add_79/n257 ) );
  XNOR2_X2 \sha1_round/add_79/U362  ( .A(\sha1_round/add_79/n254 ), .B(
        \sha1_round/add_79/n15 ), .ZN(\sha1_round/N273 ) );
  INV_X4 \sha1_round/add_79/U361  ( .A(\sha1_round/add_79/n240 ), .ZN(
        \sha1_round/add_79/n253 ) );
  INV_X4 \sha1_round/add_79/U360  ( .A(\sha1_round/add_79/n251 ), .ZN(
        \sha1_round/add_79/n242 ) );
  NAND2_X2 \sha1_round/add_79/U359  ( .A1(\sha1_round/add_79/n248 ), .A2(
        \sha1_round/add_79/n249 ), .ZN(\sha1_round/add_79/n245 ) );
  INV_X4 \sha1_round/add_79/U358  ( .A(\sha1_round/f [22]), .ZN(
        \sha1_round/add_79/n247 ) );
  NAND2_X2 \sha1_round/add_79/U357  ( .A1(\sha1_round/add_79/n91 ), .A2(
        \sha1_round/add_79/n247 ), .ZN(\sha1_round/add_79/n241 ) );
  NAND2_X2 \sha1_round/add_79/U356  ( .A1(\sha1_round/n3370 ), .A2(
        \sha1_round/f [22]), .ZN(\sha1_round/add_79/n243 ) );
  NAND2_X2 \sha1_round/add_79/U355  ( .A1(\sha1_round/add_79/n241 ), .A2(
        \sha1_round/add_79/n243 ), .ZN(\sha1_round/add_79/n246 ) );
  NAND2_X2 \sha1_round/add_79/U354  ( .A1(\sha1_round/add_79/n219 ), .A2(
        \sha1_round/add_79/n222 ), .ZN(\sha1_round/add_79/n228 ) );
  INV_X4 \sha1_round/add_79/U353  ( .A(\sha1_round/add_79/n243 ), .ZN(
        \sha1_round/add_79/n227 ) );
  INV_X4 \sha1_round/add_79/U352  ( .A(\sha1_round/add_79/n237 ), .ZN(
        \sha1_round/add_79/n230 ) );
  INV_X4 \sha1_round/add_79/U351  ( .A(\sha1_round/add_79/n213 ), .ZN(
        \sha1_round/add_79/n222 ) );
  NAND2_X2 \sha1_round/add_79/U350  ( .A1(\sha1_round/add_79/n221 ), .A2(
        \sha1_round/add_79/n222 ), .ZN(\sha1_round/add_79/n220 ) );
  NAND2_X2 \sha1_round/add_79/U349  ( .A1(\sha1_round/add_79/n219 ), .A2(
        \sha1_round/add_79/n220 ), .ZN(\sha1_round/add_79/n217 ) );
  NAND2_X2 \sha1_round/add_79/U348  ( .A1(\sha1_round/f [24]), .A2(
        \sha1_round/add_79/n89 ), .ZN(\sha1_round/add_79/n196 ) );
  XNOR2_X2 \sha1_round/add_79/U347  ( .A(\sha1_round/add_79/n217 ), .B(
        \sha1_round/add_79/n218 ), .ZN(\sha1_round/add_79/n216 ) );
  INV_X4 \sha1_round/add_79/U346  ( .A(\sha1_round/add_79/n216 ), .ZN(
        \sha1_round/N276 ) );
  INV_X4 \sha1_round/add_79/U345  ( .A(\sha1_round/add_79/n196 ), .ZN(
        \sha1_round/add_79/n214 ) );
  INV_X4 \sha1_round/add_79/U344  ( .A(\sha1_round/add_79/n197 ), .ZN(
        \sha1_round/add_79/n215 ) );
  INV_X4 \sha1_round/add_79/U343  ( .A(\sha1_round/f [25]), .ZN(
        \sha1_round/add_79/n209 ) );
  NAND2_X2 \sha1_round/add_79/U342  ( .A1(\sha1_round/add_79/n55 ), .A2(
        \sha1_round/add_79/n209 ), .ZN(\sha1_round/add_79/n193 ) );
  NAND2_X2 \sha1_round/add_79/U341  ( .A1(\sha1_round/add_79/n193 ), .A2(
        \sha1_round/add_79/n198 ), .ZN(\sha1_round/add_79/n208 ) );
  XNOR2_X2 \sha1_round/add_79/U340  ( .A(\sha1_round/add_79/n207 ), .B(
        \sha1_round/add_79/n208 ), .ZN(\sha1_round/N277 ) );
  NAND2_X2 \sha1_round/add_79/U339  ( .A1(\sha1_round/add_79/n206 ), .A2(
        \sha1_round/add_79/n193 ), .ZN(\sha1_round/add_79/n203 ) );
  NAND2_X2 \sha1_round/add_79/U338  ( .A1(\sha1_round/f [26]), .A2(
        \sha1_round/k_26 ), .ZN(\sha1_round/add_79/n192 ) );
  INV_X4 \sha1_round/add_79/U337  ( .A(\sha1_round/f [26]), .ZN(
        \sha1_round/add_79/n202 ) );
  NAND2_X2 \sha1_round/add_79/U336  ( .A1(\sha1_round/add_79/n201 ), .A2(
        \sha1_round/add_79/n202 ), .ZN(\sha1_round/add_79/n194 ) );
  NAND2_X2 \sha1_round/add_79/U335  ( .A1(\sha1_round/add_79/n192 ), .A2(
        \sha1_round/add_79/n194 ), .ZN(\sha1_round/add_79/n200 ) );
  XNOR2_X2 \sha1_round/add_79/U334  ( .A(\sha1_round/add_79/n199 ), .B(
        \sha1_round/add_79/n200 ), .ZN(\sha1_round/N278 ) );
  NAND2_X2 \sha1_round/add_79/U333  ( .A1(\sha1_round/add_79/n1 ), .A2(
        \sha1_round/add_79/n194 ), .ZN(\sha1_round/add_79/n187 ) );
  NAND2_X2 \sha1_round/add_79/U332  ( .A1(\sha1_round/add_79/n191 ), .A2(
        \sha1_round/add_79/n192 ), .ZN(\sha1_round/add_79/n183 ) );
  INV_X4 \sha1_round/add_79/U331  ( .A(\sha1_round/f [27]), .ZN(
        \sha1_round/add_79/n189 ) );
  NAND2_X2 \sha1_round/add_79/U330  ( .A1(\sha1_round/add_79/n55 ), .A2(
        \sha1_round/add_79/n189 ), .ZN(\sha1_round/add_79/n184 ) );
  XNOR2_X2 \sha1_round/add_79/U329  ( .A(\sha1_round/add_79/n188 ), .B(
        \sha1_round/add_79/n22 ), .ZN(\sha1_round/N279 ) );
  INV_X4 \sha1_round/add_79/U328  ( .A(\sha1_round/add_79/n187 ), .ZN(
        \sha1_round/add_79/n186 ) );
  NAND2_X2 \sha1_round/add_79/U327  ( .A1(\sha1_round/add_79/n186 ), .A2(
        \sha1_round/add_79/n184 ), .ZN(\sha1_round/add_79/n146 ) );
  NAND2_X2 \sha1_round/add_79/U326  ( .A1(\sha1_round/add_79/n183 ), .A2(
        \sha1_round/add_79/n184 ), .ZN(\sha1_round/add_79/n176 ) );
  NAND2_X2 \sha1_round/add_79/U325  ( .A1(\sha1_round/add_79/n176 ), .A2(
        \sha1_round/add_79/n152 ), .ZN(\sha1_round/add_79/n182 ) );
  NAND2_X2 \sha1_round/add_79/U324  ( .A1(\sha1_round/n511 ), .A2(
        \sha1_round/f [28]), .ZN(\sha1_round/add_79/n161 ) );
  INV_X4 \sha1_round/add_79/U323  ( .A(\sha1_round/f [28]), .ZN(
        \sha1_round/add_79/n180 ) );
  NAND2_X2 \sha1_round/add_79/U322  ( .A1(\sha1_round/add_79/n88 ), .A2(
        \sha1_round/add_79/n180 ), .ZN(\sha1_round/add_79/n175 ) );
  NAND2_X2 \sha1_round/add_79/U321  ( .A1(\sha1_round/add_79/n161 ), .A2(
        \sha1_round/add_79/n175 ), .ZN(\sha1_round/add_79/n179 ) );
  INV_X4 \sha1_round/add_79/U320  ( .A(\sha1_round/add_79/n161 ), .ZN(
        \sha1_round/add_79/n177 ) );
  INV_X4 \sha1_round/add_79/U319  ( .A(\sha1_round/add_79/n175 ), .ZN(
        \sha1_round/add_79/n164 ) );
  INV_X4 \sha1_round/add_79/U318  ( .A(\sha1_round/add_79/n176 ), .ZN(
        \sha1_round/add_79/n141 ) );
  NAND2_X2 \sha1_round/add_79/U317  ( .A1(\sha1_round/add_79/n141 ), .A2(
        \sha1_round/add_79/n175 ), .ZN(\sha1_round/add_79/n174 ) );
  NAND2_X2 \sha1_round/add_79/U316  ( .A1(\sha1_round/f [29]), .A2(
        \sha1_round/n825 ), .ZN(\sha1_round/add_79/n162 ) );
  NAND2_X2 \sha1_round/add_79/U315  ( .A1(\sha1_round/add_79/n162 ), .A2(
        \sha1_round/add_79/n165 ), .ZN(\sha1_round/add_79/n171 ) );
  XNOR2_X2 \sha1_round/add_79/U314  ( .A(\sha1_round/add_79/n170 ), .B(
        \sha1_round/add_79/n171 ), .ZN(\sha1_round/N281 ) );
  NAND2_X2 \sha1_round/add_79/U313  ( .A1(\sha1_round/add_79/n169 ), .A2(
        \sha1_round/add_79/n311 ), .ZN(\sha1_round/add_79/n166 ) );
  XNOR2_X2 \sha1_round/add_79/U312  ( .A(\sha1_round/add_79/n166 ), .B(
        \sha1_round/add_79/n134 ), .ZN(\sha1_round/N254 ) );
  INV_X4 \sha1_round/add_79/U311  ( .A(\sha1_round/add_79/n165 ), .ZN(
        \sha1_round/add_79/n160 ) );
  INV_X4 \sha1_round/add_79/U310  ( .A(\sha1_round/add_79/n151 ), .ZN(
        \sha1_round/add_79/n163 ) );
  INV_X4 \sha1_round/add_79/U309  ( .A(\sha1_round/add_79/n148 ), .ZN(
        \sha1_round/add_79/n159 ) );
  NAND2_X2 \sha1_round/add_79/U308  ( .A1(\sha1_round/add_79/n141 ), .A2(
        \sha1_round/add_79/n151 ), .ZN(\sha1_round/add_79/n157 ) );
  NAND2_X2 \sha1_round/add_79/U307  ( .A1(\sha1_round/f [30]), .A2(
        \sha1_round/k_30 ), .ZN(\sha1_round/add_79/n150 ) );
  NAND2_X2 \sha1_round/add_79/U306  ( .A1(\sha1_round/add_79/n150 ), .A2(
        \sha1_round/add_79/n149 ), .ZN(\sha1_round/add_79/n154 ) );
  XNOR2_X2 \sha1_round/add_79/U305  ( .A(\sha1_round/add_79/n153 ), .B(
        \sha1_round/add_79/n154 ), .ZN(\sha1_round/N282 ) );
  NAND2_X2 \sha1_round/add_79/U304  ( .A1(\sha1_round/add_79/n151 ), .A2(
        \sha1_round/add_79/n149 ), .ZN(\sha1_round/add_79/n143 ) );
  INV_X4 \sha1_round/add_79/U303  ( .A(\sha1_round/add_79/n149 ), .ZN(
        \sha1_round/add_79/n147 ) );
  INV_X4 \sha1_round/add_79/U302  ( .A(\sha1_round/add_79/n146 ), .ZN(
        \sha1_round/add_79/n144 ) );
  INV_X4 \sha1_round/add_79/U301  ( .A(\sha1_round/add_79/n143 ), .ZN(
        \sha1_round/add_79/n142 ) );
  NAND2_X2 \sha1_round/add_79/U300  ( .A1(\sha1_round/add_79/n141 ), .A2(
        \sha1_round/add_79/n142 ), .ZN(\sha1_round/add_79/n140 ) );
  NAND4_X2 \sha1_round/add_79/U299  ( .A1(\sha1_round/add_79/n137 ), .A2(
        \sha1_round/add_79/n138 ), .A3(\sha1_round/add_79/n139 ), .A4(
        \sha1_round/add_79/n140 ), .ZN(\sha1_round/add_79/n135 ) );
  XNOR2_X2 \sha1_round/add_79/U298  ( .A(\sha1_round/f [31]), .B(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n136 ) );
  XNOR2_X2 \sha1_round/add_79/U297  ( .A(\sha1_round/add_79/n135 ), .B(
        \sha1_round/add_79/n136 ), .ZN(\sha1_round/N283 ) );
  INV_X4 \sha1_round/add_79/U296  ( .A(\sha1_round/add_79/n134 ), .ZN(
        \sha1_round/add_79/n133 ) );
  INV_X4 \sha1_round/add_79/U295  ( .A(\sha1_round/add_79/n311 ), .ZN(
        \sha1_round/add_79/n131 ) );
  XNOR2_X2 \sha1_round/add_79/U294  ( .A(\sha1_round/add_79/n127 ), .B(
        \sha1_round/add_79/n128 ), .ZN(\sha1_round/N255 ) );
  XNOR2_X2 \sha1_round/add_79/U293  ( .A(\sha1_round/add_79/n126 ), .B(
        \sha1_round/add_79/n63 ), .ZN(\sha1_round/N256 ) );
  NAND2_X2 \sha1_round/add_79/U292  ( .A1(\sha1_round/add_79/n125 ), .A2(
        \sha1_round/add_79/n119 ), .ZN(\sha1_round/add_79/n122 ) );
  INV_X4 \sha1_round/add_79/U291  ( .A(\sha1_round/add_79/n124 ), .ZN(
        \sha1_round/add_79/n123 ) );
  XNOR2_X2 \sha1_round/add_79/U290  ( .A(\sha1_round/add_79/n122 ), .B(
        \sha1_round/add_79/n123 ), .ZN(\sha1_round/N257 ) );
  INV_X4 \sha1_round/add_79/U289  ( .A(\sha1_round/add_79/n120 ), .ZN(
        \sha1_round/add_79/n117 ) );
  XNOR2_X2 \sha1_round/add_79/U288  ( .A(\sha1_round/add_79/n115 ), .B(
        \sha1_round/add_79/n116 ), .ZN(\sha1_round/N258 ) );
  NAND2_X2 \sha1_round/add_79/U287  ( .A1(\sha1_round/add_79/n104 ), .A2(
        \sha1_round/add_79/n105 ), .ZN(\sha1_round/add_79/n102 ) );
  INV_X4 \sha1_round/add_79/U286  ( .A(\sha1_round/add_79/n100 ), .ZN(
        \sha1_round/add_79/n103 ) );
  INV_X4 \sha1_round/add_79/U285  ( .A(\sha1_round/add_79/n96 ), .ZN(
        \sha1_round/add_79/n95 ) );
  XNOR2_X2 \sha1_round/add_79/U284  ( .A(\sha1_round/add_79/n93 ), .B(
        \sha1_round/add_79/n94 ), .ZN(\sha1_round/N261 ) );
  NAND2_X1 \sha1_round/add_79/U283  ( .A1(\sha1_round/n2 ), .A2(
        \sha1_round/f [4]), .ZN(\sha1_round/add_79/n119 ) );
  NAND2_X1 \sha1_round/add_79/U282  ( .A1(\sha1_round/f [17]), .A2(
        \sha1_round/n2 ), .ZN(\sha1_round/add_79/n275 ) );
  NAND3_X2 \sha1_round/add_79/U281  ( .A1(\sha1_round/add_79/n109 ), .A2(
        \sha1_round/add_79/n31 ), .A3(\sha1_round/add_79/n110 ), .ZN(
        \sha1_round/add_79/n332 ) );
  NAND3_X1 \sha1_round/add_79/U280  ( .A1(\sha1_round/add_79/n31 ), .A2(
        \sha1_round/add_79/n107 ), .A3(\sha1_round/add_79/n106 ), .ZN(
        \sha1_round/add_79/n338 ) );
  NOR2_X1 \sha1_round/add_79/U279  ( .A1(\sha1_round/add_79/n26 ), .A2(
        \sha1_round/add_79/n129 ), .ZN(\sha1_round/add_79/n128 ) );
  NAND3_X2 \sha1_round/add_79/U278  ( .A1(\sha1_round/add_79/n107 ), .A2(
        \sha1_round/add_79/n121 ), .A3(\sha1_round/add_79/n8 ), .ZN(
        \sha1_round/add_79/n120 ) );
  NAND3_X1 \sha1_round/add_79/U277  ( .A1(\sha1_round/add_79/n151 ), .A2(
        \sha1_round/add_79/n144 ), .A3(\sha1_round/add_79/n145 ), .ZN(
        \sha1_round/add_79/n156 ) );
  NAND3_X1 \sha1_round/add_79/U276  ( .A1(\sha1_round/add_79/n142 ), .A2(
        \sha1_round/add_79/n144 ), .A3(\sha1_round/add_79/n145 ), .ZN(
        \sha1_round/add_79/n139 ) );
  NAND2_X4 \sha1_round/add_79/U275  ( .A1(\sha1_round/add_79/n354 ), .A2(
        \sha1_round/add_79/n355 ), .ZN(\sha1_round/add_79/n340 ) );
  INV_X2 \sha1_round/add_79/U274  ( .A(\sha1_round/add_79/n167 ), .ZN(
        \sha1_round/add_79/n269 ) );
  NAND2_X2 \sha1_round/add_79/U273  ( .A1(\sha1_round/add_79/n1 ), .A2(
        \sha1_round/add_79/n145 ), .ZN(\sha1_round/add_79/n204 ) );
  NAND2_X2 \sha1_round/add_79/U272  ( .A1(\sha1_round/add_79/n205 ), .A2(
        \sha1_round/add_79/n145 ), .ZN(\sha1_round/add_79/n211 ) );
  INV_X2 \sha1_round/add_79/U271  ( .A(\sha1_round/add_79/n101 ), .ZN(
        \sha1_round/add_79/n97 ) );
  NOR2_X2 \sha1_round/add_79/U270  ( .A1(\sha1_round/f [7]), .A2(
        \sha1_round/k_27 ), .ZN(\sha1_round/add_79/n111 ) );
  NAND2_X1 \sha1_round/add_79/U269  ( .A1(\sha1_round/add_79/n2 ), .A2(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n375 ) );
  NAND3_X2 \sha1_round/add_79/U268  ( .A1(\sha1_round/add_79/n234 ), .A2(
        \sha1_round/add_79/n235 ), .A3(\sha1_round/add_79/n236 ), .ZN(
        \sha1_round/add_79/n226 ) );
  NOR2_X1 \sha1_round/add_79/U267  ( .A1(\sha1_round/f [0]), .A2(
        \sha1_round/k_23 ), .ZN(\sha1_round/add_79/n271 ) );
  NAND2_X1 \sha1_round/add_79/U266  ( .A1(\sha1_round/add_79/n359 ), .A2(
        \sha1_round/add_79/n344 ), .ZN(\sha1_round/add_79/n361 ) );
  NAND3_X1 \sha1_round/add_79/U265  ( .A1(\sha1_round/add_79/n144 ), .A2(
        \sha1_round/add_79/n175 ), .A3(\sha1_round/add_79/n145 ), .ZN(
        \sha1_round/add_79/n173 ) );
  INV_X4 \sha1_round/add_79/U264  ( .A(\sha1_round/f [18]), .ZN(
        \sha1_round/add_79/n262 ) );
  NAND2_X2 \sha1_round/add_79/U263  ( .A1(\sha1_round/add_79/n266 ), .A2(
        \sha1_round/add_79/n267 ), .ZN(\sha1_round/add_79/n263 ) );
  AND2_X2 \sha1_round/add_79/U262  ( .A1(\sha1_round/k_27 ), .A2(
        \sha1_round/f [7]), .ZN(\sha1_round/add_79/n83 ) );
  NOR3_X2 \sha1_round/add_79/U261  ( .A1(\sha1_round/add_79/n310 ), .A2(
        \sha1_round/add_79/n269 ), .A3(\sha1_round/add_79/n129 ), .ZN(
        \sha1_round/add_79/n309 ) );
  NAND3_X1 \sha1_round/add_79/U260  ( .A1(\sha1_round/f [18]), .A2(
        \sha1_round/add_79/n27 ), .A3(\sha1_round/add_79/n250 ), .ZN(
        \sha1_round/add_79/n267 ) );
  NAND3_X2 \sha1_round/add_79/U259  ( .A1(\sha1_round/add_79/n294 ), .A2(
        \sha1_round/add_79/n295 ), .A3(\sha1_round/add_79/n24 ), .ZN(
        \sha1_round/add_79/n288 ) );
  AND2_X2 \sha1_round/add_79/U258  ( .A1(\sha1_round/add_79/n257 ), .A2(
        \sha1_round/add_79/n258 ), .ZN(\sha1_round/add_79/n82 ) );
  AND2_X2 \sha1_round/add_79/U257  ( .A1(\sha1_round/add_79/n2 ), .A2(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n81 ) );
  NOR2_X2 \sha1_round/add_79/U256  ( .A1(\sha1_round/f [8]), .A2(
        \sha1_round/k_30 ), .ZN(\sha1_round/add_79/n348 ) );
  AND2_X2 \sha1_round/add_79/U255  ( .A1(\sha1_round/n825 ), .A2(
        \sha1_round/add_79/n33 ), .ZN(\sha1_round/add_79/n80 ) );
  NOR2_X1 \sha1_round/add_79/U254  ( .A1(\sha1_round/n2 ), .A2(
        \sha1_round/f [17]), .ZN(\sha1_round/add_79/n79 ) );
  NAND3_X1 \sha1_round/add_79/U253  ( .A1(\sha1_round/f [23]), .A2(
        \sha1_round/add_79/n25 ), .A3(\sha1_round/k_23 ), .ZN(
        \sha1_round/add_79/n197 ) );
  NOR2_X1 \sha1_round/add_79/U252  ( .A1(\sha1_round/f [23]), .A2(
        \sha1_round/k_23 ), .ZN(\sha1_round/add_79/n213 ) );
  NOR2_X2 \sha1_round/add_79/U251  ( .A1(\sha1_round/add_79/n381 ), .A2(
        \sha1_round/add_79/n271 ), .ZN(\sha1_round/N252 ) );
  INV_X1 \sha1_round/add_79/U250  ( .A(\sha1_round/n511 ), .ZN(
        \sha1_round/add_79/n88 ) );
  INV_X1 \sha1_round/add_79/U249  ( .A(\sha1_round/n3370 ), .ZN(
        \sha1_round/add_79/n91 ) );
  OR2_X2 \sha1_round/add_79/U248  ( .A1(\sha1_round/add_79/n152 ), .A2(
        \sha1_round/add_79/n143 ), .ZN(\sha1_round/add_79/n137 ) );
  INV_X4 \sha1_round/add_79/U247  ( .A(\sha1_round/add_79/n86 ), .ZN(
        \sha1_round/add_79/n87 ) );
  OR2_X4 \sha1_round/add_79/U246  ( .A1(\sha1_round/add_79/n348 ), .A2(
        \sha1_round/add_79/n103 ), .ZN(\sha1_round/add_79/n77 ) );
  XNOR2_X2 \sha1_round/add_79/U245  ( .A(\sha1_round/add_79/n102 ), .B(
        \sha1_round/add_79/n77 ), .ZN(\sha1_round/N260 ) );
  NOR2_X2 \sha1_round/add_79/U244  ( .A1(\sha1_round/add_79/n212 ), .A2(
        \sha1_round/add_79/n214 ), .ZN(\sha1_round/add_79/n218 ) );
  OR2_X4 \sha1_round/add_79/U243  ( .A1(\sha1_round/add_79/n147 ), .A2(
        \sha1_round/add_79/n148 ), .ZN(\sha1_round/add_79/n75 ) );
  AND2_X2 \sha1_round/add_79/U242  ( .A1(\sha1_round/add_79/n150 ), .A2(
        \sha1_round/add_79/n75 ), .ZN(\sha1_round/add_79/n138 ) );
  NAND3_X2 \sha1_round/add_79/U241  ( .A1(\sha1_round/add_79/n230 ), .A2(
        \sha1_round/add_79/n231 ), .A3(\sha1_round/add_79/n232 ), .ZN(
        \sha1_round/add_79/n225 ) );
  NOR2_X1 \sha1_round/add_79/U240  ( .A1(\sha1_round/add_79/n74 ), .A2(
        \sha1_round/add_79/n227 ), .ZN(\sha1_round/add_79/n223 ) );
  NAND3_X1 \sha1_round/add_79/U239  ( .A1(\sha1_round/add_79/n242 ), .A2(
        \sha1_round/add_79/n240 ), .A3(\sha1_round/add_79/n250 ), .ZN(
        \sha1_round/add_79/n249 ) );
  OR2_X4 \sha1_round/add_79/U238  ( .A1(\sha1_round/add_79/n160 ), .A2(
        \sha1_round/add_79/n161 ), .ZN(\sha1_round/add_79/n73 ) );
  AND2_X2 \sha1_round/add_79/U237  ( .A1(\sha1_round/add_79/n162 ), .A2(
        \sha1_round/add_79/n73 ), .ZN(\sha1_round/add_79/n148 ) );
  XNOR2_X2 \sha1_round/add_79/U236  ( .A(\sha1_round/add_79/n263 ), .B(
        \sha1_round/add_79/n264 ), .ZN(\sha1_round/N272 ) );
  NOR2_X2 \sha1_round/add_79/U235  ( .A1(\sha1_round/add_79/n163 ), .A2(
        \sha1_round/add_79/n152 ), .ZN(\sha1_round/add_79/n158 ) );
  NOR2_X2 \sha1_round/add_79/U234  ( .A1(\sha1_round/add_79/n164 ), .A2(
        \sha1_round/add_79/n152 ), .ZN(\sha1_round/add_79/n178 ) );
  NOR2_X1 \sha1_round/add_79/U233  ( .A1(\sha1_round/add_79/n349 ), .A2(
        \sha1_round/add_79/n346 ), .ZN(\sha1_round/add_79/n357 ) );
  NOR2_X2 \sha1_round/add_79/U232  ( .A1(\sha1_round/add_79/n212 ), .A2(
        \sha1_round/add_79/n213 ), .ZN(\sha1_round/add_79/n205 ) );
  OR2_X2 \sha1_round/add_79/U231  ( .A1(\sha1_round/add_79/n253 ), .A2(
        \sha1_round/add_79/n82 ), .ZN(\sha1_round/add_79/n69 ) );
  NAND3_X2 \sha1_round/add_79/U230  ( .A1(\sha1_round/add_79/n196 ), .A2(
        \sha1_round/add_79/n197 ), .A3(\sha1_round/add_79/n198 ), .ZN(
        \sha1_round/add_79/n195 ) );
  NAND3_X2 \sha1_round/add_79/U229  ( .A1(\sha1_round/add_79/n193 ), .A2(
        \sha1_round/add_79/n194 ), .A3(\sha1_round/add_79/n195 ), .ZN(
        \sha1_round/add_79/n191 ) );
  NOR2_X2 \sha1_round/add_79/U228  ( .A1(\sha1_round/add_79/n214 ), .A2(
        \sha1_round/add_79/n215 ), .ZN(\sha1_round/add_79/n210 ) );
  NOR2_X2 \sha1_round/add_79/U227  ( .A1(\sha1_round/add_79/n158 ), .A2(
        \sha1_round/add_79/n159 ), .ZN(\sha1_round/add_79/n155 ) );
  NAND3_X2 \sha1_round/add_79/U226  ( .A1(\sha1_round/add_79/n155 ), .A2(
        \sha1_round/add_79/n156 ), .A3(\sha1_round/add_79/n157 ), .ZN(
        \sha1_round/add_79/n153 ) );
  NOR2_X2 \sha1_round/add_79/U225  ( .A1(\sha1_round/add_79/n177 ), .A2(
        \sha1_round/add_79/n178 ), .ZN(\sha1_round/add_79/n172 ) );
  NAND3_X2 \sha1_round/add_79/U224  ( .A1(\sha1_round/add_79/n172 ), .A2(
        \sha1_round/add_79/n173 ), .A3(\sha1_round/add_79/n174 ), .ZN(
        \sha1_round/add_79/n170 ) );
  NOR2_X2 \sha1_round/add_79/U223  ( .A1(\sha1_round/add_79/n308 ), .A2(
        \sha1_round/add_79/n129 ), .ZN(\sha1_round/add_79/n367 ) );
  INV_X1 \sha1_round/add_79/U222  ( .A(\sha1_round/n512 ), .ZN(
        \sha1_round/add_79/n90 ) );
  XNOR2_X2 \sha1_round/add_79/U221  ( .A(\sha1_round/add_79/n245 ), .B(
        \sha1_round/add_79/n246 ), .ZN(\sha1_round/N274 ) );
  NAND3_X2 \sha1_round/add_79/U220  ( .A1(\sha1_round/add_79/n235 ), .A2(
        \sha1_round/add_79/n297 ), .A3(\sha1_round/add_79/n236 ), .ZN(
        \sha1_round/add_79/n287 ) );
  NOR2_X1 \sha1_round/add_79/U219  ( .A1(\sha1_round/add_79/n185 ), .A2(
        \sha1_round/add_79/n146 ), .ZN(\sha1_round/add_79/n181 ) );
  NOR2_X2 \sha1_round/add_79/U218  ( .A1(\sha1_round/add_79/n160 ), .A2(
        \sha1_round/add_79/n164 ), .ZN(\sha1_round/add_79/n151 ) );
  INV_X4 \sha1_round/add_79/U217  ( .A(\sha1_round/add_79/n90 ), .ZN(
        \sha1_round/add_79/n89 ) );
  NAND2_X4 \sha1_round/add_79/U216  ( .A1(\sha1_round/add_79/n362 ), .A2(
        \sha1_round/add_79/n90 ), .ZN(\sha1_round/add_79/n359 ) );
  INV_X1 \sha1_round/add_79/U215  ( .A(\sha1_round/add_79/n270 ), .ZN(
        \sha1_round/add_79/n381 ) );
  OR2_X4 \sha1_round/add_79/U214  ( .A1(\sha1_round/n825 ), .A2(
        \sha1_round/f [29]), .ZN(\sha1_round/add_79/n165 ) );
  OR2_X4 \sha1_round/add_79/U213  ( .A1(\sha1_round/k_30 ), .A2(
        \sha1_round/f [30]), .ZN(\sha1_round/add_79/n149 ) );
  NOR2_X2 \sha1_round/add_79/U212  ( .A1(\sha1_round/add_79/n309 ), .A2(
        \sha1_round/add_79/n108 ), .ZN(\sha1_round/add_79/n304 ) );
  OR2_X4 \sha1_round/add_79/U211  ( .A1(\sha1_round/n824 ), .A2(
        \sha1_round/f [21]), .ZN(\sha1_round/add_79/n240 ) );
  NOR2_X2 \sha1_round/add_79/U210  ( .A1(\sha1_round/add_79/n181 ), .A2(
        \sha1_round/add_79/n182 ), .ZN(\sha1_round/add_79/n64 ) );
  XOR2_X2 \sha1_round/add_79/U209  ( .A(\sha1_round/add_79/n64 ), .B(
        \sha1_round/add_79/n179 ), .Z(\sha1_round/N280 ) );
  AND2_X4 \sha1_round/add_79/U208  ( .A1(\sha1_round/add_79/n244 ), .A2(
        \sha1_round/add_79/n241 ), .ZN(\sha1_round/add_79/n74 ) );
  INV_X1 \sha1_round/add_79/U207  ( .A(\sha1_round/add_79/n308 ), .ZN(
        \sha1_round/add_79/n307 ) );
  NAND3_X1 \sha1_round/add_79/U206  ( .A1(\sha1_round/add_79/n198 ), .A2(
        \sha1_round/add_79/n196 ), .A3(\sha1_round/add_79/n197 ), .ZN(
        \sha1_round/add_79/n206 ) );
  NOR2_X2 \sha1_round/add_79/U205  ( .A1(\sha1_round/add_79/n12 ), .A2(
        \sha1_round/add_79/n238 ), .ZN(\sha1_round/add_79/n277 ) );
  NAND4_X1 \sha1_round/add_79/U204  ( .A1(\sha1_round/add_79/n223 ), .A2(
        \sha1_round/add_79/n224 ), .A3(\sha1_round/add_79/n225 ), .A4(
        \sha1_round/add_79/n226 ), .ZN(\sha1_round/add_79/n221 ) );
  NOR2_X1 \sha1_round/add_79/U203  ( .A1(\sha1_round/add_79/n79 ), .A2(
        \sha1_round/add_79/n278 ), .ZN(\sha1_round/add_79/n231 ) );
  OR2_X4 \sha1_round/add_79/U202  ( .A1(\sha1_round/add_79/n168 ), .A2(
        \sha1_round/add_79/n270 ), .ZN(\sha1_round/add_79/n68 ) );
  NOR2_X1 \sha1_round/add_79/U201  ( .A1(\sha1_round/add_79/n380 ), .A2(
        \sha1_round/add_79/n119 ), .ZN(\sha1_round/add_79/n118 ) );
  NOR2_X1 \sha1_round/add_79/U200  ( .A1(\sha1_round/add_79/n347 ), .A2(
        \sha1_round/add_79/n345 ), .ZN(\sha1_round/add_79/n353 ) );
  NAND3_X2 \sha1_round/add_79/U199  ( .A1(\sha1_round/add_79/n277 ), .A2(
        \sha1_round/add_79/n235 ), .A3(\sha1_round/add_79/n236 ), .ZN(
        \sha1_round/add_79/n276 ) );
  INV_X1 \sha1_round/add_79/U198  ( .A(\sha1_round/n517 ), .ZN(
        \sha1_round/add_79/n92 ) );
  NOR2_X1 \sha1_round/add_79/U197  ( .A1(\sha1_round/f [24]), .A2(
        \sha1_round/add_79/n89 ), .ZN(\sha1_round/add_79/n212 ) );
  NAND3_X2 \sha1_round/add_79/U196  ( .A1(\sha1_round/add_79/n313 ), .A2(
        \sha1_round/add_79/n314 ), .A3(\sha1_round/add_79/n315 ), .ZN(
        \sha1_round/add_79/n238 ) );
  INV_X4 \sha1_round/add_79/U195  ( .A(\sha1_round/add_79/n60 ), .ZN(
        \sha1_round/add_79/n61 ) );
  NAND2_X2 \sha1_round/add_79/U194  ( .A1(\sha1_round/add_79/n13 ), .A2(
        \sha1_round/add_79/n319 ), .ZN(\sha1_round/add_79/n235 ) );
  INV_X1 \sha1_round/add_79/U193  ( .A(\sha1_round/add_79/n317 ), .ZN(
        \sha1_round/add_79/n327 ) );
  NOR2_X1 \sha1_round/add_79/U192  ( .A1(\sha1_round/add_79/n185 ), .A2(
        \sha1_round/add_79/n187 ), .ZN(\sha1_round/add_79/n190 ) );
  NAND2_X1 \sha1_round/add_79/U191  ( .A1(\sha1_round/add_79/n233 ), .A2(
        \sha1_round/add_79/n280 ), .ZN(\sha1_round/add_79/n291 ) );
  INV_X2 \sha1_round/add_79/U190  ( .A(\sha1_round/add_79/n291 ), .ZN(
        \sha1_round/add_79/n57 ) );
  INV_X4 \sha1_round/add_79/U189  ( .A(\sha1_round/add_79/n290 ), .ZN(
        \sha1_round/add_79/n56 ) );
  NAND2_X4 \sha1_round/add_79/U188  ( .A1(\sha1_round/add_79/n58 ), .A2(
        \sha1_round/add_79/n59 ), .ZN(\sha1_round/N268 ) );
  NAND2_X4 \sha1_round/add_79/U187  ( .A1(\sha1_round/add_79/n56 ), .A2(
        \sha1_round/add_79/n57 ), .ZN(\sha1_round/add_79/n59 ) );
  NAND2_X2 \sha1_round/add_79/U186  ( .A1(\sha1_round/add_79/n291 ), .A2(
        \sha1_round/add_79/n290 ), .ZN(\sha1_round/add_79/n58 ) );
  NAND2_X4 \sha1_round/add_79/U185  ( .A1(\sha1_round/add_79/n322 ), .A2(
        \sha1_round/add_79/n294 ), .ZN(\sha1_round/add_79/n320 ) );
  NAND3_X2 \sha1_round/add_79/U184  ( .A1(\sha1_round/add_79/n104 ), .A2(
        \sha1_round/add_79/n298 ), .A3(\sha1_round/add_79/n299 ), .ZN(
        \sha1_round/add_79/n236 ) );
  NAND2_X1 \sha1_round/add_79/U183  ( .A1(\sha1_round/n517 ), .A2(
        \sha1_round/f [3]), .ZN(\sha1_round/add_79/n306 ) );
  NAND2_X1 \sha1_round/add_79/U182  ( .A1(\sha1_round/add_79/n87 ), .A2(
        \sha1_round/f [2]), .ZN(\sha1_round/add_79/n311 ) );
  NOR2_X4 \sha1_round/add_79/U181  ( .A1(\sha1_round/f [5]), .A2(
        \sha1_round/n825 ), .ZN(\sha1_round/add_79/n380 ) );
  NAND2_X2 \sha1_round/add_79/U180  ( .A1(\sha1_round/add_79/n4 ), .A2(
        \sha1_round/add_79/n101 ), .ZN(\sha1_round/add_79/n364 ) );
  XNOR2_X2 \sha1_round/add_79/U179  ( .A(\sha1_round/add_79/n325 ), .B(
        \sha1_round/add_79/n326 ), .ZN(\sha1_round/N266 ) );
  NOR2_X4 \sha1_round/add_79/U178  ( .A1(\sha1_round/f [9]), .A2(
        \sha1_round/n825 ), .ZN(\sha1_round/add_79/n349 ) );
  NAND2_X1 \sha1_round/add_79/U177  ( .A1(\sha1_round/f [9]), .A2(
        \sha1_round/n825 ), .ZN(\sha1_round/add_79/n96 ) );
  NAND3_X2 \sha1_round/add_79/U176  ( .A1(\sha1_round/add_79/n33 ), .A2(
        \sha1_round/add_79/n85 ), .A3(\sha1_round/n825 ), .ZN(
        \sha1_round/add_79/n374 ) );
  NOR2_X2 \sha1_round/add_79/U175  ( .A1(\sha1_round/add_79/n115 ), .A2(
        \sha1_round/add_79/n379 ), .ZN(\sha1_round/add_79/n114 ) );
  OR2_X4 \sha1_round/add_79/U174  ( .A1(\sha1_round/add_79/n84 ), .A2(
        \sha1_round/add_79/n312 ), .ZN(\sha1_round/add_79/n78 ) );
  NAND2_X4 \sha1_round/add_79/U173  ( .A1(\sha1_round/add_79/n53 ), .A2(
        \sha1_round/add_79/n54 ), .ZN(\sha1_round/N267 ) );
  NAND2_X4 \sha1_round/add_79/U172  ( .A1(\sha1_round/add_79/n51 ), .A2(
        \sha1_round/add_79/n52 ), .ZN(\sha1_round/add_79/n54 ) );
  INV_X4 \sha1_round/add_79/U171  ( .A(\sha1_round/add_79/n49 ), .ZN(
        \sha1_round/add_79/n50 ) );
  NAND2_X4 \sha1_round/add_79/U170  ( .A1(\sha1_round/add_79/n50 ), .A2(
        \sha1_round/add_79/n226 ), .ZN(\sha1_round/add_79/n145 ) );
  NAND2_X4 \sha1_round/add_79/U169  ( .A1(\sha1_round/add_79/n23 ), .A2(
        \sha1_round/add_79/n35 ), .ZN(\sha1_round/add_79/n303 ) );
  NAND2_X4 \sha1_round/add_79/U168  ( .A1(\sha1_round/add_79/n61 ), .A2(
        \sha1_round/add_79/n63 ), .ZN(\sha1_round/add_79/n101 ) );
  NAND2_X4 \sha1_round/add_79/U167  ( .A1(\sha1_round/add_79/n48 ), .A2(
        \sha1_round/add_79/n47 ), .ZN(\sha1_round/N259 ) );
  NAND2_X4 \sha1_round/add_79/U166  ( .A1(\sha1_round/add_79/n45 ), .A2(
        \sha1_round/add_79/n46 ), .ZN(\sha1_round/add_79/n48 ) );
  INV_X2 \sha1_round/add_79/U165  ( .A(\sha1_round/add_79/n361 ), .ZN(
        \sha1_round/add_79/n42 ) );
  NAND2_X4 \sha1_round/add_79/U164  ( .A1(\sha1_round/add_79/n43 ), .A2(
        \sha1_round/add_79/n44 ), .ZN(\sha1_round/N262 ) );
  NAND2_X4 \sha1_round/add_79/U163  ( .A1(\sha1_round/add_79/n41 ), .A2(
        \sha1_round/add_79/n42 ), .ZN(\sha1_round/add_79/n44 ) );
  NOR2_X2 \sha1_round/add_79/U162  ( .A1(\sha1_round/add_79/n239 ), .A2(
        \sha1_round/add_79/n79 ), .ZN(\sha1_round/add_79/n283 ) );
  INV_X4 \sha1_round/add_79/U161  ( .A(\sha1_round/add_79/n283 ), .ZN(
        \sha1_round/add_79/n38 ) );
  NAND2_X4 \sha1_round/add_79/U160  ( .A1(\sha1_round/add_79/n39 ), .A2(
        \sha1_round/add_79/n40 ), .ZN(\sha1_round/add_79/n281 ) );
  NAND2_X4 \sha1_round/add_79/U159  ( .A1(\sha1_round/add_79/n37 ), .A2(
        \sha1_round/add_79/n38 ), .ZN(\sha1_round/add_79/n40 ) );
  NAND2_X2 \sha1_round/add_79/U158  ( .A1(\sha1_round/add_79/n282 ), .A2(
        \sha1_round/add_79/n283 ), .ZN(\sha1_round/add_79/n39 ) );
  INV_X2 \sha1_round/add_79/U157  ( .A(\sha1_round/add_79/n348 ), .ZN(
        \sha1_round/add_79/n366 ) );
  NAND2_X2 \sha1_round/add_79/U156  ( .A1(\sha1_round/f [1]), .A2(
        \sha1_round/n824 ), .ZN(\sha1_round/add_79/n370 ) );
  NAND2_X2 \sha1_round/add_79/U155  ( .A1(\sha1_round/n824 ), .A2(
        \sha1_round/f [1]), .ZN(\sha1_round/add_79/n167 ) );
  NAND2_X1 \sha1_round/add_79/U154  ( .A1(\sha1_round/f [13]), .A2(
        \sha1_round/k[13] ), .ZN(\sha1_round/add_79/n323 ) );
  NAND2_X4 \sha1_round/add_79/U153  ( .A1(\sha1_round/add_79/n109 ), .A2(
        \sha1_round/add_79/n21 ), .ZN(\sha1_round/add_79/n99 ) );
  NAND3_X2 \sha1_round/add_79/U152  ( .A1(\sha1_round/add_79/n36 ), .A2(
        \sha1_round/add_79/n344 ), .A3(\sha1_round/add_79/n343 ), .ZN(
        \sha1_round/add_79/n35 ) );
  NOR3_X2 \sha1_round/add_79/U151  ( .A1(\sha1_round/add_79/n78 ), .A2(
        \sha1_round/add_79/n132 ), .A3(\sha1_round/add_79/n168 ), .ZN(
        \sha1_round/add_79/n369 ) );
  NAND3_X2 \sha1_round/add_79/U150  ( .A1(\sha1_round/add_79/n101 ), .A2(
        \sha1_round/add_79/n99 ), .A3(\sha1_round/add_79/n14 ), .ZN(
        \sha1_round/add_79/n358 ) );
  INV_X1 \sha1_round/add_79/U149  ( .A(\sha1_round/add_79/n82 ), .ZN(
        \sha1_round/add_79/n256 ) );
  INV_X2 \sha1_round/add_79/U148  ( .A(\sha1_round/add_79/n132 ), .ZN(
        \sha1_round/add_79/n169 ) );
  NAND2_X2 \sha1_round/add_79/U147  ( .A1(\sha1_round/add_79/n112 ), .A2(
        \sha1_round/add_79/n113 ), .ZN(\sha1_round/add_79/n47 ) );
  INV_X4 \sha1_round/add_79/U146  ( .A(\sha1_round/add_79/n113 ), .ZN(
        \sha1_round/add_79/n46 ) );
  NOR2_X2 \sha1_round/add_79/U145  ( .A1(\sha1_round/add_79/n111 ), .A2(
        \sha1_round/add_79/n83 ), .ZN(\sha1_round/add_79/n113 ) );
  INV_X2 \sha1_round/add_79/U144  ( .A(\sha1_round/add_79/n111 ), .ZN(
        \sha1_round/add_79/n110 ) );
  OR2_X4 \sha1_round/add_79/U143  ( .A1(\sha1_round/k[15] ), .A2(
        \sha1_round/f [15]), .ZN(\sha1_round/add_79/n289 ) );
  NAND2_X1 \sha1_round/add_79/U142  ( .A1(\sha1_round/add_79/n295 ), .A2(
        \sha1_round/add_79/n289 ), .ZN(\sha1_round/add_79/n321 ) );
  NOR2_X1 \sha1_round/add_79/U141  ( .A1(\sha1_round/add_79/n269 ), .A2(
        \sha1_round/add_79/n168 ), .ZN(\sha1_round/add_79/n268 ) );
  INV_X2 \sha1_round/add_79/U140  ( .A(\sha1_round/n3170 ), .ZN(
        \sha1_round/add_79/n86 ) );
  NAND2_X1 \sha1_round/add_79/U139  ( .A1(\sha1_round/f [21]), .A2(
        \sha1_round/n824 ), .ZN(\sha1_round/add_79/n252 ) );
  NOR2_X4 \sha1_round/add_79/U138  ( .A1(\sha1_round/add_79/n300 ), .A2(
        \sha1_round/add_79/n301 ), .ZN(\sha1_round/add_79/n299 ) );
  INV_X4 \sha1_round/add_79/U137  ( .A(\sha1_round/add_79/n324 ), .ZN(
        \sha1_round/add_79/n328 ) );
  INV_X4 \sha1_round/add_79/U136  ( .A(\sha1_round/add_79/n282 ), .ZN(
        \sha1_round/add_79/n37 ) );
  NAND2_X4 \sha1_round/add_79/U135  ( .A1(\sha1_round/f [11]), .A2(
        \sha1_round/k[13] ), .ZN(\sha1_round/add_79/n343 ) );
  NOR2_X2 \sha1_round/add_79/U134  ( .A1(\sha1_round/add_79/n260 ), .A2(
        \sha1_round/add_79/n251 ), .ZN(\sha1_round/add_79/n255 ) );
  INV_X4 \sha1_round/add_79/U133  ( .A(\sha1_round/add_79/n250 ), .ZN(
        \sha1_round/add_79/n260 ) );
  NAND2_X4 \sha1_round/add_79/U132  ( .A1(\sha1_round/f [10]), .A2(
        \sha1_round/add_79/n89 ), .ZN(\sha1_round/add_79/n344 ) );
  NOR2_X4 \sha1_round/add_79/U131  ( .A1(\sha1_round/add_79/n117 ), .A2(
        \sha1_round/add_79/n18 ), .ZN(\sha1_round/add_79/n115 ) );
  NAND2_X1 \sha1_round/add_79/U130  ( .A1(\sha1_round/add_79/n311 ), .A2(
        \sha1_round/add_79/n312 ), .ZN(\sha1_round/add_79/n310 ) );
  OR2_X4 \sha1_round/add_79/U129  ( .A1(\sha1_round/add_79/n261 ), .A2(
        \sha1_round/add_79/n272 ), .ZN(\sha1_round/add_79/n34 ) );
  XNOR2_X2 \sha1_round/add_79/U128  ( .A(\sha1_round/add_79/n273 ), .B(
        \sha1_round/add_79/n34 ), .ZN(\sha1_round/N271 ) );
  NOR2_X1 \sha1_round/add_79/U127  ( .A1(\sha1_round/add_79/n80 ), .A2(
        \sha1_round/add_79/n380 ), .ZN(\sha1_round/add_79/n124 ) );
  INV_X2 \sha1_round/add_79/U126  ( .A(\sha1_round/add_79/n359 ), .ZN(
        \sha1_round/add_79/n346 ) );
  NAND2_X2 \sha1_round/add_79/U125  ( .A1(\sha1_round/add_79/n365 ), .A2(
        \sha1_round/add_79/n359 ), .ZN(\sha1_round/add_79/n36 ) );
  INV_X1 \sha1_round/add_79/U124  ( .A(\sha1_round/add_79/n244 ), .ZN(
        \sha1_round/add_79/n248 ) );
  NAND2_X4 \sha1_round/add_79/U123  ( .A1(\sha1_round/add_79/n68 ), .A2(
        \sha1_round/add_79/n167 ), .ZN(\sha1_round/add_79/n134 ) );
  NAND2_X2 \sha1_round/add_79/U122  ( .A1(\sha1_round/n825 ), .A2(
        \sha1_round/f [9]), .ZN(\sha1_round/add_79/n342 ) );
  NAND2_X2 \sha1_round/add_79/U121  ( .A1(\sha1_round/add_79/n336 ), .A2(
        \sha1_round/add_79/n313 ), .ZN(\sha1_round/add_79/n335 ) );
  INV_X4 \sha1_round/add_79/U120  ( .A(\sha1_round/add_79/n32 ), .ZN(
        \sha1_round/add_79/n33 ) );
  INV_X1 \sha1_round/add_79/U119  ( .A(\sha1_round/f [5]), .ZN(
        \sha1_round/add_79/n32 ) );
  NAND2_X1 \sha1_round/add_79/U118  ( .A1(\sha1_round/f [23]), .A2(
        \sha1_round/k_23 ), .ZN(\sha1_round/add_79/n219 ) );
  NAND2_X1 \sha1_round/add_79/U117  ( .A1(\sha1_round/f [16]), .A2(
        \sha1_round/k_26 ), .ZN(\sha1_round/add_79/n233 ) );
  NAND2_X1 \sha1_round/add_79/U116  ( .A1(\sha1_round/f [19]), .A2(
        \sha1_round/k_26 ), .ZN(\sha1_round/add_79/n266 ) );
  NAND2_X1 \sha1_round/add_79/U115  ( .A1(\sha1_round/k_30 ), .A2(
        \sha1_round/f [8]), .ZN(\sha1_round/add_79/n100 ) );
  OR2_X2 \sha1_round/add_79/U114  ( .A1(\sha1_round/f [6]), .A2(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n85 ) );
  OR3_X1 \sha1_round/add_79/U113  ( .A1(\sha1_round/add_79/n132 ), .A2(
        \sha1_round/add_79/n26 ), .A3(\sha1_round/add_79/n168 ), .ZN(
        \sha1_round/add_79/n70 ) );
  NAND2_X2 \sha1_round/add_79/U112  ( .A1(\sha1_round/add_79/n203 ), .A2(
        \sha1_round/add_79/n204 ), .ZN(\sha1_round/add_79/n199 ) );
  XNOR2_X1 \sha1_round/add_79/U111  ( .A(\sha1_round/add_79/n228 ), .B(
        \sha1_round/add_79/n145 ), .ZN(\sha1_round/N275 ) );
  NOR3_X2 \sha1_round/add_79/U110  ( .A1(\sha1_round/add_79/n349 ), .A2(
        \sha1_round/add_79/n348 ), .A3(\sha1_round/add_79/n71 ), .ZN(
        \sha1_round/add_79/n31 ) );
  NAND2_X4 \sha1_round/add_79/U109  ( .A1(\sha1_round/add_79/n210 ), .A2(
        \sha1_round/add_79/n211 ), .ZN(\sha1_round/add_79/n207 ) );
  NAND2_X2 \sha1_round/add_79/U108  ( .A1(\sha1_round/f [12]), .A2(
        \sha1_round/n3300 ), .ZN(\sha1_round/add_79/n302 ) );
  INV_X4 \sha1_round/add_79/U107  ( .A(\sha1_round/add_79/n112 ), .ZN(
        \sha1_round/add_79/n45 ) );
  NOR2_X2 \sha1_round/add_79/U106  ( .A1(\sha1_round/add_79/n255 ), .A2(
        \sha1_round/add_79/n256 ), .ZN(\sha1_round/add_79/n254 ) );
  NAND2_X2 \sha1_round/add_79/U105  ( .A1(\sha1_round/add_79/n69 ), .A2(
        \sha1_round/add_79/n252 ), .ZN(\sha1_round/add_79/n244 ) );
  AND2_X2 \sha1_round/add_79/U104  ( .A1(\sha1_round/add_79/n252 ), .A2(
        \sha1_round/add_79/n243 ), .ZN(\sha1_round/add_79/n30 ) );
  OR2_X2 \sha1_round/add_79/U103  ( .A1(\sha1_round/add_79/n227 ), .A2(
        \sha1_round/add_79/n241 ), .ZN(\sha1_round/add_79/n29 ) );
  NAND2_X2 \sha1_round/add_79/U102  ( .A1(\sha1_round/add_79/n28 ), .A2(
        \sha1_round/add_79/n29 ), .ZN(\sha1_round/add_79/n229 ) );
  NAND2_X2 \sha1_round/add_79/U101  ( .A1(\sha1_round/add_79/n69 ), .A2(
        \sha1_round/add_79/n30 ), .ZN(\sha1_round/add_79/n28 ) );
  INV_X1 \sha1_round/add_79/U100  ( .A(\sha1_round/add_79/n27 ), .ZN(
        \sha1_round/add_79/n261 ) );
  NOR2_X2 \sha1_round/add_79/U99  ( .A1(\sha1_round/add_79/n262 ), .A2(
        \sha1_round/add_79/n260 ), .ZN(\sha1_round/add_79/n273 ) );
  NAND2_X2 \sha1_round/add_79/U98  ( .A1(\sha1_round/n2 ), .A2(
        \sha1_round/f [4]), .ZN(\sha1_round/add_79/n378 ) );
  INV_X4 \sha1_round/add_79/U97  ( .A(\sha1_round/add_79/n320 ), .ZN(
        \sha1_round/add_79/n51 ) );
  INV_X2 \sha1_round/add_79/U96  ( .A(\sha1_round/f [10]), .ZN(
        \sha1_round/add_79/n362 ) );
  NAND2_X2 \sha1_round/add_79/U95  ( .A1(\sha1_round/add_79/n360 ), .A2(
        \sha1_round/add_79/n361 ), .ZN(\sha1_round/add_79/n43 ) );
  NAND2_X2 \sha1_round/add_79/U94  ( .A1(\sha1_round/add_79/n99 ), .A2(
        \sha1_round/add_79/n100 ), .ZN(\sha1_round/add_79/n98 ) );
  NOR2_X4 \sha1_round/add_79/U93  ( .A1(\sha1_round/add_79/n97 ), .A2(
        \sha1_round/add_79/n98 ), .ZN(\sha1_round/add_79/n93 ) );
  NAND2_X2 \sha1_round/add_79/U92  ( .A1(\sha1_round/add_79/n325 ), .A2(
        \sha1_round/add_79/n327 ), .ZN(\sha1_round/add_79/n322 ) );
  NAND2_X2 \sha1_round/add_79/U91  ( .A1(\sha1_round/add_79/n320 ), .A2(
        \sha1_round/add_79/n321 ), .ZN(\sha1_round/add_79/n53 ) );
  NOR2_X2 \sha1_round/add_79/U90  ( .A1(\sha1_round/add_79/n316 ), .A2(
        \sha1_round/add_79/n317 ), .ZN(\sha1_round/add_79/n315 ) );
  NOR2_X2 \sha1_round/add_79/U89  ( .A1(\sha1_round/n517 ), .A2(
        \sha1_round/f [3]), .ZN(\sha1_round/add_79/n26 ) );
  OR2_X4 \sha1_round/add_79/U88  ( .A1(\sha1_round/f [24]), .A2(
        \sha1_round/add_79/n89 ), .ZN(\sha1_round/add_79/n25 ) );
  AND2_X4 \sha1_round/add_79/U87  ( .A1(\sha1_round/add_79/n340 ), .A2(
        \sha1_round/add_79/n339 ), .ZN(\sha1_round/add_79/n23 ) );
  AND2_X4 \sha1_round/add_79/U86  ( .A1(\sha1_round/add_79/n152 ), .A2(
        \sha1_round/add_79/n184 ), .ZN(\sha1_round/add_79/n22 ) );
  AND2_X4 \sha1_round/add_79/U85  ( .A1(\sha1_round/add_79/n366 ), .A2(
        \sha1_round/add_79/n110 ), .ZN(\sha1_round/add_79/n21 ) );
  OR2_X4 \sha1_round/add_79/U84  ( .A1(\sha1_round/add_79/n334 ), .A2(
        \sha1_round/add_79/n318 ), .ZN(\sha1_round/add_79/n20 ) );
  OR2_X4 \sha1_round/add_79/U83  ( .A1(\sha1_round/add_79/n318 ), .A2(
        \sha1_round/add_79/n302 ), .ZN(\sha1_round/add_79/n19 ) );
  OR2_X4 \sha1_round/add_79/U82  ( .A1(\sha1_round/add_79/n118 ), .A2(
        \sha1_round/add_79/n80 ), .ZN(\sha1_round/add_79/n18 ) );
  OR2_X4 \sha1_round/add_79/U81  ( .A1(\sha1_round/add_79/n26 ), .A2(
        \sha1_round/add_79/n370 ), .ZN(\sha1_round/add_79/n17 ) );
  OR2_X4 \sha1_round/add_79/U80  ( .A1(\sha1_round/add_79/n318 ), .A2(
        \sha1_round/add_79/n330 ), .ZN(\sha1_round/add_79/n16 ) );
  AND2_X4 \sha1_round/add_79/U79  ( .A1(\sha1_round/add_79/n252 ), .A2(
        \sha1_round/add_79/n240 ), .ZN(\sha1_round/add_79/n15 ) );
  AND2_X4 \sha1_round/add_79/U78  ( .A1(\sha1_round/add_79/n96 ), .A2(
        \sha1_round/add_79/n100 ), .ZN(\sha1_round/add_79/n14 ) );
  OR2_X2 \sha1_round/add_79/U77  ( .A1(\sha1_round/add_79/n79 ), .A2(
        \sha1_round/add_79/n278 ), .ZN(\sha1_round/add_79/n12 ) );
  AND2_X4 \sha1_round/add_79/U76  ( .A1(\sha1_round/add_79/n323 ), .A2(
        \sha1_round/add_79/n19 ), .ZN(\sha1_round/add_79/n11 ) );
  INV_X1 \sha1_round/add_79/U75  ( .A(\sha1_round/k_27 ), .ZN(
        \sha1_round/add_79/n55 ) );
  OR2_X4 \sha1_round/add_79/U74  ( .A1(\sha1_round/f [4]), .A2(\sha1_round/n2 ), .ZN(\sha1_round/add_79/n8 ) );
  NAND2_X1 \sha1_round/add_79/U73  ( .A1(\sha1_round/add_79/n119 ), .A2(
        \sha1_round/add_79/n8 ), .ZN(\sha1_round/add_79/n126 ) );
  NAND2_X1 \sha1_round/add_79/U72  ( .A1(\sha1_round/f [2]), .A2(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n371 ) );
  NOR2_X2 \sha1_round/add_79/U71  ( .A1(\sha1_round/add_79/n26 ), .A2(
        \sha1_round/add_79/n371 ), .ZN(\sha1_round/add_79/n308 ) );
  AND2_X2 \sha1_round/add_79/U70  ( .A1(\sha1_round/add_79/n302 ), .A2(
        \sha1_round/add_79/n303 ), .ZN(\sha1_round/add_79/n13 ) );
  NAND2_X1 \sha1_round/add_79/U69  ( .A1(\sha1_round/add_79/n332 ), .A2(
        \sha1_round/add_79/n303 ), .ZN(\sha1_round/add_79/n331 ) );
  NOR2_X2 \sha1_round/add_79/U68  ( .A1(\sha1_round/add_79/n67 ), .A2(
        \sha1_round/add_79/n331 ), .ZN(\sha1_round/add_79/n329 ) );
  NAND2_X1 \sha1_round/add_79/U67  ( .A1(\sha1_round/f [14]), .A2(
        \sha1_round/k_30 ), .ZN(\sha1_round/add_79/n294 ) );
  NOR2_X1 \sha1_round/add_79/U66  ( .A1(\sha1_round/add_79/n95 ), .A2(
        \sha1_round/add_79/n349 ), .ZN(\sha1_round/add_79/n94 ) );
  INV_X1 \sha1_round/add_79/U65  ( .A(\sha1_round/add_79/n145 ), .ZN(
        \sha1_round/add_79/n185 ) );
  NAND2_X1 \sha1_round/add_79/U64  ( .A1(\sha1_round/add_79/n106 ), .A2(
        \sha1_round/add_79/n107 ), .ZN(\sha1_round/add_79/n105 ) );
  NOR2_X2 \sha1_round/add_79/U63  ( .A1(\sha1_round/add_79/n329 ), .A2(
        \sha1_round/add_79/n16 ), .ZN(\sha1_round/add_79/n324 ) );
  NOR2_X2 \sha1_round/add_79/U62  ( .A1(\sha1_round/f [14]), .A2(
        \sha1_round/k_30 ), .ZN(\sha1_round/add_79/n317 ) );
  NAND2_X2 \sha1_round/add_79/U61  ( .A1(\sha1_round/k_26 ), .A2(
        \sha1_round/f [20]), .ZN(\sha1_round/add_79/n258 ) );
  NAND2_X2 \sha1_round/add_79/U60  ( .A1(\sha1_round/add_79/n109 ), .A2(
        \sha1_round/add_79/n110 ), .ZN(\sha1_round/add_79/n104 ) );
  NOR2_X2 \sha1_round/add_79/U59  ( .A1(\sha1_round/f [1]), .A2(
        \sha1_round/n824 ), .ZN(\sha1_round/add_79/n168 ) );
  NAND2_X2 \sha1_round/add_79/U58  ( .A1(\sha1_round/add_79/n293 ), .A2(
        \sha1_round/add_79/n233 ), .ZN(\sha1_round/add_79/n232 ) );
  NAND2_X2 \sha1_round/add_79/U57  ( .A1(\sha1_round/add_79/n239 ), .A2(
        \sha1_round/add_79/n230 ), .ZN(\sha1_round/add_79/n224 ) );
  NOR2_X2 \sha1_round/add_79/U56  ( .A1(\sha1_round/add_79/n190 ), .A2(
        \sha1_round/add_79/n183 ), .ZN(\sha1_round/add_79/n188 ) );
  NAND3_X2 \sha1_round/add_79/U55  ( .A1(\sha1_round/f [18]), .A2(
        \sha1_round/add_79/n259 ), .A3(\sha1_round/add_79/n27 ), .ZN(
        \sha1_round/add_79/n251 ) );
  INV_X4 \sha1_round/add_79/U54  ( .A(\sha1_round/add_79/n360 ), .ZN(
        \sha1_round/add_79/n41 ) );
  NAND2_X2 \sha1_round/add_79/U53  ( .A1(\sha1_round/add_79/n364 ), .A2(
        \sha1_round/add_79/n365 ), .ZN(\sha1_round/add_79/n363 ) );
  NOR2_X2 \sha1_round/add_79/U52  ( .A1(\sha1_round/add_79/n132 ), .A2(
        \sha1_round/add_79/n133 ), .ZN(\sha1_round/add_79/n130 ) );
  NOR2_X2 \sha1_round/add_79/U51  ( .A1(\sha1_round/add_79/n130 ), .A2(
        \sha1_round/add_79/n131 ), .ZN(\sha1_round/add_79/n127 ) );
  INV_X4 \sha1_round/add_79/U50  ( .A(\sha1_round/add_79/n349 ), .ZN(
        \sha1_round/add_79/n365 ) );
  NOR2_X2 \sha1_round/add_79/U49  ( .A1(\sha1_round/f [7]), .A2(
        \sha1_round/k_27 ), .ZN(\sha1_round/add_79/n373 ) );
  NAND3_X2 \sha1_round/add_79/U48  ( .A1(\sha1_round/add_79/n372 ), .A2(
        \sha1_round/add_79/n8 ), .A3(\sha1_round/add_79/n121 ), .ZN(
        \sha1_round/add_79/n108 ) );
  NOR2_X2 \sha1_round/add_79/U47  ( .A1(\sha1_round/add_79/n379 ), .A2(
        \sha1_round/add_79/n373 ), .ZN(\sha1_round/add_79/n372 ) );
  NOR2_X1 \sha1_round/add_79/U46  ( .A1(\sha1_round/add_79/n81 ), .A2(
        \sha1_round/add_79/n379 ), .ZN(\sha1_round/add_79/n116 ) );
  INV_X4 \sha1_round/add_79/U45  ( .A(\sha1_round/add_79/n108 ), .ZN(
        \sha1_round/add_79/n106 ) );
  NOR2_X4 \sha1_round/add_79/U44  ( .A1(\sha1_round/f [6]), .A2(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n379 ) );
  INV_X2 \sha1_round/add_79/U43  ( .A(\sha1_round/add_79/n287 ), .ZN(
        \sha1_round/add_79/n286 ) );
  NAND2_X1 \sha1_round/add_79/U42  ( .A1(\sha1_round/add_79/n287 ), .A2(
        \sha1_round/add_79/n293 ), .ZN(\sha1_round/add_79/n290 ) );
  NOR2_X1 \sha1_round/add_79/U41  ( .A1(\sha1_round/n517 ), .A2(
        \sha1_round/f [3]), .ZN(\sha1_round/add_79/n84 ) );
  NAND2_X4 \sha1_round/add_79/U40  ( .A1(\sha1_round/add_79/n285 ), .A2(
        \sha1_round/add_79/n284 ), .ZN(\sha1_round/add_79/n282 ) );
  NAND2_X4 \sha1_round/add_79/U39  ( .A1(\sha1_round/add_79/n5 ), .A2(
        \sha1_round/add_79/n338 ), .ZN(\sha1_round/add_79/n336 ) );
  NAND3_X4 \sha1_round/add_79/U38  ( .A1(\sha1_round/add_79/n240 ), .A2(
        \sha1_round/add_79/n241 ), .A3(\sha1_round/add_79/n242 ), .ZN(
        \sha1_round/add_79/n237 ) );
  NOR3_X4 \sha1_round/add_79/U37  ( .A1(\sha1_round/add_79/n237 ), .A2(
        \sha1_round/add_79/n12 ), .A3(\sha1_round/add_79/n238 ), .ZN(
        \sha1_round/add_79/n234 ) );
  NAND2_X1 \sha1_round/add_79/U36  ( .A1(\sha1_round/f [27]), .A2(
        \sha1_round/k_27 ), .ZN(\sha1_round/add_79/n152 ) );
  NAND2_X1 \sha1_round/add_79/U35  ( .A1(\sha1_round/f [25]), .A2(
        \sha1_round/k_27 ), .ZN(\sha1_round/add_79/n198 ) );
  OR2_X2 \sha1_round/add_79/U34  ( .A1(\sha1_round/add_79/n317 ), .A2(
        \sha1_round/add_79/n296 ), .ZN(\sha1_round/add_79/n24 ) );
  NOR2_X1 \sha1_round/add_79/U33  ( .A1(\sha1_round/f [13]), .A2(
        \sha1_round/k[13] ), .ZN(\sha1_round/add_79/n318 ) );
  OR2_X4 \sha1_round/add_79/U32  ( .A1(\sha1_round/f [19]), .A2(
        \sha1_round/k_26 ), .ZN(\sha1_round/add_79/n27 ) );
  INV_X1 \sha1_round/add_79/U31  ( .A(\sha1_round/add_79/n340 ), .ZN(
        \sha1_round/add_79/n347 ) );
  NAND2_X2 \sha1_round/add_79/U30  ( .A1(\sha1_round/add_79/n286 ), .A2(
        \sha1_round/add_79/n280 ), .ZN(\sha1_round/add_79/n285 ) );
  NAND2_X2 \sha1_round/add_79/U29  ( .A1(\sha1_round/add_79/n358 ), .A2(
        \sha1_round/add_79/n357 ), .ZN(\sha1_round/add_79/n356 ) );
  AND2_X4 \sha1_round/add_79/U28  ( .A1(\sha1_round/add_79/n100 ), .A2(
        \sha1_round/add_79/n99 ), .ZN(\sha1_round/add_79/n4 ) );
  INV_X4 \sha1_round/add_79/U27  ( .A(\sha1_round/add_79/n281 ), .ZN(
        \sha1_round/N269 ) );
  INV_X4 \sha1_round/add_79/U26  ( .A(\sha1_round/add_79/n321 ), .ZN(
        \sha1_round/add_79/n52 ) );
  NAND2_X2 \sha1_round/add_79/U25  ( .A1(\sha1_round/add_79/n335 ), .A2(
        \sha1_round/add_79/n302 ), .ZN(\sha1_round/add_79/n333 ) );
  NAND3_X2 \sha1_round/add_79/U24  ( .A1(\sha1_round/add_79/n225 ), .A2(
        \sha1_round/add_79/n229 ), .A3(\sha1_round/add_79/n224 ), .ZN(
        \sha1_round/add_79/n49 ) );
  NAND2_X2 \sha1_round/add_79/U23  ( .A1(\sha1_round/add_79/n328 ), .A2(
        \sha1_round/add_79/n11 ), .ZN(\sha1_round/add_79/n325 ) );
  NAND2_X2 \sha1_round/add_79/U22  ( .A1(\sha1_round/add_79/n367 ), .A2(
        \sha1_round/add_79/n368 ), .ZN(\sha1_round/add_79/n63 ) );
  NAND2_X2 \sha1_round/add_79/U21  ( .A1(\sha1_round/add_79/n368 ), .A2(
        \sha1_round/add_79/n367 ), .ZN(\sha1_round/add_79/n107 ) );
  NAND2_X2 \sha1_round/add_79/U20  ( .A1(\sha1_round/add_79/n359 ), .A2(
        \sha1_round/add_79/n340 ), .ZN(\sha1_round/add_79/n71 ) );
  NOR2_X2 \sha1_round/add_79/U19  ( .A1(\sha1_round/add_79/n369 ), .A2(
        \sha1_round/add_79/n62 ), .ZN(\sha1_round/add_79/n368 ) );
  NAND2_X2 \sha1_round/add_79/U18  ( .A1(\sha1_round/add_79/n366 ), .A2(
        \sha1_round/add_79/n106 ), .ZN(\sha1_round/add_79/n60 ) );
  NAND2_X2 \sha1_round/add_79/U17  ( .A1(\sha1_round/add_79/n288 ), .A2(
        \sha1_round/add_79/n289 ), .ZN(\sha1_round/add_79/n293 ) );
  NAND2_X2 \sha1_round/add_79/U16  ( .A1(\sha1_round/f [0]), .A2(
        \sha1_round/k_23 ), .ZN(\sha1_round/add_79/n312 ) );
  NAND3_X4 \sha1_round/add_79/U15  ( .A1(\sha1_round/add_79/n274 ), .A2(
        \sha1_round/add_79/n275 ), .A3(\sha1_round/add_79/n276 ), .ZN(
        \sha1_round/add_79/n250 ) );
  NOR2_X4 \sha1_round/add_79/U14  ( .A1(\sha1_round/add_79/n114 ), .A2(
        \sha1_round/add_79/n81 ), .ZN(\sha1_round/add_79/n112 ) );
  INV_X2 \sha1_round/add_79/U13  ( .A(\sha1_round/add_79/n31 ), .ZN(
        \sha1_round/add_79/n319 ) );
  NAND2_X4 \sha1_round/add_79/U12  ( .A1(\sha1_round/add_79/n363 ), .A2(
        \sha1_round/add_79/n96 ), .ZN(\sha1_round/add_79/n360 ) );
  NOR3_X2 \sha1_round/add_79/U11  ( .A1(\sha1_round/add_79/n378 ), .A2(
        \sha1_round/add_79/n379 ), .A3(\sha1_round/add_79/n380 ), .ZN(
        \sha1_round/add_79/n377 ) );
  NAND2_X1 \sha1_round/add_79/U10  ( .A1(\sha1_round/add_79/n8 ), .A2(
        \sha1_round/add_79/n63 ), .ZN(\sha1_round/add_79/n125 ) );
  AND3_X4 \sha1_round/add_79/U9  ( .A1(\sha1_round/add_79/n107 ), .A2(
        \sha1_round/add_79/n31 ), .A3(\sha1_round/add_79/n106 ), .ZN(
        \sha1_round/add_79/n67 ) );
  INV_X8 \sha1_round/add_79/U8  ( .A(\sha1_round/add_79/n351 ), .ZN(
        \sha1_round/N263 ) );
  CLKBUF_X2 \sha1_round/add_79/U7  ( .A(\sha1_round/f [6]), .Z(
        \sha1_round/add_79/n2 ) );
  NOR2_X2 \sha1_round/add_79/U6  ( .A1(\sha1_round/add_79/n17 ), .A2(
        \sha1_round/add_79/n132 ), .ZN(\sha1_round/add_79/n62 ) );
  AND2_X2 \sha1_round/add_79/U5  ( .A1(\sha1_round/add_79/n303 ), .A2(
        \sha1_round/add_79/n332 ), .ZN(\sha1_round/add_79/n5 ) );
  AND2_X4 \sha1_round/add_79/U4  ( .A1(\sha1_round/add_79/n205 ), .A2(
        \sha1_round/add_79/n193 ), .ZN(\sha1_round/add_79/n1 ) );
  NOR2_X4 \sha1_round/add_79/U3  ( .A1(\sha1_round/f [2]), .A2(
        \sha1_round/add_79/n87 ), .ZN(\sha1_round/add_79/n132 ) );
  NAND2_X2 \sha1_round/add_79/U2  ( .A1(\sha1_round/add_79/n356 ), .A2(
        \sha1_round/add_79/n344 ), .ZN(\sha1_round/add_79/n352 ) );
  NAND2_X2 \sha1_round/add_79_2/U405  ( .A1(w[0]), .A2(rnd_q[0]), .ZN(
        \sha1_round/add_79_2/n223 ) );
  INV_X4 \sha1_round/add_79_2/U404  ( .A(\sha1_round/add_79_2/n223 ), .ZN(
        \sha1_round/add_79_2/n299 ) );
  NAND2_X2 \sha1_round/add_79_2/U403  ( .A1(w[9]), .A2(rnd_q[9]), .ZN(
        \sha1_round/add_79_2/n349 ) );
  INV_X4 \sha1_round/add_79_2/U402  ( .A(\sha1_round/add_79_2/n349 ), .ZN(
        \sha1_round/add_79_2/n40 ) );
  INV_X4 \sha1_round/add_79_2/U401  ( .A(\sha1_round/add_79_2/n83 ), .ZN(
        \sha1_round/add_79_2/n298 ) );
  NAND2_X2 \sha1_round/add_79_2/U400  ( .A1(rnd_q[2]), .A2(w[2]), .ZN(
        \sha1_round/add_79_2/n374 ) );
  INV_X4 \sha1_round/add_79_2/U399  ( .A(\sha1_round/add_79_2/n107 ), .ZN(
        \sha1_round/add_79_2/n370 ) );
  NAND2_X2 \sha1_round/add_79_2/U398  ( .A1(w[3]), .A2(rnd_q[3]), .ZN(
        \sha1_round/add_79_2/n72 ) );
  NAND2_X2 \sha1_round/add_79_2/U397  ( .A1(w[0]), .A2(rnd_q[0]), .ZN(
        \sha1_round/add_79_2/n372 ) );
  NAND2_X2 \sha1_round/add_79_2/U396  ( .A1(w[1]), .A2(rnd_q[1]), .ZN(
        \sha1_round/add_79_2/n373 ) );
  NAND2_X2 \sha1_round/add_79_2/U395  ( .A1(\sha1_round/add_79_2/n372 ), .A2(
        \sha1_round/add_79_2/n373 ), .ZN(\sha1_round/add_79_2/n369 ) );
  INV_X4 \sha1_round/add_79_2/U394  ( .A(\sha1_round/add_79_2/n61 ), .ZN(
        \sha1_round/add_79_2/n363 ) );
  INV_X4 \sha1_round/add_79_2/U393  ( .A(w[4]), .ZN(\sha1_round/add_79_2/n366 ) );
  INV_X4 \sha1_round/add_79_2/U392  ( .A(rnd_q[4]), .ZN(
        \sha1_round/add_79_2/n367 ) );
  NAND2_X2 \sha1_round/add_79_2/U391  ( .A1(\sha1_round/add_79_2/n366 ), .A2(
        \sha1_round/add_79_2/n367 ), .ZN(\sha1_round/add_79_2/n71 ) );
  INV_X4 \sha1_round/add_79_2/U390  ( .A(\sha1_round/add_79_2/n262 ), .ZN(
        \sha1_round/add_79_2/n56 ) );
  NAND2_X2 \sha1_round/add_79_2/U389  ( .A1(rnd_q[6]), .A2(w[6]), .ZN(
        \sha1_round/add_79_2/n362 ) );
  INV_X4 \sha1_round/add_79_2/U388  ( .A(\sha1_round/add_79_2/n276 ), .ZN(
        \sha1_round/add_79_2/n358 ) );
  NAND2_X2 \sha1_round/add_79_2/U387  ( .A1(w[7]), .A2(rnd_q[7]), .ZN(
        \sha1_round/add_79_2/n269 ) );
  NAND2_X2 \sha1_round/add_79_2/U386  ( .A1(w[4]), .A2(rnd_q[4]), .ZN(
        \sha1_round/add_79_2/n81 ) );
  NAND2_X2 \sha1_round/add_79_2/U385  ( .A1(w[5]), .A2(rnd_q[5]), .ZN(
        \sha1_round/add_79_2/n69 ) );
  NAND2_X2 \sha1_round/add_79_2/U384  ( .A1(\sha1_round/add_79_2/n81 ), .A2(
        \sha1_round/add_79_2/n69 ), .ZN(\sha1_round/add_79_2/n360 ) );
  INV_X4 \sha1_round/add_79_2/U383  ( .A(\sha1_round/add_79_2/n47 ), .ZN(
        \sha1_round/add_79_2/n321 ) );
  NAND2_X2 \sha1_round/add_79_2/U382  ( .A1(w[8]), .A2(rnd_q[8]), .ZN(
        \sha1_round/add_79_2/n52 ) );
  NAND2_X2 \sha1_round/add_79_2/U381  ( .A1(\sha1_round/add_79_2/n321 ), .A2(
        \sha1_round/add_79_2/n52 ), .ZN(\sha1_round/add_79_2/n357 ) );
  XNOR2_X2 \sha1_round/add_79_2/U380  ( .A(\sha1_round/add_79_2/n352 ), .B(
        \sha1_round/add_79_2/n353 ), .ZN(\sha1_round/N294 ) );
  INV_X4 \sha1_round/add_79_2/U379  ( .A(\sha1_round/add_79_2/n285 ), .ZN(
        \sha1_round/add_79_2/n340 ) );
  XNOR2_X2 \sha1_round/add_79_2/U378  ( .A(\sha1_round/add_79_2/n344 ), .B(
        \sha1_round/add_79_2/n345 ), .ZN(\sha1_round/N295 ) );
  INV_X4 \sha1_round/add_79_2/U377  ( .A(w[12]), .ZN(
        \sha1_round/add_79_2/n342 ) );
  INV_X4 \sha1_round/add_79_2/U376  ( .A(rnd_q[12]), .ZN(
        \sha1_round/add_79_2/n343 ) );
  NAND2_X2 \sha1_round/add_79_2/U375  ( .A1(\sha1_round/add_79_2/n342 ), .A2(
        \sha1_round/add_79_2/n343 ), .ZN(\sha1_round/add_79_2/n301 ) );
  NAND2_X2 \sha1_round/add_79_2/U374  ( .A1(w[12]), .A2(rnd_q[12]), .ZN(
        \sha1_round/add_79_2/n292 ) );
  NAND2_X2 \sha1_round/add_79_2/U373  ( .A1(\sha1_round/add_79_2/n301 ), .A2(
        \sha1_round/add_79_2/n292 ), .ZN(\sha1_round/add_79_2/n329 ) );
  INV_X4 \sha1_round/add_79_2/U372  ( .A(\sha1_round/add_79_2/n44 ), .ZN(
        \sha1_round/add_79_2/n338 ) );
  INV_X4 \sha1_round/add_79_2/U371  ( .A(\sha1_round/add_79_2/n264 ), .ZN(
        \sha1_round/add_79_2/n268 ) );
  NAND2_X2 \sha1_round/add_79_2/U370  ( .A1(\sha1_round/add_79_2/n268 ), .A2(
        \sha1_round/add_79_2/n47 ), .ZN(\sha1_round/add_79_2/n330 ) );
  INV_X4 \sha1_round/add_79_2/U369  ( .A(\sha1_round/add_79_2/n41 ), .ZN(
        \sha1_round/add_79_2/n336 ) );
  INV_X4 \sha1_round/add_79_2/U368  ( .A(\sha1_round/add_79_2/n335 ), .ZN(
        \sha1_round/add_79_2/n337 ) );
  NAND4_X2 \sha1_round/add_79_2/U367  ( .A1(w[8]), .A2(rnd_q[8]), .A3(
        \sha1_round/add_79_2/n336 ), .A4(\sha1_round/add_79_2/n337 ), .ZN(
        \sha1_round/add_79_2/n332 ) );
  NAND2_X2 \sha1_round/add_79_2/U366  ( .A1(\sha1_round/add_79_2/n286 ), .A2(
        \sha1_round/add_79_2/n285 ), .ZN(\sha1_round/add_79_2/n322 ) );
  INV_X4 \sha1_round/add_79_2/U365  ( .A(\sha1_round/add_79_2/n49 ), .ZN(
        \sha1_round/add_79_2/n273 ) );
  NAND2_X2 \sha1_round/add_79_2/U364  ( .A1(\sha1_round/add_79_2/n273 ), .A2(
        \sha1_round/add_79_2/n268 ), .ZN(\sha1_round/add_79_2/n331 ) );
  XNOR2_X2 \sha1_round/add_79_2/U363  ( .A(\sha1_round/add_79_2/n329 ), .B(
        \sha1_round/add_79_2/n328 ), .ZN(\sha1_round/N296 ) );
  NAND2_X2 \sha1_round/add_79_2/U362  ( .A1(\sha1_round/add_79_2/n328 ), .A2(
        \sha1_round/add_79_2/n301 ), .ZN(\sha1_round/add_79_2/n327 ) );
  NAND2_X2 \sha1_round/add_79_2/U361  ( .A1(\sha1_round/add_79_2/n327 ), .A2(
        \sha1_round/add_79_2/n292 ), .ZN(\sha1_round/add_79_2/n323 ) );
  NAND2_X2 \sha1_round/add_79_2/U360  ( .A1(w[13]), .A2(rnd_q[13]), .ZN(
        \sha1_round/add_79_2/n279 ) );
  INV_X4 \sha1_round/add_79_2/U359  ( .A(w[13]), .ZN(
        \sha1_round/add_79_2/n325 ) );
  INV_X4 \sha1_round/add_79_2/U358  ( .A(rnd_q[13]), .ZN(
        \sha1_round/add_79_2/n326 ) );
  NAND2_X2 \sha1_round/add_79_2/U357  ( .A1(\sha1_round/add_79_2/n325 ), .A2(
        \sha1_round/add_79_2/n326 ), .ZN(\sha1_round/add_79_2/n300 ) );
  NAND2_X2 \sha1_round/add_79_2/U356  ( .A1(\sha1_round/add_79_2/n279 ), .A2(
        \sha1_round/add_79_2/n300 ), .ZN(\sha1_round/add_79_2/n324 ) );
  XNOR2_X2 \sha1_round/add_79_2/U355  ( .A(\sha1_round/add_79_2/n323 ), .B(
        \sha1_round/add_79_2/n324 ), .ZN(\sha1_round/N297 ) );
  INV_X4 \sha1_round/add_79_2/U354  ( .A(\sha1_round/add_79_2/n322 ), .ZN(
        \sha1_round/add_79_2/n319 ) );
  INV_X4 \sha1_round/add_79_2/U353  ( .A(\sha1_round/add_79_2/n76 ), .ZN(
        \sha1_round/add_79_2/n275 ) );
  NAND2_X2 \sha1_round/add_79_2/U352  ( .A1(\sha1_round/add_79_2/n317 ), .A2(
        \sha1_round/add_79_2/n318 ), .ZN(\sha1_round/add_79_2/n316 ) );
  NAND2_X2 \sha1_round/add_79_2/U351  ( .A1(\sha1_round/add_79_2/n315 ), .A2(
        \sha1_round/add_79_2/n316 ), .ZN(\sha1_round/add_79_2/n314 ) );
  NAND2_X2 \sha1_round/add_79_2/U350  ( .A1(\sha1_round/add_79_2/n314 ), .A2(
        \sha1_round/add_79_2/n301 ), .ZN(\sha1_round/add_79_2/n307 ) );
  NAND2_X2 \sha1_round/add_79_2/U349  ( .A1(\sha1_round/add_79_2/n307 ), .A2(
        \sha1_round/add_79_2/n292 ), .ZN(\sha1_round/add_79_2/n313 ) );
  NAND2_X2 \sha1_round/add_79_2/U348  ( .A1(\sha1_round/add_79_2/n313 ), .A2(
        \sha1_round/add_79_2/n300 ), .ZN(\sha1_round/add_79_2/n312 ) );
  NAND2_X2 \sha1_round/add_79_2/U347  ( .A1(\sha1_round/add_79_2/n279 ), .A2(
        \sha1_round/add_79_2/n312 ), .ZN(\sha1_round/add_79_2/n308 ) );
  INV_X4 \sha1_round/add_79_2/U346  ( .A(w[14]), .ZN(
        \sha1_round/add_79_2/n310 ) );
  INV_X4 \sha1_round/add_79_2/U345  ( .A(rnd_q[14]), .ZN(
        \sha1_round/add_79_2/n311 ) );
  NAND2_X2 \sha1_round/add_79_2/U344  ( .A1(\sha1_round/add_79_2/n310 ), .A2(
        \sha1_round/add_79_2/n311 ), .ZN(\sha1_round/add_79_2/n281 ) );
  NAND2_X2 \sha1_round/add_79_2/U343  ( .A1(w[14]), .A2(rnd_q[14]), .ZN(
        \sha1_round/add_79_2/n280 ) );
  NAND2_X2 \sha1_round/add_79_2/U342  ( .A1(\sha1_round/add_79_2/n281 ), .A2(
        \sha1_round/add_79_2/n280 ), .ZN(\sha1_round/add_79_2/n309 ) );
  XNOR2_X2 \sha1_round/add_79_2/U341  ( .A(\sha1_round/add_79_2/n308 ), .B(
        \sha1_round/add_79_2/n309 ), .ZN(\sha1_round/N298 ) );
  INV_X4 \sha1_round/add_79_2/U340  ( .A(\sha1_round/add_79_2/n280 ), .ZN(
        \sha1_round/add_79_2/n306 ) );
  NAND2_X2 \sha1_round/add_79_2/U339  ( .A1(w[15]), .A2(rnd_q[15]), .ZN(
        \sha1_round/add_79_2/n284 ) );
  INV_X4 \sha1_round/add_79_2/U338  ( .A(w[15]), .ZN(
        \sha1_round/add_79_2/n303 ) );
  INV_X4 \sha1_round/add_79_2/U337  ( .A(rnd_q[15]), .ZN(
        \sha1_round/add_79_2/n304 ) );
  NAND2_X2 \sha1_round/add_79_2/U336  ( .A1(\sha1_round/add_79_2/n303 ), .A2(
        \sha1_round/add_79_2/n304 ), .ZN(\sha1_round/add_79_2/n282 ) );
  NAND2_X2 \sha1_round/add_79_2/U335  ( .A1(\sha1_round/add_79_2/n284 ), .A2(
        \sha1_round/add_79_2/n282 ), .ZN(\sha1_round/add_79_2/n302 ) );
  NAND2_X2 \sha1_round/add_79_2/U334  ( .A1(w[16]), .A2(rnd_q[16]), .ZN(
        \sha1_round/add_79_2/n251 ) );
  NAND2_X2 \sha1_round/add_79_2/U333  ( .A1(\sha1_round/add_79_2/n251 ), .A2(
        \sha1_round/add_79_2/n253 ), .ZN(\sha1_round/add_79_2/n254 ) );
  NAND2_X2 \sha1_round/add_79_2/U332  ( .A1(\sha1_round/add_79_2/n261 ), .A2(
        \sha1_round/add_79_2/n268 ), .ZN(\sha1_round/add_79_2/n294 ) );
  NAND2_X2 \sha1_round/add_79_2/U331  ( .A1(w[1]), .A2(rnd_q[1]), .ZN(
        \sha1_round/add_79_2/n108 ) );
  INV_X4 \sha1_round/add_79_2/U330  ( .A(\sha1_round/add_79_2/n108 ), .ZN(
        \sha1_round/add_79_2/n222 ) );
  NAND2_X2 \sha1_round/add_79_2/U329  ( .A1(\sha1_round/add_79_2/n296 ), .A2(
        \sha1_round/add_79_2/n273 ), .ZN(\sha1_round/add_79_2/n295 ) );
  NAND3_X2 \sha1_round/add_79_2/U328  ( .A1(\sha1_round/add_79_2/n261 ), .A2(
        \sha1_round/add_79_2/n273 ), .A3(\sha1_round/add_79_2/n293 ), .ZN(
        \sha1_round/add_79_2/n289 ) );
  INV_X4 \sha1_round/add_79_2/U327  ( .A(\sha1_round/add_79_2/n292 ), .ZN(
        \sha1_round/add_79_2/n291 ) );
  NAND2_X2 \sha1_round/add_79_2/U326  ( .A1(\sha1_round/add_79_2/n291 ), .A2(
        \sha1_round/add_79_2/n261 ), .ZN(\sha1_round/add_79_2/n290 ) );
  NAND2_X2 \sha1_round/add_79_2/U325  ( .A1(\sha1_round/add_79_2/n289 ), .A2(
        \sha1_round/add_79_2/n290 ), .ZN(\sha1_round/add_79_2/n288 ) );
  NAND2_X2 \sha1_round/add_79_2/U324  ( .A1(\sha1_round/add_79_2/n279 ), .A2(
        \sha1_round/add_79_2/n280 ), .ZN(\sha1_round/add_79_2/n278 ) );
  NAND2_X2 \sha1_round/add_79_2/U323  ( .A1(\sha1_round/add_79_2/n277 ), .A2(
        \sha1_round/add_79_2/n278 ), .ZN(\sha1_round/add_79_2/n270 ) );
  NAND3_X2 \sha1_round/add_79_2/U322  ( .A1(\sha1_round/add_79_2/n276 ), .A2(
        \sha1_round/add_79_2/n261 ), .A3(\sha1_round/add_79_2/n268 ), .ZN(
        \sha1_round/add_79_2/n271 ) );
  NAND3_X2 \sha1_round/add_79_2/U321  ( .A1(\sha1_round/add_79_2/n261 ), .A2(
        \sha1_round/add_79_2/n273 ), .A3(\sha1_round/add_79_2/n274 ), .ZN(
        \sha1_round/add_79_2/n272 ) );
  NAND3_X2 \sha1_round/add_79_2/U320  ( .A1(\sha1_round/add_79_2/n270 ), .A2(
        \sha1_round/add_79_2/n271 ), .A3(\sha1_round/add_79_2/n272 ), .ZN(
        \sha1_round/add_79_2/n257 ) );
  INV_X4 \sha1_round/add_79_2/U319  ( .A(\sha1_round/add_79_2/n269 ), .ZN(
        \sha1_round/add_79_2/n57 ) );
  NAND3_X2 \sha1_round/add_79_2/U318  ( .A1(\sha1_round/add_79_2/n57 ), .A2(
        \sha1_round/add_79_2/n261 ), .A3(\sha1_round/add_79_2/n268 ), .ZN(
        \sha1_round/add_79_2/n259 ) );
  NAND2_X2 \sha1_round/add_79_2/U317  ( .A1(\sha1_round/add_79_2/n81 ), .A2(
        \sha1_round/add_79_2/n69 ), .ZN(\sha1_round/add_79_2/n267 ) );
  NAND2_X2 \sha1_round/add_79_2/U316  ( .A1(\sha1_round/add_79_2/n266 ), .A2(
        \sha1_round/add_79_2/n267 ), .ZN(\sha1_round/add_79_2/n265 ) );
  NAND2_X2 \sha1_round/add_79_2/U315  ( .A1(\sha1_round/add_79_2/n259 ), .A2(
        \sha1_round/add_79_2/n260 ), .ZN(\sha1_round/add_79_2/n258 ) );
  NOR2_X2 \sha1_round/add_79_2/U314  ( .A1(\sha1_round/add_79_2/n257 ), .A2(
        \sha1_round/add_79_2/n258 ), .ZN(\sha1_round/add_79_2/n256 ) );
  XNOR2_X2 \sha1_round/add_79_2/U313  ( .A(\sha1_round/add_79_2/n254 ), .B(
        \sha1_round/add_79_2/n118 ), .ZN(\sha1_round/N300 ) );
  INV_X4 \sha1_round/add_79_2/U312  ( .A(\sha1_round/add_79_2/n231 ), .ZN(
        \sha1_round/add_79_2/n253 ) );
  NAND2_X2 \sha1_round/add_79_2/U311  ( .A1(\sha1_round/add_79_2/n118 ), .A2(
        \sha1_round/add_79_2/n253 ), .ZN(\sha1_round/add_79_2/n252 ) );
  NAND2_X2 \sha1_round/add_79_2/U310  ( .A1(\sha1_round/add_79_2/n251 ), .A2(
        \sha1_round/add_79_2/n252 ), .ZN(\sha1_round/add_79_2/n246 ) );
  INV_X4 \sha1_round/add_79_2/U309  ( .A(w[17]), .ZN(
        \sha1_round/add_79_2/n249 ) );
  INV_X4 \sha1_round/add_79_2/U308  ( .A(rnd_q[17]), .ZN(
        \sha1_round/add_79_2/n250 ) );
  NAND2_X2 \sha1_round/add_79_2/U307  ( .A1(\sha1_round/add_79_2/n249 ), .A2(
        \sha1_round/add_79_2/n250 ), .ZN(\sha1_round/add_79_2/n244 ) );
  INV_X4 \sha1_round/add_79_2/U306  ( .A(\sha1_round/add_79_2/n244 ), .ZN(
        \sha1_round/add_79_2/n233 ) );
  NAND2_X2 \sha1_round/add_79_2/U305  ( .A1(w[17]), .A2(rnd_q[17]), .ZN(
        \sha1_round/add_79_2/n243 ) );
  INV_X4 \sha1_round/add_79_2/U304  ( .A(\sha1_round/add_79_2/n243 ), .ZN(
        \sha1_round/add_79_2/n248 ) );
  INV_X4 \sha1_round/add_79_2/U303  ( .A(\sha1_round/add_79_2/n118 ), .ZN(
        \sha1_round/add_79_2/n245 ) );
  NAND2_X2 \sha1_round/add_79_2/U302  ( .A1(\sha1_round/add_79_2/n242 ), .A2(
        \sha1_round/add_79_2/n243 ), .ZN(\sha1_round/add_79_2/n237 ) );
  NAND2_X2 \sha1_round/add_79_2/U301  ( .A1(w[18]), .A2(rnd_q[18]), .ZN(
        \sha1_round/add_79_2/n236 ) );
  INV_X4 \sha1_round/add_79_2/U300  ( .A(w[18]), .ZN(
        \sha1_round/add_79_2/n239 ) );
  INV_X4 \sha1_round/add_79_2/U299  ( .A(rnd_q[18]), .ZN(
        \sha1_round/add_79_2/n240 ) );
  NAND2_X2 \sha1_round/add_79_2/U298  ( .A1(\sha1_round/add_79_2/n239 ), .A2(
        \sha1_round/add_79_2/n240 ), .ZN(\sha1_round/add_79_2/n234 ) );
  NAND2_X2 \sha1_round/add_79_2/U297  ( .A1(\sha1_round/add_79_2/n236 ), .A2(
        \sha1_round/add_79_2/n234 ), .ZN(\sha1_round/add_79_2/n238 ) );
  NAND2_X2 \sha1_round/add_79_2/U296  ( .A1(\sha1_round/add_79_2/n237 ), .A2(
        \sha1_round/add_79_2/n234 ), .ZN(\sha1_round/add_79_2/n235 ) );
  NAND2_X2 \sha1_round/add_79_2/U295  ( .A1(\sha1_round/add_79_2/n235 ), .A2(
        \sha1_round/add_79_2/n236 ), .ZN(\sha1_round/add_79_2/n185 ) );
  INV_X4 \sha1_round/add_79_2/U294  ( .A(\sha1_round/add_79_2/n185 ), .ZN(
        \sha1_round/add_79_2/n229 ) );
  INV_X4 \sha1_round/add_79_2/U293  ( .A(\sha1_round/add_79_2/n234 ), .ZN(
        \sha1_round/add_79_2/n232 ) );
  NAND2_X2 \sha1_round/add_79_2/U292  ( .A1(\sha1_round/add_79_2/n219 ), .A2(
        \sha1_round/add_79_2/n118 ), .ZN(\sha1_round/add_79_2/n230 ) );
  NAND2_X2 \sha1_round/add_79_2/U291  ( .A1(\sha1_round/add_79_2/n229 ), .A2(
        \sha1_round/add_79_2/n230 ), .ZN(\sha1_round/add_79_2/n225 ) );
  INV_X4 \sha1_round/add_79_2/U290  ( .A(w[19]), .ZN(
        \sha1_round/add_79_2/n227 ) );
  INV_X4 \sha1_round/add_79_2/U289  ( .A(rnd_q[19]), .ZN(
        \sha1_round/add_79_2/n228 ) );
  NAND2_X2 \sha1_round/add_79_2/U288  ( .A1(\sha1_round/add_79_2/n227 ), .A2(
        \sha1_round/add_79_2/n228 ), .ZN(\sha1_round/add_79_2/n186 ) );
  NAND2_X2 \sha1_round/add_79_2/U287  ( .A1(w[19]), .A2(rnd_q[19]), .ZN(
        \sha1_round/add_79_2/n220 ) );
  NAND2_X2 \sha1_round/add_79_2/U286  ( .A1(\sha1_round/add_79_2/n186 ), .A2(
        \sha1_round/add_79_2/n220 ), .ZN(\sha1_round/add_79_2/n226 ) );
  XNOR2_X2 \sha1_round/add_79_2/U285  ( .A(\sha1_round/add_79_2/n225 ), .B(
        \sha1_round/add_79_2/n226 ), .ZN(\sha1_round/N303 ) );
  XNOR2_X2 \sha1_round/add_79_2/U284  ( .A(\sha1_round/add_79_2/n223 ), .B(
        \sha1_round/add_79_2/n221 ), .ZN(\sha1_round/N285 ) );
  INV_X4 \sha1_round/add_79_2/U283  ( .A(\sha1_round/add_79_2/n220 ), .ZN(
        \sha1_round/add_79_2/n119 ) );
  NAND2_X2 \sha1_round/add_79_2/U282  ( .A1(\sha1_round/add_79_2/n217 ), .A2(
        \sha1_round/add_79_2/n218 ), .ZN(\sha1_round/add_79_2/n205 ) );
  INV_X4 \sha1_round/add_79_2/U281  ( .A(\sha1_round/add_79_2/n205 ), .ZN(
        \sha1_round/add_79_2/n197 ) );
  XNOR2_X2 \sha1_round/add_79_2/U280  ( .A(\sha1_round/add_79_2/n197 ), .B(
        \sha1_round/add_79_2/n216 ), .ZN(\sha1_round/N304 ) );
  NAND2_X2 \sha1_round/add_79_2/U279  ( .A1(w[21]), .A2(rnd_q[21]), .ZN(
        \sha1_round/add_79_2/n209 ) );
  INV_X4 \sha1_round/add_79_2/U278  ( .A(\sha1_round/add_79_2/n209 ), .ZN(
        \sha1_round/add_79_2/n212 ) );
  XNOR2_X2 \sha1_round/add_79_2/U277  ( .A(\sha1_round/add_79_2/n210 ), .B(
        \sha1_round/add_79_2/n211 ), .ZN(\sha1_round/N305 ) );
  NAND2_X2 \sha1_round/add_79_2/U276  ( .A1(\sha1_round/add_79_2/n208 ), .A2(
        \sha1_round/add_79_2/n209 ), .ZN(\sha1_round/add_79_2/n195 ) );
  INV_X4 \sha1_round/add_79_2/U275  ( .A(\sha1_round/add_79_2/n195 ), .ZN(
        \sha1_round/add_79_2/n203 ) );
  NAND2_X2 \sha1_round/add_79_2/U274  ( .A1(\sha1_round/add_79_2/n198 ), .A2(
        \sha1_round/add_79_2/n205 ), .ZN(\sha1_round/add_79_2/n204 ) );
  NAND2_X2 \sha1_round/add_79_2/U273  ( .A1(\sha1_round/add_79_2/n203 ), .A2(
        \sha1_round/add_79_2/n204 ), .ZN(\sha1_round/add_79_2/n199 ) );
  NAND2_X2 \sha1_round/add_79_2/U272  ( .A1(w[22]), .A2(rnd_q[22]), .ZN(
        \sha1_round/add_79_2/n194 ) );
  INV_X4 \sha1_round/add_79_2/U271  ( .A(w[22]), .ZN(
        \sha1_round/add_79_2/n201 ) );
  INV_X4 \sha1_round/add_79_2/U270  ( .A(rnd_q[22]), .ZN(
        \sha1_round/add_79_2/n202 ) );
  NAND2_X2 \sha1_round/add_79_2/U269  ( .A1(\sha1_round/add_79_2/n201 ), .A2(
        \sha1_round/add_79_2/n202 ), .ZN(\sha1_round/add_79_2/n196 ) );
  NAND2_X2 \sha1_round/add_79_2/U268  ( .A1(\sha1_round/add_79_2/n194 ), .A2(
        \sha1_round/add_79_2/n196 ), .ZN(\sha1_round/add_79_2/n200 ) );
  XNOR2_X2 \sha1_round/add_79_2/U267  ( .A(\sha1_round/add_79_2/n199 ), .B(
        \sha1_round/add_79_2/n200 ), .ZN(\sha1_round/N306 ) );
  NAND2_X2 \sha1_round/add_79_2/U266  ( .A1(\sha1_round/add_79_2/n198 ), .A2(
        \sha1_round/add_79_2/n196 ), .ZN(\sha1_round/add_79_2/n188 ) );
  NAND2_X2 \sha1_round/add_79_2/U265  ( .A1(\sha1_round/add_79_2/n195 ), .A2(
        \sha1_round/add_79_2/n196 ), .ZN(\sha1_round/add_79_2/n193 ) );
  NAND2_X2 \sha1_round/add_79_2/U264  ( .A1(\sha1_round/add_79_2/n193 ), .A2(
        \sha1_round/add_79_2/n194 ), .ZN(\sha1_round/add_79_2/n183 ) );
  INV_X4 \sha1_round/add_79_2/U263  ( .A(w[23]), .ZN(
        \sha1_round/add_79_2/n190 ) );
  INV_X4 \sha1_round/add_79_2/U262  ( .A(rnd_q[23]), .ZN(
        \sha1_round/add_79_2/n191 ) );
  NAND2_X2 \sha1_round/add_79_2/U261  ( .A1(\sha1_round/add_79_2/n190 ), .A2(
        \sha1_round/add_79_2/n191 ), .ZN(\sha1_round/add_79_2/n184 ) );
  NAND2_X2 \sha1_round/add_79_2/U260  ( .A1(w[23]), .A2(rnd_q[23]), .ZN(
        \sha1_round/add_79_2/n129 ) );
  NAND2_X2 \sha1_round/add_79_2/U259  ( .A1(\sha1_round/add_79_2/n184 ), .A2(
        \sha1_round/add_79_2/n129 ), .ZN(\sha1_round/add_79_2/n189 ) );
  INV_X4 \sha1_round/add_79_2/U258  ( .A(\sha1_round/add_79_2/n188 ), .ZN(
        \sha1_round/add_79_2/n187 ) );
  NAND2_X2 \sha1_round/add_79_2/U257  ( .A1(\sha1_round/add_79_2/n119 ), .A2(
        \sha1_round/add_79_2/n2 ), .ZN(\sha1_round/add_79_2/n170 ) );
  NAND2_X2 \sha1_round/add_79_2/U256  ( .A1(\sha1_round/add_79_2/n169 ), .A2(
        \sha1_round/add_79_2/n170 ), .ZN(\sha1_round/add_79_2/n181 ) );
  NAND2_X2 \sha1_round/add_79_2/U255  ( .A1(\sha1_round/add_79_2/n183 ), .A2(
        \sha1_round/add_79_2/n184 ), .ZN(\sha1_round/add_79_2/n122 ) );
  NAND2_X2 \sha1_round/add_79_2/U254  ( .A1(\sha1_round/add_79_2/n122 ), .A2(
        \sha1_round/add_79_2/n129 ), .ZN(\sha1_round/add_79_2/n182 ) );
  NOR2_X2 \sha1_round/add_79_2/U253  ( .A1(\sha1_round/add_79_2/n181 ), .A2(
        \sha1_round/add_79_2/n182 ), .ZN(\sha1_round/add_79_2/n180 ) );
  NAND2_X2 \sha1_round/add_79_2/U252  ( .A1(w[24]), .A2(rnd_q[24]), .ZN(
        \sha1_round/add_79_2/n175 ) );
  INV_X4 \sha1_round/add_79_2/U251  ( .A(\sha1_round/add_79_2/n175 ), .ZN(
        \sha1_round/add_79_2/n166 ) );
  NAND2_X2 \sha1_round/add_79_2/U250  ( .A1(\sha1_round/add_79_2/n169 ), .A2(
        \sha1_round/add_79_2/n170 ), .ZN(\sha1_round/add_79_2/n177 ) );
  NAND2_X2 \sha1_round/add_79_2/U249  ( .A1(\sha1_round/add_79_2/n122 ), .A2(
        \sha1_round/add_79_2/n129 ), .ZN(\sha1_round/add_79_2/n178 ) );
  NOR2_X2 \sha1_round/add_79_2/U248  ( .A1(\sha1_round/add_79_2/n177 ), .A2(
        \sha1_round/add_79_2/n178 ), .ZN(\sha1_round/add_79_2/n176 ) );
  NAND2_X2 \sha1_round/add_79_2/U247  ( .A1(\sha1_round/add_79_2/n174 ), .A2(
        \sha1_round/add_79_2/n175 ), .ZN(\sha1_round/add_79_2/n172 ) );
  INV_X4 \sha1_round/add_79_2/U246  ( .A(\sha1_round/add_79_2/n171 ), .ZN(
        \sha1_round/add_79_2/n167 ) );
  NAND4_X2 \sha1_round/add_79_2/U245  ( .A1(\sha1_round/add_79_2/n122 ), .A2(
        \sha1_round/add_79_2/n129 ), .A3(\sha1_round/add_79_2/n169 ), .A4(
        \sha1_round/add_79_2/n170 ), .ZN(\sha1_round/add_79_2/n168 ) );
  NAND2_X2 \sha1_round/add_79_2/U244  ( .A1(w[26]), .A2(rnd_q[26]), .ZN(
        \sha1_round/add_79_2/n140 ) );
  INV_X4 \sha1_round/add_79_2/U243  ( .A(w[26]), .ZN(
        \sha1_round/add_79_2/n160 ) );
  INV_X4 \sha1_round/add_79_2/U242  ( .A(rnd_q[26]), .ZN(
        \sha1_round/add_79_2/n161 ) );
  NAND2_X2 \sha1_round/add_79_2/U241  ( .A1(\sha1_round/add_79_2/n160 ), .A2(
        \sha1_round/add_79_2/n161 ), .ZN(\sha1_round/add_79_2/n158 ) );
  NAND2_X2 \sha1_round/add_79_2/U240  ( .A1(\sha1_round/add_79_2/n140 ), .A2(
        \sha1_round/add_79_2/n158 ), .ZN(\sha1_round/add_79_2/n159 ) );
  INV_X4 \sha1_round/add_79_2/U239  ( .A(\sha1_round/add_79_2/n140 ), .ZN(
        \sha1_round/add_79_2/n151 ) );
  INV_X4 \sha1_round/add_79_2/U238  ( .A(\sha1_round/add_79_2/n158 ), .ZN(
        \sha1_round/add_79_2/n149 ) );
  NAND2_X2 \sha1_round/add_79_2/U237  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(
        \sha1_round/add_79_2/n155 ) );
  NAND2_X2 \sha1_round/add_79_2/U236  ( .A1(w[24]), .A2(rnd_q[24]), .ZN(
        \sha1_round/add_79_2/n156 ) );
  NAND2_X2 \sha1_round/add_79_2/U235  ( .A1(\sha1_round/add_79_2/n155 ), .A2(
        \sha1_round/add_79_2/n156 ), .ZN(\sha1_round/add_79_2/n154 ) );
  NAND2_X2 \sha1_round/add_79_2/U234  ( .A1(\sha1_round/add_79_2/n153 ), .A2(
        \sha1_round/add_79_2/n154 ), .ZN(\sha1_round/add_79_2/n139 ) );
  INV_X4 \sha1_round/add_79_2/U233  ( .A(\sha1_round/add_79_2/n139 ), .ZN(
        \sha1_round/add_79_2/n152 ) );
  NAND2_X2 \sha1_round/add_79_2/U232  ( .A1(\sha1_round/add_79_2/n141 ), .A2(
        \sha1_round/add_79_2/n131 ), .ZN(\sha1_round/add_79_2/n147 ) );
  NAND2_X2 \sha1_round/add_79_2/U231  ( .A1(\sha1_round/add_79_2/n146 ), .A2(
        \sha1_round/add_79_2/n147 ), .ZN(\sha1_round/add_79_2/n142 ) );
  INV_X4 \sha1_round/add_79_2/U230  ( .A(w[27]), .ZN(
        \sha1_round/add_79_2/n144 ) );
  INV_X4 \sha1_round/add_79_2/U229  ( .A(rnd_q[27]), .ZN(
        \sha1_round/add_79_2/n145 ) );
  NAND2_X2 \sha1_round/add_79_2/U228  ( .A1(\sha1_round/add_79_2/n144 ), .A2(
        \sha1_round/add_79_2/n145 ), .ZN(\sha1_round/add_79_2/n130 ) );
  NAND2_X2 \sha1_round/add_79_2/U227  ( .A1(w[27]), .A2(rnd_q[27]), .ZN(
        \sha1_round/add_79_2/n137 ) );
  NAND2_X2 \sha1_round/add_79_2/U226  ( .A1(\sha1_round/add_79_2/n130 ), .A2(
        \sha1_round/add_79_2/n137 ), .ZN(\sha1_round/add_79_2/n143 ) );
  XNOR2_X2 \sha1_round/add_79_2/U225  ( .A(\sha1_round/add_79_2/n142 ), .B(
        \sha1_round/add_79_2/n143 ), .ZN(\sha1_round/N311 ) );
  NAND2_X2 \sha1_round/add_79_2/U224  ( .A1(\sha1_round/add_79_2/n139 ), .A2(
        \sha1_round/add_79_2/n140 ), .ZN(\sha1_round/add_79_2/n138 ) );
  NAND2_X2 \sha1_round/add_79_2/U223  ( .A1(\sha1_round/add_79_2/n138 ), .A2(
        \sha1_round/add_79_2/n130 ), .ZN(\sha1_round/add_79_2/n136 ) );
  NAND2_X2 \sha1_round/add_79_2/U222  ( .A1(\sha1_round/add_79_2/n136 ), .A2(
        \sha1_round/add_79_2/n137 ), .ZN(\sha1_round/add_79_2/n125 ) );
  INV_X4 \sha1_round/add_79_2/U221  ( .A(w[28]), .ZN(
        \sha1_round/add_79_2/n134 ) );
  INV_X4 \sha1_round/add_79_2/U220  ( .A(rnd_q[28]), .ZN(
        \sha1_round/add_79_2/n135 ) );
  NAND2_X2 \sha1_round/add_79_2/U219  ( .A1(\sha1_round/add_79_2/n134 ), .A2(
        \sha1_round/add_79_2/n135 ), .ZN(\sha1_round/add_79_2/n126 ) );
  NAND2_X2 \sha1_round/add_79_2/U218  ( .A1(w[28]), .A2(rnd_q[28]), .ZN(
        \sha1_round/add_79_2/n132 ) );
  NAND2_X2 \sha1_round/add_79_2/U217  ( .A1(\sha1_round/add_79_2/n126 ), .A2(
        \sha1_round/add_79_2/n132 ), .ZN(\sha1_round/add_79_2/n133 ) );
  INV_X4 \sha1_round/add_79_2/U216  ( .A(\sha1_round/add_79_2/n132 ), .ZN(
        \sha1_round/add_79_2/n127 ) );
  NAND2_X2 \sha1_round/add_79_2/U215  ( .A1(\sha1_round/add_79_2/n125 ), .A2(
        \sha1_round/add_79_2/n126 ), .ZN(\sha1_round/add_79_2/n124 ) );
  NAND2_X2 \sha1_round/add_79_2/U214  ( .A1(\sha1_round/add_79_2/n123 ), .A2(
        \sha1_round/add_79_2/n124 ), .ZN(\sha1_round/add_79_2/n97 ) );
  INV_X4 \sha1_round/add_79_2/U213  ( .A(\sha1_round/add_79_2/n122 ), .ZN(
        \sha1_round/add_79_2/n120 ) );
  INV_X4 \sha1_round/add_79_2/U212  ( .A(\sha1_round/add_79_2/n121 ), .ZN(
        \sha1_round/add_79_2/n115 ) );
  NAND2_X2 \sha1_round/add_79_2/U211  ( .A1(\sha1_round/add_79_2/n116 ), .A2(
        \sha1_round/add_79_2/n117 ), .ZN(\sha1_round/add_79_2/n94 ) );
  NAND2_X2 \sha1_round/add_79_2/U210  ( .A1(\sha1_round/add_79_2/n94 ), .A2(
        \sha1_round/add_79_2/n3 ), .ZN(\sha1_round/add_79_2/n114 ) );
  NAND2_X2 \sha1_round/add_79_2/U209  ( .A1(\sha1_round/add_79_2/n113 ), .A2(
        \sha1_round/add_79_2/n114 ), .ZN(\sha1_round/add_79_2/n109 ) );
  NAND2_X2 \sha1_round/add_79_2/U208  ( .A1(w[29]), .A2(rnd_q[29]), .ZN(
        \sha1_round/add_79_2/n96 ) );
  INV_X4 \sha1_round/add_79_2/U207  ( .A(w[29]), .ZN(
        \sha1_round/add_79_2/n111 ) );
  INV_X4 \sha1_round/add_79_2/U206  ( .A(rnd_q[29]), .ZN(
        \sha1_round/add_79_2/n112 ) );
  NAND2_X2 \sha1_round/add_79_2/U205  ( .A1(\sha1_round/add_79_2/n111 ), .A2(
        \sha1_round/add_79_2/n112 ), .ZN(\sha1_round/add_79_2/n99 ) );
  NAND2_X2 \sha1_round/add_79_2/U204  ( .A1(\sha1_round/add_79_2/n96 ), .A2(
        \sha1_round/add_79_2/n99 ), .ZN(\sha1_round/add_79_2/n110 ) );
  XNOR2_X2 \sha1_round/add_79_2/U203  ( .A(\sha1_round/add_79_2/n109 ), .B(
        \sha1_round/add_79_2/n110 ), .ZN(\sha1_round/N313 ) );
  XNOR2_X2 \sha1_round/add_79_2/U202  ( .A(\sha1_round/add_79_2/n86 ), .B(
        \sha1_round/add_79_2/n106 ), .ZN(\sha1_round/N286 ) );
  NAND2_X2 \sha1_round/add_79_2/U201  ( .A1(\sha1_round/add_79_2/n97 ), .A2(
        \sha1_round/add_79_2/n99 ), .ZN(\sha1_round/add_79_2/n103 ) );
  NAND2_X2 \sha1_round/add_79_2/U200  ( .A1(\sha1_round/add_79_2/n1 ), .A2(
        \sha1_round/add_79_2/n99 ), .ZN(\sha1_round/add_79_2/n104 ) );
  NAND4_X2 \sha1_round/add_79_2/U199  ( .A1(\sha1_round/add_79_2/n103 ), .A2(
        \sha1_round/add_79_2/n96 ), .A3(\sha1_round/add_79_2/n104 ), .A4(
        \sha1_round/add_79_2/n105 ), .ZN(\sha1_round/add_79_2/n100 ) );
  INV_X4 \sha1_round/add_79_2/U198  ( .A(w[30]), .ZN(
        \sha1_round/add_79_2/n101 ) );
  INV_X4 \sha1_round/add_79_2/U197  ( .A(rnd_q[30]), .ZN(
        \sha1_round/add_79_2/n102 ) );
  INV_X4 \sha1_round/add_79_2/U196  ( .A(\sha1_round/add_79_2/n99 ), .ZN(
        \sha1_round/add_79_2/n98 ) );
  NAND2_X2 \sha1_round/add_79_2/U195  ( .A1(\sha1_round/add_79_2/n93 ), .A2(
        \sha1_round/add_79_2/n97 ), .ZN(\sha1_round/add_79_2/n89 ) );
  NAND2_X2 \sha1_round/add_79_2/U194  ( .A1(\sha1_round/add_79_2/n93 ), .A2(
        \sha1_round/add_79_2/n1 ), .ZN(\sha1_round/add_79_2/n91 ) );
  NAND4_X2 \sha1_round/add_79_2/U193  ( .A1(\sha1_round/add_79_2/n89 ), .A2(
        \sha1_round/add_79_2/n90 ), .A3(\sha1_round/add_79_2/n91 ), .A4(
        \sha1_round/add_79_2/n92 ), .ZN(\sha1_round/add_79_2/n87 ) );
  XNOR2_X2 \sha1_round/add_79_2/U192  ( .A(w[31]), .B(rnd_q[31]), .ZN(
        \sha1_round/add_79_2/n88 ) );
  XNOR2_X2 \sha1_round/add_79_2/U191  ( .A(\sha1_round/add_79_2/n87 ), .B(
        \sha1_round/add_79_2/n88 ), .ZN(\sha1_round/N315 ) );
  NAND2_X2 \sha1_round/add_79_2/U190  ( .A1(\sha1_round/add_79_2/n72 ), .A2(
        \sha1_round/add_79_2/n83 ), .ZN(\sha1_round/add_79_2/n82 ) );
  INV_X4 \sha1_round/add_79_2/U189  ( .A(\sha1_round/add_79_2/n71 ), .ZN(
        \sha1_round/add_79_2/n64 ) );
  INV_X4 \sha1_round/add_79_2/U188  ( .A(\sha1_round/add_79_2/n81 ), .ZN(
        \sha1_round/add_79_2/n75 ) );
  XNOR2_X2 \sha1_round/add_79_2/U187  ( .A(\sha1_round/add_79_2/n48 ), .B(
        \sha1_round/add_79_2/n80 ), .ZN(\sha1_round/N288 ) );
  INV_X4 \sha1_round/add_79_2/U186  ( .A(\sha1_round/add_79_2/n69 ), .ZN(
        \sha1_round/add_79_2/n62 ) );
  XNOR2_X2 \sha1_round/add_79_2/U185  ( .A(\sha1_round/add_79_2/n77 ), .B(
        \sha1_round/add_79_2/n78 ), .ZN(\sha1_round/N289 ) );
  INV_X4 \sha1_round/add_79_2/U184  ( .A(\sha1_round/add_79_2/n60 ), .ZN(
        \sha1_round/add_79_2/n70 ) );
  NAND2_X2 \sha1_round/add_79_2/U183  ( .A1(\sha1_round/add_79_2/n68 ), .A2(
        \sha1_round/add_79_2/n69 ), .ZN(\sha1_round/add_79_2/n67 ) );
  INV_X4 \sha1_round/add_79_2/U182  ( .A(\sha1_round/add_79_2/n66 ), .ZN(
        \sha1_round/add_79_2/n65 ) );
  XNOR2_X2 \sha1_round/add_79_2/U181  ( .A(\sha1_round/add_79_2/n54 ), .B(
        \sha1_round/add_79_2/n55 ), .ZN(\sha1_round/N291 ) );
  INV_X4 \sha1_round/add_79_2/U180  ( .A(\sha1_round/add_79_2/n52 ), .ZN(
        \sha1_round/add_79_2/n43 ) );
  XNOR2_X2 \sha1_round/add_79_2/U179  ( .A(\sha1_round/add_79_2/n50 ), .B(
        \sha1_round/add_79_2/n51 ), .ZN(\sha1_round/N292 ) );
  XNOR2_X2 \sha1_round/add_79_2/U178  ( .A(\sha1_round/add_79_2/n38 ), .B(
        \sha1_round/add_79_2/n39 ), .ZN(\sha1_round/N293 ) );
  NAND2_X2 \sha1_round/add_79_2/U177  ( .A1(\sha1_round/add_79_2/n72 ), .A2(
        \sha1_round/add_79_2/n73 ), .ZN(\sha1_round/add_79_2/n368 ) );
  AND2_X2 \sha1_round/add_79_2/U176  ( .A1(w[11]), .A2(rnd_q[11]), .ZN(
        \sha1_round/add_79_2/n37 ) );
  AND2_X2 \sha1_round/add_79_2/U175  ( .A1(w[2]), .A2(rnd_q[2]), .ZN(
        \sha1_round/add_79_2/n36 ) );
  AND2_X2 \sha1_round/add_79_2/U174  ( .A1(w[6]), .A2(rnd_q[6]), .ZN(
        \sha1_round/add_79_2/n35 ) );
  NOR2_X2 \sha1_round/add_79_2/U173  ( .A1(rnd_q[20]), .A2(w[20]), .ZN(
        \sha1_round/add_79_2/n207 ) );
  NOR2_X2 \sha1_round/add_79_2/U172  ( .A1(rnd_q[21]), .A2(w[21]), .ZN(
        \sha1_round/add_79_2/n206 ) );
  NOR2_X2 \sha1_round/add_79_2/U171  ( .A1(\sha1_round/add_79_2/n206 ), .A2(
        \sha1_round/add_79_2/n207 ), .ZN(\sha1_round/add_79_2/n198 ) );
  NOR2_X2 \sha1_round/add_79_2/U170  ( .A1(rnd_q[10]), .A2(w[10]), .ZN(
        \sha1_round/add_79_2/n341 ) );
  AND2_X2 \sha1_round/add_79_2/U169  ( .A1(w[10]), .A2(rnd_q[10]), .ZN(
        \sha1_round/add_79_2/n34 ) );
  OR2_X2 \sha1_round/add_79_2/U168  ( .A1(w[3]), .A2(rnd_q[3]), .ZN(
        \sha1_round/add_79_2/n83 ) );
  NOR2_X2 \sha1_round/add_79_2/U167  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(
        \sha1_round/add_79_2/n157 ) );
  NOR2_X2 \sha1_round/add_79_2/U166  ( .A1(\sha1_round/add_79_2/n149 ), .A2(
        \sha1_round/add_79_2/n157 ), .ZN(\sha1_round/add_79_2/n153 ) );
  NAND3_X2 \sha1_round/add_79_2/U165  ( .A1(rnd_q[20]), .A2(
        \sha1_round/add_79_2/n11 ), .A3(w[20]), .ZN(\sha1_round/add_79_2/n208 ) );
  NAND3_X2 \sha1_round/add_79_2/U164  ( .A1(rnd_q[16]), .A2(w[16]), .A3(
        \sha1_round/add_79_2/n244 ), .ZN(\sha1_round/add_79_2/n242 ) );
  NOR2_X2 \sha1_round/add_79_2/U163  ( .A1(rnd_q[20]), .A2(w[20]), .ZN(
        \sha1_round/add_79_2/n215 ) );
  NOR2_X2 \sha1_round/add_79_2/U162  ( .A1(rnd_q[5]), .A2(w[5]), .ZN(
        \sha1_round/add_79_2/n365 ) );
  NOR2_X2 \sha1_round/add_79_2/U161  ( .A1(\sha1_round/add_79_2/n56 ), .A2(
        \sha1_round/add_79_2/n365 ), .ZN(\sha1_round/add_79_2/n364 ) );
  NOR2_X2 \sha1_round/add_79_2/U160  ( .A1(\sha1_round/add_79_2/n9 ), .A2(
        \sha1_round/add_79_2/n95 ), .ZN(\sha1_round/add_79_2/n90 ) );
  NOR2_X2 \sha1_round/add_79_2/U159  ( .A1(\sha1_round/add_79_2/n298 ), .A2(
        \sha1_round/add_79_2/n374 ), .ZN(\sha1_round/add_79_2/n76 ) );
  NOR2_X2 \sha1_round/add_79_2/U158  ( .A1(rnd_q[0]), .A2(w[0]), .ZN(
        \sha1_round/add_79_2/n224 ) );
  NOR2_X2 \sha1_round/add_79_2/U157  ( .A1(\sha1_round/add_79_2/n299 ), .A2(
        \sha1_round/add_79_2/n224 ), .ZN(\sha1_round/N284 ) );
  NOR2_X2 \sha1_round/add_79_2/U156  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(
        \sha1_round/add_79_2/n164 ) );
  NAND3_X2 \sha1_round/add_79_2/U155  ( .A1(rnd_q[9]), .A2(w[9]), .A3(
        \sha1_round/add_79_2/n337 ), .ZN(\sha1_round/add_79_2/n333 ) );
  NOR2_X2 \sha1_round/add_79_2/U154  ( .A1(\sha1_round/add_79_2/n34 ), .A2(
        \sha1_round/add_79_2/n37 ), .ZN(\sha1_round/add_79_2/n334 ) );
  NAND3_X2 \sha1_round/add_79_2/U153  ( .A1(\sha1_round/add_79_2/n332 ), .A2(
        \sha1_round/add_79_2/n333 ), .A3(\sha1_round/add_79_2/n334 ), .ZN(
        \sha1_round/add_79_2/n286 ) );
  NOR2_X2 \sha1_round/add_79_2/U152  ( .A1(rnd_q[10]), .A2(w[10]), .ZN(
        \sha1_round/add_79_2/n335 ) );
  NOR2_X2 \sha1_round/add_79_2/U151  ( .A1(rnd_q[21]), .A2(w[21]), .ZN(
        \sha1_round/add_79_2/n213 ) );
  NOR2_X2 \sha1_round/add_79_2/U150  ( .A1(\sha1_round/add_79_2/n214 ), .A2(
        \sha1_round/add_79_2/n7 ), .ZN(\sha1_round/add_79_2/n210 ) );
  NOR2_X2 \sha1_round/add_79_2/U149  ( .A1(\sha1_round/add_79_2/n212 ), .A2(
        \sha1_round/add_79_2/n213 ), .ZN(\sha1_round/add_79_2/n211 ) );
  NOR2_X2 \sha1_round/add_79_2/U148  ( .A1(rnd_q[9]), .A2(w[9]), .ZN(
        \sha1_round/add_79_2/n41 ) );
  NOR2_X2 \sha1_round/add_79_2/U147  ( .A1(rnd_q[8]), .A2(w[8]), .ZN(
        \sha1_round/add_79_2/n44 ) );
  NOR2_X2 \sha1_round/add_79_2/U146  ( .A1(rnd_q[16]), .A2(w[16]), .ZN(
        \sha1_round/add_79_2/n231 ) );
  OR2_X2 \sha1_round/add_79_2/U145  ( .A1(w[11]), .A2(rnd_q[11]), .ZN(
        \sha1_round/add_79_2/n285 ) );
  NOR2_X2 \sha1_round/add_79_2/U144  ( .A1(rnd_q[24]), .A2(w[24]), .ZN(
        \sha1_round/add_79_2/n148 ) );
  NOR2_X2 \sha1_round/add_79_2/U143  ( .A1(rnd_q[1]), .A2(w[1]), .ZN(
        \sha1_round/add_79_2/n107 ) );
  NOR2_X2 \sha1_round/add_79_2/U142  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(
        \sha1_round/add_79_2/n150 ) );
  NOR3_X2 \sha1_round/add_79_2/U141  ( .A1(\sha1_round/add_79_2/n148 ), .A2(
        \sha1_round/add_79_2/n149 ), .A3(\sha1_round/add_79_2/n150 ), .ZN(
        \sha1_round/add_79_2/n131 ) );
  NOR2_X2 \sha1_round/add_79_2/U140  ( .A1(rnd_q[2]), .A2(w[2]), .ZN(
        \sha1_round/add_79_2/n85 ) );
  NOR2_X2 \sha1_round/add_79_2/U139  ( .A1(rnd_q[6]), .A2(w[6]), .ZN(
        \sha1_round/add_79_2/n61 ) );
  NOR2_X2 \sha1_round/add_79_2/U138  ( .A1(rnd_q[5]), .A2(w[5]), .ZN(
        \sha1_round/add_79_2/n60 ) );
  OR2_X2 \sha1_round/add_79_2/U137  ( .A1(w[7]), .A2(rnd_q[7]), .ZN(
        \sha1_round/add_79_2/n262 ) );
  NOR2_X2 \sha1_round/add_79_2/U136  ( .A1(\sha1_round/add_79_2/n4 ), .A2(
        \sha1_round/add_79_2/n96 ), .ZN(\sha1_round/add_79_2/n95 ) );
  NOR2_X2 \sha1_round/add_79_2/U135  ( .A1(\sha1_round/add_79_2/n4 ), .A2(
        \sha1_round/add_79_2/n98 ), .ZN(\sha1_round/add_79_2/n93 ) );
  OR2_X2 \sha1_round/add_79_2/U134  ( .A1(\sha1_round/add_79_2/n60 ), .A2(
        \sha1_round/add_79_2/n61 ), .ZN(\sha1_round/add_79_2/n33 ) );
  AND3_X2 \sha1_round/add_79_2/U133  ( .A1(\sha1_round/add_79_2/n131 ), .A2(
        \sha1_round/add_79_2/n130 ), .A3(\sha1_round/add_79_2/n141 ), .ZN(
        \sha1_round/add_79_2/n32 ) );
  OR2_X2 \sha1_round/add_79_2/U132  ( .A1(\sha1_round/add_79_2/n44 ), .A2(
        \sha1_round/add_79_2/n41 ), .ZN(\sha1_round/add_79_2/n31 ) );
  AND2_X2 \sha1_round/add_79_2/U131  ( .A1(\sha1_round/add_79_2/n282 ), .A2(
        \sha1_round/add_79_2/n281 ), .ZN(\sha1_round/add_79_2/n277 ) );
  NOR2_X2 \sha1_round/add_79_2/U130  ( .A1(\sha1_round/add_79_2/n340 ), .A2(
        \sha1_round/add_79_2/n341 ), .ZN(\sha1_round/add_79_2/n339 ) );
  NAND3_X2 \sha1_round/add_79_2/U129  ( .A1(\sha1_round/add_79_2/n336 ), .A2(
        \sha1_round/add_79_2/n338 ), .A3(\sha1_round/add_79_2/n339 ), .ZN(
        \sha1_round/add_79_2/n264 ) );
  NAND3_X2 \sha1_round/add_79_2/U128  ( .A1(\sha1_round/add_79_2/n70 ), .A2(
        \sha1_round/add_79_2/n71 ), .A3(\sha1_round/add_79_2/n66 ), .ZN(
        \sha1_round/add_79_2/n68 ) );
  NAND3_X2 \sha1_round/add_79_2/U127  ( .A1(\sha1_round/add_79_2/n3 ), .A2(
        \sha1_round/add_79_2/n99 ), .A3(\sha1_round/add_79_2/n94 ), .ZN(
        \sha1_round/add_79_2/n105 ) );
  NOR2_X2 \sha1_round/add_79_2/U126  ( .A1(\sha1_round/add_79_2/n222 ), .A2(
        \sha1_round/add_79_2/n107 ), .ZN(\sha1_round/add_79_2/n221 ) );
  NOR2_X2 \sha1_round/add_79_2/U125  ( .A1(\sha1_round/add_79_2/n61 ), .A2(
        \sha1_round/add_79_2/n60 ), .ZN(\sha1_round/add_79_2/n266 ) );
  NOR2_X2 \sha1_round/add_79_2/U124  ( .A1(\sha1_round/add_79_2/n48 ), .A2(
        \sha1_round/add_79_2/n49 ), .ZN(\sha1_round/add_79_2/n356 ) );
  NOR2_X2 \sha1_round/add_79_2/U123  ( .A1(\sha1_round/add_79_2/n356 ), .A2(
        \sha1_round/add_79_2/n357 ), .ZN(\sha1_round/add_79_2/n355 ) );
  NOR2_X2 \sha1_round/add_79_2/U122  ( .A1(\sha1_round/add_79_2/n48 ), .A2(
        \sha1_round/add_79_2/n49 ), .ZN(\sha1_round/add_79_2/n350 ) );
  NAND3_X2 \sha1_round/add_79_2/U121  ( .A1(\sha1_round/add_79_2/n52 ), .A2(
        \sha1_round/add_79_2/n349 ), .A3(\sha1_round/add_79_2/n321 ), .ZN(
        \sha1_round/add_79_2/n351 ) );
  NOR2_X2 \sha1_round/add_79_2/U120  ( .A1(\sha1_round/add_79_2/n350 ), .A2(
        \sha1_round/add_79_2/n351 ), .ZN(\sha1_round/add_79_2/n347 ) );
  NOR2_X2 \sha1_round/add_79_2/U119  ( .A1(\sha1_round/add_79_2/n48 ), .A2(
        \sha1_round/add_79_2/n49 ), .ZN(\sha1_round/add_79_2/n46 ) );
  NOR2_X2 \sha1_round/add_79_2/U118  ( .A1(\sha1_round/add_79_2/n46 ), .A2(
        \sha1_round/add_79_2/n47 ), .ZN(\sha1_round/add_79_2/n45 ) );
  NAND3_X2 \sha1_round/add_79_2/U117  ( .A1(\sha1_round/add_79_2/n73 ), .A2(
        \sha1_round/add_79_2/n72 ), .A3(\sha1_round/add_79_2/n275 ), .ZN(
        \sha1_round/add_79_2/n318 ) );
  NOR4_X2 \sha1_round/add_79_2/U116  ( .A1(\sha1_round/add_79_2/n297 ), .A2(
        \sha1_round/add_79_2/n298 ), .A3(\sha1_round/add_79_2/n85 ), .A4(
        \sha1_round/add_79_2/n107 ), .ZN(\sha1_round/add_79_2/n296 ) );
  NOR2_X2 \sha1_round/add_79_2/U115  ( .A1(\sha1_round/add_79_2/n294 ), .A2(
        \sha1_round/add_79_2/n295 ), .ZN(\sha1_round/add_79_2/n287 ) );
  NOR2_X2 \sha1_round/add_79_2/U114  ( .A1(\sha1_round/add_79_2/n121 ), .A2(
        \sha1_round/add_79_2/n129 ), .ZN(\sha1_round/add_79_2/n128 ) );
  NOR2_X2 \sha1_round/add_79_2/U113  ( .A1(\sha1_round/add_79_2/n151 ), .A2(
        \sha1_round/add_79_2/n152 ), .ZN(\sha1_round/add_79_2/n146 ) );
  NOR2_X2 \sha1_round/add_79_2/U112  ( .A1(\sha1_round/add_79_2/n166 ), .A2(
        \sha1_round/add_79_2/n6 ), .ZN(\sha1_round/add_79_2/n165 ) );
  NOR2_X2 \sha1_round/add_79_2/U111  ( .A1(\sha1_round/add_79_2/n164 ), .A2(
        \sha1_round/add_79_2/n165 ), .ZN(\sha1_round/add_79_2/n163 ) );
  NOR2_X2 \sha1_round/add_79_2/U110  ( .A1(\sha1_round/add_79_2/n85 ), .A2(
        \sha1_round/add_79_2/n86 ), .ZN(\sha1_round/add_79_2/n84 ) );
  NAND3_X2 \sha1_round/add_79_2/U109  ( .A1(\sha1_round/add_79_2/n185 ), .A2(
        \sha1_round/add_79_2/n186 ), .A3(\sha1_round/add_79_2/n2 ), .ZN(
        \sha1_round/add_79_2/n169 ) );
  NOR2_X2 \sha1_round/add_79_2/U108  ( .A1(\sha1_round/add_79_2/n75 ), .A2(
        \sha1_round/add_79_2/n76 ), .ZN(\sha1_round/add_79_2/n74 ) );
  NAND3_X2 \sha1_round/add_79_2/U107  ( .A1(\sha1_round/add_79_2/n73 ), .A2(
        \sha1_round/add_79_2/n74 ), .A3(\sha1_round/add_79_2/n72 ), .ZN(
        \sha1_round/add_79_2/n66 ) );
  NOR2_X2 \sha1_round/add_79_2/U106  ( .A1(\sha1_round/add_79_2/n298 ), .A2(
        \sha1_round/add_79_2/n85 ), .ZN(\sha1_round/add_79_2/n371 ) );
  NAND3_X2 \sha1_round/add_79_2/U105  ( .A1(\sha1_round/add_79_2/n369 ), .A2(
        \sha1_round/add_79_2/n370 ), .A3(\sha1_round/add_79_2/n371 ), .ZN(
        \sha1_round/add_79_2/n73 ) );
  NAND3_X2 \sha1_round/add_79_2/U104  ( .A1(\sha1_round/add_79_2/n358 ), .A2(
        \sha1_round/add_79_2/n269 ), .A3(\sha1_round/add_79_2/n359 ), .ZN(
        \sha1_round/add_79_2/n47 ) );
  AND2_X4 \sha1_round/add_79_2/U103  ( .A1(\sha1_round/add_79_2/n31 ), .A2(
        \sha1_round/add_79_2/n349 ), .ZN(\sha1_round/add_79_2/n29 ) );
  OR2_X2 \sha1_round/add_79_2/U102  ( .A1(\sha1_round/add_79_2/n29 ), .A2(
        \sha1_round/add_79_2/n335 ), .ZN(\sha1_round/add_79_2/n348 ) );
  NAND3_X2 \sha1_round/add_79_2/U101  ( .A1(\sha1_round/add_79_2/n130 ), .A2(
        \sha1_round/add_79_2/n126 ), .A3(\sha1_round/add_79_2/n131 ), .ZN(
        \sha1_round/add_79_2/n121 ) );
  NOR3_X2 \sha1_round/add_79_2/U100  ( .A1(\sha1_round/add_79_2/n245 ), .A2(
        \sha1_round/add_79_2/n233 ), .A3(\sha1_round/add_79_2/n231 ), .ZN(
        \sha1_round/add_79_2/n241 ) );
  NOR2_X2 \sha1_round/add_79_2/U99  ( .A1(\sha1_round/add_79_2/n60 ), .A2(
        \sha1_round/add_79_2/n61 ), .ZN(\sha1_round/add_79_2/n361 ) );
  OR2_X4 \sha1_round/add_79_2/U98  ( .A1(\sha1_round/add_79_2/n107 ), .A2(
        \sha1_round/add_79_2/n223 ), .ZN(\sha1_round/add_79_2/n28 ) );
  AND2_X2 \sha1_round/add_79_2/U97  ( .A1(\sha1_round/add_79_2/n108 ), .A2(
        \sha1_round/add_79_2/n28 ), .ZN(\sha1_round/add_79_2/n86 ) );
  NOR3_X2 \sha1_round/add_79_2/U96  ( .A1(\sha1_round/add_79_2/n231 ), .A2(
        \sha1_round/add_79_2/n232 ), .A3(\sha1_round/add_79_2/n233 ), .ZN(
        \sha1_round/add_79_2/n219 ) );
  OR2_X4 \sha1_round/add_79_2/U95  ( .A1(\sha1_round/add_79_2/n4 ), .A2(
        \sha1_round/add_79_2/n9 ), .ZN(\sha1_round/add_79_2/n27 ) );
  XNOR2_X2 \sha1_round/add_79_2/U94  ( .A(\sha1_round/add_79_2/n100 ), .B(
        \sha1_round/add_79_2/n27 ), .ZN(\sha1_round/N314 ) );
  NOR2_X2 \sha1_round/add_79_2/U93  ( .A1(\sha1_round/add_79_2/n319 ), .A2(
        \sha1_round/add_79_2/n320 ), .ZN(\sha1_round/add_79_2/n315 ) );
  NOR2_X2 \sha1_round/add_79_2/U92  ( .A1(\sha1_round/add_79_2/n127 ), .A2(
        \sha1_round/add_79_2/n128 ), .ZN(\sha1_round/add_79_2/n123 ) );
  NOR2_X2 \sha1_round/add_79_2/U91  ( .A1(\sha1_round/add_79_2/n164 ), .A2(
        \sha1_round/add_79_2/n6 ), .ZN(\sha1_round/add_79_2/n173 ) );
  XOR2_X2 \sha1_round/add_79_2/U90  ( .A(\sha1_round/add_79_2/n172 ), .B(
        \sha1_round/add_79_2/n173 ), .Z(\sha1_round/N309 ) );
  NOR2_X2 \sha1_round/add_79_2/U89  ( .A1(\sha1_round/add_79_2/n355 ), .A2(
        \sha1_round/add_79_2/n31 ), .ZN(\sha1_round/add_79_2/n354 ) );
  NOR2_X2 \sha1_round/add_79_2/U88  ( .A1(\sha1_round/add_79_2/n40 ), .A2(
        \sha1_round/add_79_2/n354 ), .ZN(\sha1_round/add_79_2/n352 ) );
  NOR2_X2 \sha1_round/add_79_2/U87  ( .A1(\sha1_round/add_79_2/n34 ), .A2(
        \sha1_round/add_79_2/n335 ), .ZN(\sha1_round/add_79_2/n353 ) );
  NOR2_X2 \sha1_round/add_79_2/U86  ( .A1(\sha1_round/add_79_2/n97 ), .A2(
        \sha1_round/add_79_2/n1 ), .ZN(\sha1_round/add_79_2/n113 ) );
  NOR2_X2 \sha1_round/add_79_2/U85  ( .A1(\sha1_round/add_79_2/n233 ), .A2(
        \sha1_round/add_79_2/n248 ), .ZN(\sha1_round/add_79_2/n247 ) );
  XOR2_X2 \sha1_round/add_79_2/U84  ( .A(\sha1_round/add_79_2/n246 ), .B(
        \sha1_round/add_79_2/n247 ), .Z(\sha1_round/N301 ) );
  OR2_X4 \sha1_round/add_79_2/U83  ( .A1(\sha1_round/add_79_2/n32 ), .A2(
        \sha1_round/add_79_2/n125 ), .ZN(\sha1_round/add_79_2/n25 ) );
  XNOR2_X2 \sha1_round/add_79_2/U82  ( .A(\sha1_round/add_79_2/n25 ), .B(
        \sha1_round/add_79_2/n133 ), .ZN(\sha1_round/N312 ) );
  NOR2_X2 \sha1_round/add_79_2/U81  ( .A1(\sha1_round/add_79_2/n148 ), .A2(
        \sha1_round/add_79_2/n166 ), .ZN(\sha1_round/add_79_2/n179 ) );
  XOR2_X2 \sha1_round/add_79_2/U80  ( .A(\sha1_round/add_79_2/n141 ), .B(
        \sha1_round/add_79_2/n179 ), .Z(\sha1_round/N308 ) );
  NOR2_X2 \sha1_round/add_79_2/U79  ( .A1(\sha1_round/add_79_2/n48 ), .A2(
        \sha1_round/add_79_2/n49 ), .ZN(\sha1_round/add_79_2/n53 ) );
  NOR2_X2 \sha1_round/add_79_2/U78  ( .A1(\sha1_round/add_79_2/n53 ), .A2(
        \sha1_round/add_79_2/n47 ), .ZN(\sha1_round/add_79_2/n50 ) );
  NOR2_X2 \sha1_round/add_79_2/U77  ( .A1(\sha1_round/add_79_2/n44 ), .A2(
        \sha1_round/add_79_2/n43 ), .ZN(\sha1_round/add_79_2/n51 ) );
  NOR2_X2 \sha1_round/add_79_2/U76  ( .A1(\sha1_round/add_79_2/n44 ), .A2(
        \sha1_round/add_79_2/n45 ), .ZN(\sha1_round/add_79_2/n42 ) );
  NOR2_X2 \sha1_round/add_79_2/U75  ( .A1(\sha1_round/add_79_2/n42 ), .A2(
        \sha1_round/add_79_2/n43 ), .ZN(\sha1_round/add_79_2/n38 ) );
  NOR2_X2 \sha1_round/add_79_2/U74  ( .A1(\sha1_round/add_79_2/n40 ), .A2(
        \sha1_round/add_79_2/n41 ), .ZN(\sha1_round/add_79_2/n39 ) );
  NOR2_X2 \sha1_round/add_79_2/U73  ( .A1(\sha1_round/add_79_2/n347 ), .A2(
        \sha1_round/add_79_2/n348 ), .ZN(\sha1_round/add_79_2/n346 ) );
  NOR2_X2 \sha1_round/add_79_2/U72  ( .A1(\sha1_round/add_79_2/n346 ), .A2(
        \sha1_round/add_79_2/n34 ), .ZN(\sha1_round/add_79_2/n344 ) );
  NOR2_X2 \sha1_round/add_79_2/U71  ( .A1(\sha1_round/add_79_2/n7 ), .A2(
        \sha1_round/add_79_2/n215 ), .ZN(\sha1_round/add_79_2/n216 ) );
  NOR2_X2 \sha1_round/add_79_2/U70  ( .A1(\sha1_round/add_79_2/n59 ), .A2(
        \sha1_round/add_79_2/n33 ), .ZN(\sha1_round/add_79_2/n58 ) );
  NOR2_X2 \sha1_round/add_79_2/U69  ( .A1(\sha1_round/add_79_2/n58 ), .A2(
        \sha1_round/add_79_2/n35 ), .ZN(\sha1_round/add_79_2/n54 ) );
  AND3_X4 \sha1_round/add_79_2/U68  ( .A1(\sha1_round/add_79_2/n281 ), .A2(
        \sha1_round/add_79_2/n282 ), .A3(\sha1_round/add_79_2/n300 ), .ZN(
        \sha1_round/add_79_2/n24 ) );
  AND2_X2 \sha1_round/add_79_2/U67  ( .A1(\sha1_round/add_79_2/n301 ), .A2(
        \sha1_round/add_79_2/n24 ), .ZN(\sha1_round/add_79_2/n261 ) );
  NOR2_X2 \sha1_round/add_79_2/U66  ( .A1(\sha1_round/add_79_2/n76 ), .A2(
        \sha1_round/add_79_2/n368 ), .ZN(\sha1_round/add_79_2/n48 ) );
  NOR2_X2 \sha1_round/add_79_2/U65  ( .A1(\sha1_round/add_79_2/n48 ), .A2(
        \sha1_round/add_79_2/n64 ), .ZN(\sha1_round/add_79_2/n79 ) );
  NOR2_X2 \sha1_round/add_79_2/U64  ( .A1(\sha1_round/add_79_2/n79 ), .A2(
        \sha1_round/add_79_2/n75 ), .ZN(\sha1_round/add_79_2/n77 ) );
  NOR2_X2 \sha1_round/add_79_2/U63  ( .A1(\sha1_round/add_79_2/n62 ), .A2(
        \sha1_round/add_79_2/n60 ), .ZN(\sha1_round/add_79_2/n78 ) );
  NOR2_X2 \sha1_round/add_79_2/U62  ( .A1(\sha1_round/add_79_2/n36 ), .A2(
        \sha1_round/add_79_2/n85 ), .ZN(\sha1_round/add_79_2/n106 ) );
  NAND3_X2 \sha1_round/add_79_2/U61  ( .A1(\sha1_round/add_79_2/n93 ), .A2(
        \sha1_round/add_79_2/n3 ), .A3(\sha1_round/add_79_2/n94 ), .ZN(
        \sha1_round/add_79_2/n92 ) );
  NAND3_X2 \sha1_round/add_79_2/U60  ( .A1(\sha1_round/add_79_2/n330 ), .A2(
        \sha1_round/add_79_2/n322 ), .A3(\sha1_round/add_79_2/n10 ), .ZN(
        \sha1_round/add_79_2/n328 ) );
  NAND3_X2 \sha1_round/add_79_2/U59  ( .A1(\sha1_round/add_79_2/n5 ), .A2(
        \sha1_round/add_79_2/n2 ), .A3(\sha1_round/add_79_2/n118 ), .ZN(
        \sha1_round/add_79_2/n171 ) );
  NOR2_X2 \sha1_round/add_79_2/U58  ( .A1(\sha1_round/add_79_2/n64 ), .A2(
        \sha1_round/add_79_2/n65 ), .ZN(\sha1_round/add_79_2/n63 ) );
  NOR2_X2 \sha1_round/add_79_2/U57  ( .A1(\sha1_round/add_79_2/n62 ), .A2(
        \sha1_round/add_79_2/n63 ), .ZN(\sha1_round/add_79_2/n59 ) );
  NOR2_X2 \sha1_round/add_79_2/U56  ( .A1(\sha1_round/add_79_2/n197 ), .A2(
        \sha1_round/add_79_2/n188 ), .ZN(\sha1_round/add_79_2/n192 ) );
  NOR2_X2 \sha1_round/add_79_2/U55  ( .A1(\sha1_round/add_79_2/n222 ), .A2(
        \sha1_round/add_79_2/n299 ), .ZN(\sha1_round/add_79_2/n297 ) );
  NOR2_X2 \sha1_round/add_79_2/U54  ( .A1(\sha1_round/add_79_2/n119 ), .A2(
        \sha1_round/add_79_2/n8 ), .ZN(\sha1_round/add_79_2/n217 ) );
  NOR2_X2 \sha1_round/add_79_2/U53  ( .A1(\sha1_round/add_79_2/n287 ), .A2(
        \sha1_round/add_79_2/n288 ), .ZN(\sha1_round/add_79_2/n255 ) );
  NAND3_X2 \sha1_round/add_79_2/U52  ( .A1(\sha1_round/add_79_2/n255 ), .A2(
        \sha1_round/add_79_2/n12 ), .A3(\sha1_round/add_79_2/n256 ), .ZN(
        \sha1_round/add_79_2/n118 ) );
  NOR2_X2 \sha1_round/add_79_2/U51  ( .A1(\sha1_round/add_79_2/n119 ), .A2(
        \sha1_round/add_79_2/n8 ), .ZN(\sha1_round/add_79_2/n116 ) );
  NOR2_X2 \sha1_round/add_79_2/U50  ( .A1(\sha1_round/add_79_2/n64 ), .A2(
        \sha1_round/add_79_2/n75 ), .ZN(\sha1_round/add_79_2/n80 ) );
  NOR2_X1 \sha1_round/add_79_2/U49  ( .A1(\sha1_round/add_79_2/n56 ), .A2(
        \sha1_round/add_79_2/n362 ), .ZN(\sha1_round/add_79_2/n276 ) );
  OR2_X4 \sha1_round/add_79_2/U48  ( .A1(\sha1_round/add_79_2/n164 ), .A2(
        \sha1_round/add_79_2/n148 ), .ZN(\sha1_round/add_79_2/n23 ) );
  NOR2_X2 \sha1_round/add_79_2/U47  ( .A1(\sha1_round/add_79_2/n167 ), .A2(
        \sha1_round/add_79_2/n168 ), .ZN(\sha1_round/add_79_2/n22 ) );
  NOR2_X2 \sha1_round/add_79_2/U46  ( .A1(\sha1_round/add_79_2/n22 ), .A2(
        \sha1_round/add_79_2/n23 ), .ZN(\sha1_round/add_79_2/n162 ) );
  AND2_X2 \sha1_round/add_79_2/U45  ( .A1(\sha1_round/add_79_2/n171 ), .A2(
        \sha1_round/add_79_2/n176 ), .ZN(\sha1_round/add_79_2/n21 ) );
  OR2_X2 \sha1_round/add_79_2/U44  ( .A1(\sha1_round/add_79_2/n21 ), .A2(
        \sha1_round/add_79_2/n148 ), .ZN(\sha1_round/add_79_2/n174 ) );
  NAND2_X2 \sha1_round/add_79_2/U43  ( .A1(\sha1_round/add_79_2/n300 ), .A2(
        \sha1_round/add_79_2/n281 ), .ZN(\sha1_round/add_79_2/n20 ) );
  AND3_X4 \sha1_round/add_79_2/U42  ( .A1(\sha1_round/add_79_2/n292 ), .A2(
        \sha1_round/add_79_2/n279 ), .A3(\sha1_round/add_79_2/n307 ), .ZN(
        \sha1_round/add_79_2/n19 ) );
  NOR2_X2 \sha1_round/add_79_2/U41  ( .A1(\sha1_round/add_79_2/n19 ), .A2(
        \sha1_round/add_79_2/n20 ), .ZN(\sha1_round/add_79_2/n305 ) );
  NAND3_X1 \sha1_round/add_79_2/U40  ( .A1(\sha1_round/add_79_2/n261 ), .A2(
        \sha1_round/add_79_2/n285 ), .A3(\sha1_round/add_79_2/n286 ), .ZN(
        \sha1_round/add_79_2/n283 ) );
  NOR2_X2 \sha1_round/add_79_2/U39  ( .A1(\sha1_round/add_79_2/n35 ), .A2(
        \sha1_round/add_79_2/n61 ), .ZN(\sha1_round/add_79_2/n18 ) );
  XOR2_X2 \sha1_round/add_79_2/U38  ( .A(\sha1_round/add_79_2/n67 ), .B(
        \sha1_round/add_79_2/n18 ), .Z(\sha1_round/N290 ) );
  NOR2_X1 \sha1_round/add_79_2/U37  ( .A1(\sha1_round/add_79_2/n215 ), .A2(
        \sha1_round/add_79_2/n197 ), .ZN(\sha1_round/add_79_2/n214 ) );
  NOR2_X1 \sha1_round/add_79_2/U36  ( .A1(\sha1_round/add_79_2/n264 ), .A2(
        \sha1_round/add_79_2/n49 ), .ZN(\sha1_round/add_79_2/n317 ) );
  NOR2_X1 \sha1_round/add_79_2/U35  ( .A1(\sha1_round/add_79_2/n264 ), .A2(
        \sha1_round/add_79_2/n72 ), .ZN(\sha1_round/add_79_2/n293 ) );
  NAND3_X1 \sha1_round/add_79_2/U34  ( .A1(\sha1_round/add_79_2/n261 ), .A2(
        \sha1_round/add_79_2/n262 ), .A3(\sha1_round/add_79_2/n263 ), .ZN(
        \sha1_round/add_79_2/n260 ) );
  NOR2_X1 \sha1_round/add_79_2/U33  ( .A1(\sha1_round/add_79_2/n264 ), .A2(
        \sha1_round/add_79_2/n265 ), .ZN(\sha1_round/add_79_2/n263 ) );
  NOR2_X2 \sha1_round/add_79_2/U32  ( .A1(\sha1_round/add_79_2/n162 ), .A2(
        \sha1_round/add_79_2/n163 ), .ZN(\sha1_round/add_79_2/n17 ) );
  XOR2_X2 \sha1_round/add_79_2/U31  ( .A(\sha1_round/add_79_2/n17 ), .B(
        \sha1_round/add_79_2/n159 ), .Z(\sha1_round/N310 ) );
  NAND2_X1 \sha1_round/add_79_2/U30  ( .A1(\sha1_round/add_79_2/n171 ), .A2(
        \sha1_round/add_79_2/n180 ), .ZN(\sha1_round/add_79_2/n141 ) );
  NOR2_X2 \sha1_round/add_79_2/U29  ( .A1(\sha1_round/add_79_2/n192 ), .A2(
        \sha1_round/add_79_2/n183 ), .ZN(\sha1_round/add_79_2/n16 ) );
  XOR2_X2 \sha1_round/add_79_2/U28  ( .A(\sha1_round/add_79_2/n16 ), .B(
        \sha1_round/add_79_2/n189 ), .Z(\sha1_round/N307 ) );
  NOR2_X2 \sha1_round/add_79_2/U27  ( .A1(\sha1_round/add_79_2/n84 ), .A2(
        \sha1_round/add_79_2/n36 ), .ZN(\sha1_round/add_79_2/n15 ) );
  XOR2_X2 \sha1_round/add_79_2/U26  ( .A(\sha1_round/add_79_2/n15 ), .B(
        \sha1_round/add_79_2/n82 ), .Z(\sha1_round/N287 ) );
  NOR2_X2 \sha1_round/add_79_2/U25  ( .A1(\sha1_round/add_79_2/n305 ), .A2(
        \sha1_round/add_79_2/n306 ), .ZN(\sha1_round/add_79_2/n14 ) );
  XOR2_X2 \sha1_round/add_79_2/U24  ( .A(\sha1_round/add_79_2/n14 ), .B(
        \sha1_round/add_79_2/n302 ), .Z(\sha1_round/N299 ) );
  NOR2_X1 \sha1_round/add_79_2/U23  ( .A1(\sha1_round/add_79_2/n340 ), .A2(
        \sha1_round/add_79_2/n37 ), .ZN(\sha1_round/add_79_2/n345 ) );
  NOR2_X2 \sha1_round/add_79_2/U22  ( .A1(\sha1_round/add_79_2/n241 ), .A2(
        \sha1_round/add_79_2/n237 ), .ZN(\sha1_round/add_79_2/n13 ) );
  XOR2_X2 \sha1_round/add_79_2/U21  ( .A(\sha1_round/add_79_2/n13 ), .B(
        \sha1_round/add_79_2/n238 ), .Z(\sha1_round/N302 ) );
  NAND3_X1 \sha1_round/add_79_2/U20  ( .A1(\sha1_round/add_79_2/n360 ), .A2(
        \sha1_round/add_79_2/n262 ), .A3(\sha1_round/add_79_2/n361 ), .ZN(
        \sha1_round/add_79_2/n359 ) );
  NOR2_X1 \sha1_round/add_79_2/U19  ( .A1(\sha1_round/add_79_2/n56 ), .A2(
        \sha1_round/add_79_2/n57 ), .ZN(\sha1_round/add_79_2/n55 ) );
  NOR2_X1 \sha1_round/add_79_2/U18  ( .A1(\sha1_round/add_79_2/n321 ), .A2(
        \sha1_round/add_79_2/n264 ), .ZN(\sha1_round/add_79_2/n320 ) );
  NOR2_X1 \sha1_round/add_79_2/U17  ( .A1(\sha1_round/add_79_2/n264 ), .A2(
        \sha1_round/add_79_2/n275 ), .ZN(\sha1_round/add_79_2/n274 ) );
  NAND2_X1 \sha1_round/add_79_2/U16  ( .A1(\sha1_round/add_79_2/n5 ), .A2(
        \sha1_round/add_79_2/n118 ), .ZN(\sha1_round/add_79_2/n218 ) );
  NAND2_X1 \sha1_round/add_79_2/U15  ( .A1(\sha1_round/add_79_2/n5 ), .A2(
        \sha1_round/add_79_2/n118 ), .ZN(\sha1_round/add_79_2/n117 ) );
  NAND3_X2 \sha1_round/add_79_2/U14  ( .A1(\sha1_round/add_79_2/n363 ), .A2(
        \sha1_round/add_79_2/n71 ), .A3(\sha1_round/add_79_2/n364 ), .ZN(
        \sha1_round/add_79_2/n49 ) );
  AND2_X4 \sha1_round/add_79_2/U13  ( .A1(\sha1_round/add_79_2/n283 ), .A2(
        \sha1_round/add_79_2/n284 ), .ZN(\sha1_round/add_79_2/n12 ) );
  OR2_X4 \sha1_round/add_79_2/U12  ( .A1(rnd_q[21]), .A2(w[21]), .ZN(
        \sha1_round/add_79_2/n11 ) );
  OR2_X4 \sha1_round/add_79_2/U11  ( .A1(\sha1_round/add_79_2/n48 ), .A2(
        \sha1_round/add_79_2/n331 ), .ZN(\sha1_round/add_79_2/n10 ) );
  AND2_X4 \sha1_round/add_79_2/U10  ( .A1(w[30]), .A2(rnd_q[30]), .ZN(
        \sha1_round/add_79_2/n9 ) );
  AND2_X4 \sha1_round/add_79_2/U9  ( .A1(\sha1_round/add_79_2/n185 ), .A2(
        \sha1_round/add_79_2/n186 ), .ZN(\sha1_round/add_79_2/n8 ) );
  AND2_X4 \sha1_round/add_79_2/U8  ( .A1(w[20]), .A2(rnd_q[20]), .ZN(
        \sha1_round/add_79_2/n7 ) );
  AND2_X4 \sha1_round/add_79_2/U7  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(
        \sha1_round/add_79_2/n6 ) );
  AND2_X4 \sha1_round/add_79_2/U6  ( .A1(\sha1_round/add_79_2/n219 ), .A2(
        \sha1_round/add_79_2/n186 ), .ZN(\sha1_round/add_79_2/n5 ) );
  AND2_X4 \sha1_round/add_79_2/U5  ( .A1(\sha1_round/add_79_2/n101 ), .A2(
        \sha1_round/add_79_2/n102 ), .ZN(\sha1_round/add_79_2/n4 ) );
  AND2_X4 \sha1_round/add_79_2/U4  ( .A1(\sha1_round/add_79_2/n2 ), .A2(
        \sha1_round/add_79_2/n115 ), .ZN(\sha1_round/add_79_2/n3 ) );
  AND2_X4 \sha1_round/add_79_2/U3  ( .A1(\sha1_round/add_79_2/n187 ), .A2(
        \sha1_round/add_79_2/n184 ), .ZN(\sha1_round/add_79_2/n2 ) );
  AND2_X4 \sha1_round/add_79_2/U2  ( .A1(\sha1_round/add_79_2/n120 ), .A2(
        \sha1_round/add_79_2/n115 ), .ZN(\sha1_round/add_79_2/n1 ) );
  AND2_X2 \rnd_cnt_reg/U15  ( .A1(rnd_cnt_d[6]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N9 ) );
  AND2_X2 \rnd_cnt_reg/U14  ( .A1(rnd_cnt_d[5]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N8 ) );
  AND2_X2 \rnd_cnt_reg/U13  ( .A1(rnd_cnt_d[4]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N7 ) );
  AND2_X2 \rnd_cnt_reg/U12  ( .A1(rnd_cnt_d[3]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N6 ) );
  INV_X4 \rnd_cnt_reg/U11  ( .A(\rnd_cnt_reg/n70 ), .ZN(rnd_cnt_q[2]) );
  INV_X4 \rnd_cnt_reg/U10  ( .A(\rnd_cnt_reg/n40 ), .ZN(rnd_cnt_q[3]) );
  INV_X1 \rnd_cnt_reg/U7  ( .A(n7117), .ZN(\rnd_cnt_reg/n12 ) );
  AND2_X4 \rnd_cnt_reg/U6  ( .A1(rnd_cnt_d[2]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N5 ) );
  INV_X4 \rnd_cnt_reg/U5  ( .A(\rnd_cnt_reg/n60 ), .ZN(rnd_cnt_q[5]) );
  INV_X4 \rnd_cnt_reg/U4  ( .A(\rnd_cnt_reg/n2 ), .ZN(rnd_cnt_q[6]) );
  INV_X8 \rnd_cnt_reg/U3  ( .A(\rnd_cnt_reg/n10 ), .ZN(rnd_cnt_q[4]) );
  DFF_X2 \rnd_cnt_reg/q_reg_5_  ( .D(\rnd_cnt_reg/N8 ), .CK(clk), .Q(), .QN(
        \rnd_cnt_reg/n60 ) );
  DFF_X2 \rnd_cnt_reg/q_reg_4_  ( .D(\rnd_cnt_reg/N7 ), .CK(clk), .Q(), .QN(
        \rnd_cnt_reg/n10 ) );
  DFF_X1 \rnd_cnt_reg/q_reg_6_  ( .D(\rnd_cnt_reg/N9 ), .CK(clk), .Q(), .QN(
        \rnd_cnt_reg/n2 ) );
  DFF_X2 \rnd_cnt_reg/q_reg_2_  ( .D(\rnd_cnt_reg/N5 ), .CK(clk), .Q(), .QN(
        \rnd_cnt_reg/n70 ) );
  AND2_X2 \rnd_cnt_reg/U9  ( .A1(rnd_cnt_d[0]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N3 ) );
  AND2_X2 \rnd_cnt_reg/U8  ( .A1(rnd_cnt_d[1]), .A2(\rnd_cnt_reg/n12 ), .ZN(
        \rnd_cnt_reg/N4 ) );
  DFF_X2 \rnd_cnt_reg/q_reg_0_  ( .D(\rnd_cnt_reg/N3 ), .CK(clk), .Q(
        rnd_cnt_q[0]), .QN() );
  DFF_X2 \rnd_cnt_reg/q_reg_1_  ( .D(\rnd_cnt_reg/N4 ), .CK(clk), .Q(
        rnd_cnt_q[1]), .QN() );
  DFF_X2 \rnd_cnt_reg/q_reg_3_  ( .D(\rnd_cnt_reg/N6 ), .CK(clk), .Q(), .QN(
        \rnd_cnt_reg/n40 ) );
  INV_X4 \state_reg/U5  ( .A(n7117), .ZN(\state_reg/n2 ) );
  AND2_X4 \state_reg/U3  ( .A1(next_state[1]), .A2(\state_reg/n2 ), .ZN(
        \state_reg/N4 ) );
  AND2_X2 \state_reg/U4  ( .A1(next_state[0]), .A2(\state_reg/n2 ), .ZN(
        \state_reg/N3 ) );
  DFF_X2 \state_reg/q_reg_0_  ( .D(\state_reg/N3 ), .CK(clk), .Q(state[0]), 
        .QN() );
  DFF_X2 \state_reg/q_reg_1_  ( .D(\state_reg/N4 ), .CK(clk), .Q(state[1]), 
        .QN() );
  AND2_X2 \w_reg/U562  ( .A1(w_d[497]), .A2(\w_reg/n610 ), .ZN(\w_reg/N500 )
         );
  AND2_X2 \w_reg/U561  ( .A1(w_d[496]), .A2(\w_reg/n610 ), .ZN(\w_reg/N499 )
         );
  AND2_X2 \w_reg/U560  ( .A1(w_d[495]), .A2(\w_reg/n610 ), .ZN(\w_reg/N498 )
         );
  AND2_X2 \w_reg/U559  ( .A1(w_d[494]), .A2(\w_reg/n610 ), .ZN(\w_reg/N497 )
         );
  AND2_X2 \w_reg/U558  ( .A1(w_d[493]), .A2(\w_reg/n610 ), .ZN(\w_reg/N496 )
         );
  AND2_X2 \w_reg/U557  ( .A1(w_d[492]), .A2(\w_reg/n610 ), .ZN(\w_reg/N495 )
         );
  AND2_X2 \w_reg/U556  ( .A1(w_d[491]), .A2(\w_reg/n610 ), .ZN(\w_reg/N494 )
         );
  AND2_X2 \w_reg/U555  ( .A1(w_d[490]), .A2(\w_reg/n600 ), .ZN(\w_reg/N493 )
         );
  AND2_X2 \w_reg/U554  ( .A1(w_d[489]), .A2(\w_reg/n600 ), .ZN(\w_reg/N492 )
         );
  AND2_X2 \w_reg/U553  ( .A1(w_d[488]), .A2(\w_reg/n600 ), .ZN(\w_reg/N491 )
         );
  AND2_X2 \w_reg/U552  ( .A1(w_d[487]), .A2(\w_reg/n600 ), .ZN(\w_reg/N490 )
         );
  AND2_X2 \w_reg/U551  ( .A1(w_d[486]), .A2(\w_reg/n600 ), .ZN(\w_reg/N489 )
         );
  AND2_X2 \w_reg/U550  ( .A1(w_d[485]), .A2(\w_reg/n600 ), .ZN(\w_reg/N488 )
         );
  AND2_X2 \w_reg/U549  ( .A1(w_d[484]), .A2(\w_reg/n600 ), .ZN(\w_reg/N487 )
         );
  AND2_X2 \w_reg/U548  ( .A1(w_d[483]), .A2(\w_reg/n600 ), .ZN(\w_reg/N486 )
         );
  AND2_X2 \w_reg/U547  ( .A1(w_d[482]), .A2(\w_reg/n600 ), .ZN(\w_reg/N485 )
         );
  AND2_X2 \w_reg/U546  ( .A1(w_d[481]), .A2(\w_reg/n600 ), .ZN(\w_reg/N484 )
         );
  AND2_X2 \w_reg/U545  ( .A1(w_d[480]), .A2(\w_reg/n600 ), .ZN(\w_reg/N483 )
         );
  INV_X4 \w_reg/U544  ( .A(reset), .ZN(\w_reg/n1070 ) );
  BUF_X4 \w_reg/U543  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1060 ) );
  BUF_X4 \w_reg/U542  ( .A(\w_reg/n1070 ), .Z(\w_reg/n660 ) );
  BUF_X4 \w_reg/U541  ( .A(\w_reg/n1070 ), .Z(\w_reg/n670 ) );
  BUF_X4 \w_reg/U540  ( .A(\w_reg/n1070 ), .Z(\w_reg/n610 ) );
  BUF_X4 \w_reg/U539  ( .A(\w_reg/n1070 ), .Z(\w_reg/n600 ) );
  BUF_X4 \w_reg/U538  ( .A(\w_reg/n1070 ), .Z(\w_reg/n680 ) );
  BUF_X4 \w_reg/U537  ( .A(\w_reg/n1070 ), .Z(\w_reg/n690 ) );
  BUF_X4 \w_reg/U536  ( .A(\w_reg/n1070 ), .Z(\w_reg/n700 ) );
  BUF_X4 \w_reg/U535  ( .A(\w_reg/n1070 ), .Z(\w_reg/n710 ) );
  BUF_X4 \w_reg/U534  ( .A(\w_reg/n1070 ), .Z(\w_reg/n720 ) );
  BUF_X4 \w_reg/U533  ( .A(\w_reg/n1070 ), .Z(\w_reg/n730 ) );
  BUF_X4 \w_reg/U532  ( .A(\w_reg/n1070 ), .Z(\w_reg/n740 ) );
  BUF_X4 \w_reg/U531  ( .A(\w_reg/n1070 ), .Z(\w_reg/n750 ) );
  BUF_X4 \w_reg/U530  ( .A(\w_reg/n1070 ), .Z(\w_reg/n760 ) );
  BUF_X4 \w_reg/U529  ( .A(\w_reg/n1070 ), .Z(\w_reg/n770 ) );
  BUF_X4 \w_reg/U528  ( .A(\w_reg/n1070 ), .Z(\w_reg/n780 ) );
  BUF_X4 \w_reg/U527  ( .A(\w_reg/n1070 ), .Z(\w_reg/n790 ) );
  BUF_X4 \w_reg/U526  ( .A(\w_reg/n1070 ), .Z(\w_reg/n800 ) );
  BUF_X4 \w_reg/U525  ( .A(\w_reg/n1070 ), .Z(\w_reg/n810 ) );
  BUF_X4 \w_reg/U524  ( .A(\w_reg/n1070 ), .Z(\w_reg/n820 ) );
  BUF_X4 \w_reg/U523  ( .A(\w_reg/n1070 ), .Z(\w_reg/n830 ) );
  BUF_X4 \w_reg/U522  ( .A(\w_reg/n1070 ), .Z(\w_reg/n840 ) );
  BUF_X4 \w_reg/U521  ( .A(\w_reg/n1070 ), .Z(\w_reg/n850 ) );
  BUF_X4 \w_reg/U520  ( .A(\w_reg/n1070 ), .Z(\w_reg/n860 ) );
  BUF_X4 \w_reg/U519  ( .A(\w_reg/n1070 ), .Z(\w_reg/n870 ) );
  BUF_X4 \w_reg/U518  ( .A(\w_reg/n1070 ), .Z(\w_reg/n880 ) );
  BUF_X4 \w_reg/U517  ( .A(\w_reg/n1070 ), .Z(\w_reg/n890 ) );
  BUF_X4 \w_reg/U516  ( .A(\w_reg/n1070 ), .Z(\w_reg/n900 ) );
  BUF_X4 \w_reg/U515  ( .A(\w_reg/n1070 ), .Z(\w_reg/n910 ) );
  BUF_X4 \w_reg/U514  ( .A(\w_reg/n1070 ), .Z(\w_reg/n920 ) );
  BUF_X4 \w_reg/U503  ( .A(\w_reg/n1070 ), .Z(\w_reg/n930 ) );
  BUF_X4 \w_reg/U492  ( .A(\w_reg/n1070 ), .Z(\w_reg/n940 ) );
  BUF_X4 \w_reg/U481  ( .A(\w_reg/n1070 ), .Z(\w_reg/n950 ) );
  BUF_X4 \w_reg/U470  ( .A(\w_reg/n1070 ), .Z(\w_reg/n960 ) );
  BUF_X4 \w_reg/U459  ( .A(\w_reg/n1070 ), .Z(\w_reg/n970 ) );
  BUF_X4 \w_reg/U448  ( .A(\w_reg/n1070 ), .Z(\w_reg/n980 ) );
  BUF_X4 \w_reg/U437  ( .A(\w_reg/n1070 ), .Z(\w_reg/n990 ) );
  BUF_X4 \w_reg/U426  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1000 ) );
  BUF_X4 \w_reg/U415  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1010 ) );
  BUF_X4 \w_reg/U404  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1020 ) );
  BUF_X4 \w_reg/U393  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1030 ) );
  BUF_X4 \w_reg/U382  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1040 ) );
  BUF_X4 \w_reg/U371  ( .A(\w_reg/n1070 ), .Z(\w_reg/n1050 ) );
  BUF_X4 \w_reg/U360  ( .A(\w_reg/n1070 ), .Z(\w_reg/n620 ) );
  BUF_X4 \w_reg/U349  ( .A(\w_reg/n1070 ), .Z(\w_reg/n630 ) );
  BUF_X4 \w_reg/U338  ( .A(\w_reg/n1070 ), .Z(\w_reg/n640 ) );
  BUF_X4 \w_reg/U327  ( .A(\w_reg/n1070 ), .Z(\w_reg/n650 ) );
  AND2_X1 \w_reg/U316  ( .A1(w_d[31]), .A2(\w_reg/n820 ), .ZN(\w_reg/N34 ) );
  AND2_X1 \w_reg/U305  ( .A1(w_d[30]), .A2(\w_reg/n830 ), .ZN(\w_reg/N33 ) );
  AND2_X1 \w_reg/U294  ( .A1(w_d[29]), .A2(\w_reg/n840 ), .ZN(\w_reg/N32 ) );
  AND2_X1 \w_reg/U293  ( .A1(w_d[28]), .A2(\w_reg/n850 ), .ZN(\w_reg/N31 ) );
  AND2_X1 \w_reg/U282  ( .A1(w_d[27]), .A2(\w_reg/n860 ), .ZN(\w_reg/N30 ) );
  AND2_X1 \w_reg/U271  ( .A1(w_d[26]), .A2(\w_reg/n870 ), .ZN(\w_reg/N29 ) );
  AND2_X1 \w_reg/U260  ( .A1(w_d[25]), .A2(\w_reg/n880 ), .ZN(\w_reg/N28 ) );
  AND2_X1 \w_reg/U249  ( .A1(w_d[24]), .A2(\w_reg/n890 ), .ZN(\w_reg/N27 ) );
  AND2_X1 \w_reg/U183  ( .A1(w_d[23]), .A2(\w_reg/n900 ), .ZN(\w_reg/N26 ) );
  AND2_X1 \w_reg/U90  ( .A1(w_d[22]), .A2(\w_reg/n910 ), .ZN(\w_reg/N25 ) );
  AND2_X1 \w_reg/U89  ( .A1(w_d[21]), .A2(\w_reg/n920 ), .ZN(\w_reg/N24 ) );
  AND2_X1 \w_reg/U88  ( .A1(w_d[20]), .A2(\w_reg/n930 ), .ZN(\w_reg/N23 ) );
  AND2_X1 \w_reg/U87  ( .A1(w_d[19]), .A2(\w_reg/n940 ), .ZN(\w_reg/N22 ) );
  AND2_X1 \w_reg/U86  ( .A1(w_d[18]), .A2(\w_reg/n950 ), .ZN(\w_reg/N21 ) );
  AND2_X1 \w_reg/U85  ( .A1(w_d[17]), .A2(\w_reg/n960 ), .ZN(\w_reg/N20 ) );
  AND2_X1 \w_reg/U84  ( .A1(w_d[16]), .A2(\w_reg/n970 ), .ZN(\w_reg/N19 ) );
  AND2_X1 \w_reg/U82  ( .A1(w_d[15]), .A2(\w_reg/n980 ), .ZN(\w_reg/N18 ) );
  AND2_X1 \w_reg/U81  ( .A1(w_d[14]), .A2(\w_reg/n990 ), .ZN(\w_reg/N17 ) );
  AND2_X1 \w_reg/U80  ( .A1(w_d[13]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N16 ) );
  AND2_X1 \w_reg/U79  ( .A1(w_d[12]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N15 ) );
  AND2_X1 \w_reg/U78  ( .A1(w_d[11]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N14 ) );
  AND2_X1 \w_reg/U77  ( .A1(w_d[10]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N13 ) );
  AND2_X1 \w_reg/U76  ( .A1(w_d[9]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N12 ) );
  AND2_X1 \w_reg/U75  ( .A1(w_d[8]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N11 ) );
  AND2_X1 \w_reg/U74  ( .A1(w_d[7]), .A2(\w_reg/n1060 ), .ZN(\w_reg/N10 ) );
  AND2_X1 \w_reg/U73  ( .A1(w_d[6]), .A2(\w_reg/n620 ), .ZN(\w_reg/N9 ) );
  AND2_X1 \w_reg/U72  ( .A1(w_d[5]), .A2(\w_reg/n630 ), .ZN(\w_reg/N8 ) );
  AND2_X1 \w_reg/U70  ( .A1(w_d[4]), .A2(\w_reg/n640 ), .ZN(\w_reg/N7 ) );
  AND2_X1 \w_reg/U46  ( .A1(w_d[3]), .A2(\w_reg/n650 ), .ZN(\w_reg/N6 ) );
  AND2_X1 \w_reg/U35  ( .A1(w_d[2]), .A2(\w_reg/n670 ), .ZN(\w_reg/N5 ) );
  AND2_X1 \w_reg/U24  ( .A1(w_d[1]), .A2(\w_reg/n760 ), .ZN(\w_reg/N4 ) );
  AND2_X1 \w_reg/U13  ( .A1(w_d[0]), .A2(\w_reg/n860 ), .ZN(\w_reg/N3 ) );
  AND2_X2 \w_reg/U513  ( .A1(w_d[97]), .A2(\w_reg/n1060 ), .ZN(\w_reg/N100 )
         );
  AND2_X2 \w_reg/U512  ( .A1(w_d[98]), .A2(\w_reg/n1060 ), .ZN(\w_reg/N101 )
         );
  AND2_X2 \w_reg/U511  ( .A1(w_d[99]), .A2(\w_reg/n1060 ), .ZN(\w_reg/N102 )
         );
  AND2_X2 \w_reg/U510  ( .A1(w_d[100]), .A2(\w_reg/n1060 ), .ZN(\w_reg/N103 )
         );
  AND2_X2 \w_reg/U509  ( .A1(w_d[101]), .A2(\w_reg/n1060 ), .ZN(\w_reg/N104 )
         );
  AND2_X2 \w_reg/U508  ( .A1(w_d[102]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N105 )
         );
  AND2_X2 \w_reg/U507  ( .A1(w_d[103]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N106 )
         );
  AND2_X2 \w_reg/U506  ( .A1(w_d[104]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N107 )
         );
  AND2_X2 \w_reg/U505  ( .A1(w_d[105]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N108 )
         );
  AND2_X2 \w_reg/U504  ( .A1(w_d[106]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N109 )
         );
  AND2_X2 \w_reg/U502  ( .A1(w_d[107]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N110 )
         );
  AND2_X2 \w_reg/U501  ( .A1(w_d[108]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N111 )
         );
  AND2_X2 \w_reg/U500  ( .A1(w_d[109]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N112 )
         );
  AND2_X2 \w_reg/U499  ( .A1(w_d[110]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N113 )
         );
  AND2_X2 \w_reg/U498  ( .A1(w_d[111]), .A2(\w_reg/n1050 ), .ZN(\w_reg/N114 )
         );
  AND2_X2 \w_reg/U497  ( .A1(w_d[112]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N115 )
         );
  AND2_X2 \w_reg/U496  ( .A1(w_d[113]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N116 )
         );
  AND2_X2 \w_reg/U495  ( .A1(w_d[114]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N117 )
         );
  AND2_X2 \w_reg/U494  ( .A1(w_d[115]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N118 )
         );
  AND2_X2 \w_reg/U493  ( .A1(w_d[116]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N119 )
         );
  AND2_X2 \w_reg/U491  ( .A1(w_d[117]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N120 )
         );
  AND2_X2 \w_reg/U490  ( .A1(w_d[118]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N121 )
         );
  AND2_X2 \w_reg/U489  ( .A1(w_d[119]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N122 )
         );
  AND2_X2 \w_reg/U488  ( .A1(w_d[120]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N123 )
         );
  AND2_X2 \w_reg/U487  ( .A1(w_d[121]), .A2(\w_reg/n1040 ), .ZN(\w_reg/N124 )
         );
  AND2_X2 \w_reg/U486  ( .A1(w_d[122]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N125 )
         );
  AND2_X2 \w_reg/U485  ( .A1(w_d[123]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N126 )
         );
  AND2_X2 \w_reg/U484  ( .A1(w_d[124]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N127 )
         );
  AND2_X2 \w_reg/U483  ( .A1(w_d[125]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N128 )
         );
  AND2_X2 \w_reg/U482  ( .A1(w_d[126]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N129 )
         );
  AND2_X2 \w_reg/U480  ( .A1(w_d[127]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N130 )
         );
  AND2_X2 \w_reg/U479  ( .A1(w_d[128]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N131 )
         );
  AND2_X2 \w_reg/U478  ( .A1(w_d[129]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N132 )
         );
  AND2_X2 \w_reg/U477  ( .A1(w_d[130]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N133 )
         );
  AND2_X2 \w_reg/U476  ( .A1(w_d[131]), .A2(\w_reg/n1030 ), .ZN(\w_reg/N134 )
         );
  AND2_X2 \w_reg/U475  ( .A1(w_d[132]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N135 )
         );
  AND2_X2 \w_reg/U474  ( .A1(w_d[133]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N136 )
         );
  AND2_X2 \w_reg/U473  ( .A1(w_d[134]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N137 )
         );
  AND2_X2 \w_reg/U472  ( .A1(w_d[135]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N138 )
         );
  AND2_X2 \w_reg/U471  ( .A1(w_d[136]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N139 )
         );
  AND2_X2 \w_reg/U469  ( .A1(w_d[137]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N140 )
         );
  AND2_X2 \w_reg/U468  ( .A1(w_d[138]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N141 )
         );
  AND2_X2 \w_reg/U467  ( .A1(w_d[139]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N142 )
         );
  AND2_X2 \w_reg/U466  ( .A1(w_d[140]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N143 )
         );
  AND2_X2 \w_reg/U465  ( .A1(w_d[141]), .A2(\w_reg/n1020 ), .ZN(\w_reg/N144 )
         );
  AND2_X2 \w_reg/U464  ( .A1(w_d[142]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N145 )
         );
  AND2_X2 \w_reg/U463  ( .A1(w_d[143]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N146 )
         );
  AND2_X2 \w_reg/U462  ( .A1(w_d[144]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N147 )
         );
  AND2_X2 \w_reg/U461  ( .A1(w_d[145]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N148 )
         );
  AND2_X2 \w_reg/U460  ( .A1(w_d[146]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N149 )
         );
  AND2_X2 \w_reg/U458  ( .A1(w_d[147]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N150 )
         );
  AND2_X2 \w_reg/U457  ( .A1(w_d[148]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N151 )
         );
  AND2_X2 \w_reg/U456  ( .A1(w_d[149]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N152 )
         );
  AND2_X2 \w_reg/U455  ( .A1(w_d[150]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N153 )
         );
  AND2_X2 \w_reg/U454  ( .A1(w_d[151]), .A2(\w_reg/n1010 ), .ZN(\w_reg/N154 )
         );
  AND2_X2 \w_reg/U453  ( .A1(w_d[152]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N155 )
         );
  AND2_X2 \w_reg/U452  ( .A1(w_d[153]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N156 )
         );
  AND2_X2 \w_reg/U451  ( .A1(w_d[154]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N157 )
         );
  AND2_X2 \w_reg/U450  ( .A1(w_d[155]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N158 )
         );
  AND2_X2 \w_reg/U449  ( .A1(w_d[156]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N159 )
         );
  AND2_X2 \w_reg/U447  ( .A1(w_d[157]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N160 )
         );
  AND2_X2 \w_reg/U446  ( .A1(w_d[158]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N161 )
         );
  AND2_X2 \w_reg/U445  ( .A1(w_d[159]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N162 )
         );
  AND2_X2 \w_reg/U444  ( .A1(w_d[160]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N163 )
         );
  AND2_X2 \w_reg/U443  ( .A1(w_d[161]), .A2(\w_reg/n1000 ), .ZN(\w_reg/N164 )
         );
  AND2_X2 \w_reg/U442  ( .A1(w_d[162]), .A2(\w_reg/n990 ), .ZN(\w_reg/N165 )
         );
  AND2_X2 \w_reg/U441  ( .A1(w_d[163]), .A2(\w_reg/n990 ), .ZN(\w_reg/N166 )
         );
  AND2_X2 \w_reg/U440  ( .A1(w_d[164]), .A2(\w_reg/n990 ), .ZN(\w_reg/N167 )
         );
  AND2_X2 \w_reg/U439  ( .A1(w_d[165]), .A2(\w_reg/n990 ), .ZN(\w_reg/N168 )
         );
  AND2_X2 \w_reg/U438  ( .A1(w_d[166]), .A2(\w_reg/n990 ), .ZN(\w_reg/N169 )
         );
  AND2_X2 \w_reg/U436  ( .A1(w_d[167]), .A2(\w_reg/n990 ), .ZN(\w_reg/N170 )
         );
  AND2_X2 \w_reg/U435  ( .A1(w_d[168]), .A2(\w_reg/n990 ), .ZN(\w_reg/N171 )
         );
  AND2_X2 \w_reg/U434  ( .A1(w_d[169]), .A2(\w_reg/n990 ), .ZN(\w_reg/N172 )
         );
  AND2_X2 \w_reg/U433  ( .A1(w_d[170]), .A2(\w_reg/n990 ), .ZN(\w_reg/N173 )
         );
  AND2_X2 \w_reg/U432  ( .A1(w_d[171]), .A2(\w_reg/n990 ), .ZN(\w_reg/N174 )
         );
  AND2_X2 \w_reg/U431  ( .A1(w_d[172]), .A2(\w_reg/n980 ), .ZN(\w_reg/N175 )
         );
  AND2_X2 \w_reg/U430  ( .A1(w_d[173]), .A2(\w_reg/n980 ), .ZN(\w_reg/N176 )
         );
  AND2_X2 \w_reg/U429  ( .A1(w_d[174]), .A2(\w_reg/n980 ), .ZN(\w_reg/N177 )
         );
  AND2_X2 \w_reg/U428  ( .A1(w_d[175]), .A2(\w_reg/n980 ), .ZN(\w_reg/N178 )
         );
  AND2_X2 \w_reg/U427  ( .A1(w_d[176]), .A2(\w_reg/n980 ), .ZN(\w_reg/N179 )
         );
  AND2_X2 \w_reg/U425  ( .A1(w_d[177]), .A2(\w_reg/n980 ), .ZN(\w_reg/N180 )
         );
  AND2_X2 \w_reg/U424  ( .A1(w_d[178]), .A2(\w_reg/n980 ), .ZN(\w_reg/N181 )
         );
  AND2_X2 \w_reg/U423  ( .A1(w_d[179]), .A2(\w_reg/n980 ), .ZN(\w_reg/N182 )
         );
  AND2_X2 \w_reg/U422  ( .A1(w_d[180]), .A2(\w_reg/n980 ), .ZN(\w_reg/N183 )
         );
  AND2_X2 \w_reg/U421  ( .A1(w_d[181]), .A2(\w_reg/n980 ), .ZN(\w_reg/N184 )
         );
  AND2_X2 \w_reg/U420  ( .A1(w_d[182]), .A2(\w_reg/n970 ), .ZN(\w_reg/N185 )
         );
  AND2_X2 \w_reg/U419  ( .A1(w_d[183]), .A2(\w_reg/n970 ), .ZN(\w_reg/N186 )
         );
  AND2_X2 \w_reg/U418  ( .A1(w_d[184]), .A2(\w_reg/n970 ), .ZN(\w_reg/N187 )
         );
  AND2_X2 \w_reg/U417  ( .A1(w_d[185]), .A2(\w_reg/n970 ), .ZN(\w_reg/N188 )
         );
  AND2_X2 \w_reg/U416  ( .A1(w_d[186]), .A2(\w_reg/n970 ), .ZN(\w_reg/N189 )
         );
  AND2_X2 \w_reg/U414  ( .A1(w_d[187]), .A2(\w_reg/n970 ), .ZN(\w_reg/N190 )
         );
  AND2_X2 \w_reg/U413  ( .A1(w_d[188]), .A2(\w_reg/n970 ), .ZN(\w_reg/N191 )
         );
  AND2_X2 \w_reg/U412  ( .A1(w_d[189]), .A2(\w_reg/n970 ), .ZN(\w_reg/N192 )
         );
  AND2_X2 \w_reg/U411  ( .A1(w_d[190]), .A2(\w_reg/n970 ), .ZN(\w_reg/N193 )
         );
  AND2_X2 \w_reg/U410  ( .A1(w_d[191]), .A2(\w_reg/n970 ), .ZN(\w_reg/N194 )
         );
  AND2_X2 \w_reg/U409  ( .A1(w_d[192]), .A2(\w_reg/n960 ), .ZN(\w_reg/N195 )
         );
  AND2_X2 \w_reg/U408  ( .A1(w_d[193]), .A2(\w_reg/n960 ), .ZN(\w_reg/N196 )
         );
  AND2_X2 \w_reg/U407  ( .A1(w_d[194]), .A2(\w_reg/n960 ), .ZN(\w_reg/N197 )
         );
  AND2_X2 \w_reg/U406  ( .A1(w_d[195]), .A2(\w_reg/n960 ), .ZN(\w_reg/N198 )
         );
  AND2_X2 \w_reg/U405  ( .A1(w_d[196]), .A2(\w_reg/n960 ), .ZN(\w_reg/N199 )
         );
  AND2_X2 \w_reg/U403  ( .A1(w_d[197]), .A2(\w_reg/n960 ), .ZN(\w_reg/N200 )
         );
  AND2_X2 \w_reg/U402  ( .A1(w_d[198]), .A2(\w_reg/n960 ), .ZN(\w_reg/N201 )
         );
  AND2_X2 \w_reg/U401  ( .A1(w_d[199]), .A2(\w_reg/n960 ), .ZN(\w_reg/N202 )
         );
  AND2_X2 \w_reg/U400  ( .A1(w_d[200]), .A2(\w_reg/n960 ), .ZN(\w_reg/N203 )
         );
  AND2_X2 \w_reg/U399  ( .A1(w_d[201]), .A2(\w_reg/n960 ), .ZN(\w_reg/N204 )
         );
  AND2_X2 \w_reg/U398  ( .A1(w_d[202]), .A2(\w_reg/n950 ), .ZN(\w_reg/N205 )
         );
  AND2_X2 \w_reg/U397  ( .A1(w_d[203]), .A2(\w_reg/n950 ), .ZN(\w_reg/N206 )
         );
  AND2_X2 \w_reg/U396  ( .A1(w_d[204]), .A2(\w_reg/n950 ), .ZN(\w_reg/N207 )
         );
  AND2_X2 \w_reg/U395  ( .A1(w_d[205]), .A2(\w_reg/n950 ), .ZN(\w_reg/N208 )
         );
  AND2_X2 \w_reg/U394  ( .A1(w_d[206]), .A2(\w_reg/n950 ), .ZN(\w_reg/N209 )
         );
  AND2_X2 \w_reg/U392  ( .A1(w_d[207]), .A2(\w_reg/n950 ), .ZN(\w_reg/N210 )
         );
  AND2_X2 \w_reg/U391  ( .A1(w_d[208]), .A2(\w_reg/n950 ), .ZN(\w_reg/N211 )
         );
  AND2_X2 \w_reg/U390  ( .A1(w_d[209]), .A2(\w_reg/n950 ), .ZN(\w_reg/N212 )
         );
  AND2_X2 \w_reg/U389  ( .A1(w_d[210]), .A2(\w_reg/n950 ), .ZN(\w_reg/N213 )
         );
  AND2_X2 \w_reg/U388  ( .A1(w_d[211]), .A2(\w_reg/n950 ), .ZN(\w_reg/N214 )
         );
  AND2_X2 \w_reg/U387  ( .A1(w_d[212]), .A2(\w_reg/n940 ), .ZN(\w_reg/N215 )
         );
  AND2_X2 \w_reg/U386  ( .A1(w_d[213]), .A2(\w_reg/n940 ), .ZN(\w_reg/N216 )
         );
  AND2_X2 \w_reg/U385  ( .A1(w_d[214]), .A2(\w_reg/n940 ), .ZN(\w_reg/N217 )
         );
  AND2_X2 \w_reg/U384  ( .A1(w_d[215]), .A2(\w_reg/n940 ), .ZN(\w_reg/N218 )
         );
  AND2_X2 \w_reg/U383  ( .A1(w_d[216]), .A2(\w_reg/n940 ), .ZN(\w_reg/N219 )
         );
  AND2_X2 \w_reg/U381  ( .A1(w_d[217]), .A2(\w_reg/n940 ), .ZN(\w_reg/N220 )
         );
  AND2_X2 \w_reg/U380  ( .A1(w_d[218]), .A2(\w_reg/n940 ), .ZN(\w_reg/N221 )
         );
  AND2_X2 \w_reg/U379  ( .A1(w_d[219]), .A2(\w_reg/n940 ), .ZN(\w_reg/N222 )
         );
  AND2_X2 \w_reg/U378  ( .A1(w_d[220]), .A2(\w_reg/n940 ), .ZN(\w_reg/N223 )
         );
  AND2_X2 \w_reg/U377  ( .A1(w_d[221]), .A2(\w_reg/n940 ), .ZN(\w_reg/N224 )
         );
  AND2_X2 \w_reg/U376  ( .A1(w_d[222]), .A2(\w_reg/n930 ), .ZN(\w_reg/N225 )
         );
  AND2_X2 \w_reg/U375  ( .A1(w_d[223]), .A2(\w_reg/n930 ), .ZN(\w_reg/N226 )
         );
  AND2_X2 \w_reg/U374  ( .A1(w_d[224]), .A2(\w_reg/n930 ), .ZN(\w_reg/N227 )
         );
  AND2_X2 \w_reg/U373  ( .A1(w_d[225]), .A2(\w_reg/n930 ), .ZN(\w_reg/N228 )
         );
  AND2_X2 \w_reg/U372  ( .A1(w_d[226]), .A2(\w_reg/n930 ), .ZN(\w_reg/N229 )
         );
  AND2_X2 \w_reg/U370  ( .A1(w_d[227]), .A2(\w_reg/n930 ), .ZN(\w_reg/N230 )
         );
  AND2_X2 \w_reg/U369  ( .A1(w_d[228]), .A2(\w_reg/n930 ), .ZN(\w_reg/N231 )
         );
  AND2_X2 \w_reg/U368  ( .A1(w_d[229]), .A2(\w_reg/n930 ), .ZN(\w_reg/N232 )
         );
  AND2_X2 \w_reg/U367  ( .A1(w_d[230]), .A2(\w_reg/n930 ), .ZN(\w_reg/N233 )
         );
  AND2_X2 \w_reg/U366  ( .A1(w_d[231]), .A2(\w_reg/n930 ), .ZN(\w_reg/N234 )
         );
  AND2_X2 \w_reg/U365  ( .A1(w_d[232]), .A2(\w_reg/n920 ), .ZN(\w_reg/N235 )
         );
  AND2_X2 \w_reg/U364  ( .A1(w_d[233]), .A2(\w_reg/n920 ), .ZN(\w_reg/N236 )
         );
  AND2_X2 \w_reg/U363  ( .A1(w_d[234]), .A2(\w_reg/n920 ), .ZN(\w_reg/N237 )
         );
  AND2_X2 \w_reg/U362  ( .A1(w_d[235]), .A2(\w_reg/n920 ), .ZN(\w_reg/N238 )
         );
  AND2_X2 \w_reg/U361  ( .A1(w_d[236]), .A2(\w_reg/n920 ), .ZN(\w_reg/N239 )
         );
  AND2_X2 \w_reg/U359  ( .A1(w_d[237]), .A2(\w_reg/n920 ), .ZN(\w_reg/N240 )
         );
  AND2_X2 \w_reg/U358  ( .A1(w_d[238]), .A2(\w_reg/n920 ), .ZN(\w_reg/N241 )
         );
  AND2_X2 \w_reg/U357  ( .A1(w_d[239]), .A2(\w_reg/n920 ), .ZN(\w_reg/N242 )
         );
  AND2_X2 \w_reg/U356  ( .A1(w_d[240]), .A2(\w_reg/n920 ), .ZN(\w_reg/N243 )
         );
  AND2_X2 \w_reg/U355  ( .A1(w_d[241]), .A2(\w_reg/n920 ), .ZN(\w_reg/N244 )
         );
  AND2_X2 \w_reg/U354  ( .A1(w_d[242]), .A2(\w_reg/n910 ), .ZN(\w_reg/N245 )
         );
  AND2_X2 \w_reg/U353  ( .A1(w_d[243]), .A2(\w_reg/n910 ), .ZN(\w_reg/N246 )
         );
  AND2_X2 \w_reg/U352  ( .A1(w_d[244]), .A2(\w_reg/n910 ), .ZN(\w_reg/N247 )
         );
  AND2_X2 \w_reg/U351  ( .A1(w_d[245]), .A2(\w_reg/n910 ), .ZN(\w_reg/N248 )
         );
  AND2_X2 \w_reg/U350  ( .A1(w_d[246]), .A2(\w_reg/n910 ), .ZN(\w_reg/N249 )
         );
  AND2_X2 \w_reg/U348  ( .A1(w_d[247]), .A2(\w_reg/n910 ), .ZN(\w_reg/N250 )
         );
  AND2_X2 \w_reg/U347  ( .A1(w_d[248]), .A2(\w_reg/n910 ), .ZN(\w_reg/N251 )
         );
  AND2_X2 \w_reg/U346  ( .A1(w_d[249]), .A2(\w_reg/n910 ), .ZN(\w_reg/N252 )
         );
  AND2_X2 \w_reg/U345  ( .A1(w_d[250]), .A2(\w_reg/n910 ), .ZN(\w_reg/N253 )
         );
  AND2_X2 \w_reg/U344  ( .A1(w_d[251]), .A2(\w_reg/n910 ), .ZN(\w_reg/N254 )
         );
  AND2_X2 \w_reg/U343  ( .A1(w_d[252]), .A2(\w_reg/n900 ), .ZN(\w_reg/N255 )
         );
  AND2_X2 \w_reg/U342  ( .A1(w_d[253]), .A2(\w_reg/n900 ), .ZN(\w_reg/N256 )
         );
  AND2_X2 \w_reg/U341  ( .A1(w_d[254]), .A2(\w_reg/n900 ), .ZN(\w_reg/N257 )
         );
  AND2_X2 \w_reg/U340  ( .A1(w_d[255]), .A2(\w_reg/n900 ), .ZN(\w_reg/N258 )
         );
  AND2_X2 \w_reg/U339  ( .A1(w_d[256]), .A2(\w_reg/n900 ), .ZN(\w_reg/N259 )
         );
  AND2_X2 \w_reg/U337  ( .A1(w_d[257]), .A2(\w_reg/n900 ), .ZN(\w_reg/N260 )
         );
  AND2_X2 \w_reg/U336  ( .A1(w_d[258]), .A2(\w_reg/n900 ), .ZN(\w_reg/N261 )
         );
  AND2_X2 \w_reg/U335  ( .A1(w_d[259]), .A2(\w_reg/n900 ), .ZN(\w_reg/N262 )
         );
  AND2_X2 \w_reg/U334  ( .A1(w_d[260]), .A2(\w_reg/n900 ), .ZN(\w_reg/N263 )
         );
  AND2_X2 \w_reg/U333  ( .A1(w_d[261]), .A2(\w_reg/n900 ), .ZN(\w_reg/N264 )
         );
  AND2_X2 \w_reg/U332  ( .A1(w_d[262]), .A2(\w_reg/n890 ), .ZN(\w_reg/N265 )
         );
  AND2_X2 \w_reg/U331  ( .A1(w_d[263]), .A2(\w_reg/n890 ), .ZN(\w_reg/N266 )
         );
  AND2_X2 \w_reg/U330  ( .A1(w_d[264]), .A2(\w_reg/n890 ), .ZN(\w_reg/N267 )
         );
  AND2_X2 \w_reg/U329  ( .A1(w_d[265]), .A2(\w_reg/n890 ), .ZN(\w_reg/N268 )
         );
  AND2_X2 \w_reg/U328  ( .A1(w_d[266]), .A2(\w_reg/n890 ), .ZN(\w_reg/N269 )
         );
  AND2_X2 \w_reg/U326  ( .A1(w_d[267]), .A2(\w_reg/n890 ), .ZN(\w_reg/N270 )
         );
  AND2_X2 \w_reg/U325  ( .A1(w_d[268]), .A2(\w_reg/n890 ), .ZN(\w_reg/N271 )
         );
  AND2_X2 \w_reg/U324  ( .A1(w_d[269]), .A2(\w_reg/n890 ), .ZN(\w_reg/N272 )
         );
  AND2_X2 \w_reg/U323  ( .A1(w_d[270]), .A2(\w_reg/n890 ), .ZN(\w_reg/N273 )
         );
  AND2_X2 \w_reg/U322  ( .A1(w_d[271]), .A2(\w_reg/n890 ), .ZN(\w_reg/N274 )
         );
  AND2_X2 \w_reg/U321  ( .A1(w_d[272]), .A2(\w_reg/n880 ), .ZN(\w_reg/N275 )
         );
  AND2_X2 \w_reg/U320  ( .A1(w_d[273]), .A2(\w_reg/n880 ), .ZN(\w_reg/N276 )
         );
  AND2_X2 \w_reg/U319  ( .A1(w_d[274]), .A2(\w_reg/n880 ), .ZN(\w_reg/N277 )
         );
  AND2_X2 \w_reg/U318  ( .A1(w_d[275]), .A2(\w_reg/n880 ), .ZN(\w_reg/N278 )
         );
  AND2_X2 \w_reg/U317  ( .A1(w_d[276]), .A2(\w_reg/n880 ), .ZN(\w_reg/N279 )
         );
  AND2_X2 \w_reg/U315  ( .A1(w_d[277]), .A2(\w_reg/n880 ), .ZN(\w_reg/N280 )
         );
  AND2_X2 \w_reg/U314  ( .A1(w_d[278]), .A2(\w_reg/n880 ), .ZN(\w_reg/N281 )
         );
  AND2_X2 \w_reg/U313  ( .A1(w_d[279]), .A2(\w_reg/n880 ), .ZN(\w_reg/N282 )
         );
  AND2_X2 \w_reg/U312  ( .A1(w_d[280]), .A2(\w_reg/n880 ), .ZN(\w_reg/N283 )
         );
  AND2_X2 \w_reg/U311  ( .A1(w_d[281]), .A2(\w_reg/n880 ), .ZN(\w_reg/N284 )
         );
  AND2_X2 \w_reg/U310  ( .A1(w_d[282]), .A2(\w_reg/n870 ), .ZN(\w_reg/N285 )
         );
  AND2_X2 \w_reg/U309  ( .A1(w_d[283]), .A2(\w_reg/n870 ), .ZN(\w_reg/N286 )
         );
  AND2_X2 \w_reg/U308  ( .A1(w_d[284]), .A2(\w_reg/n870 ), .ZN(\w_reg/N287 )
         );
  AND2_X2 \w_reg/U307  ( .A1(w_d[285]), .A2(\w_reg/n870 ), .ZN(\w_reg/N288 )
         );
  AND2_X2 \w_reg/U306  ( .A1(w_d[286]), .A2(\w_reg/n870 ), .ZN(\w_reg/N289 )
         );
  AND2_X2 \w_reg/U304  ( .A1(w_d[287]), .A2(\w_reg/n870 ), .ZN(\w_reg/N290 )
         );
  AND2_X2 \w_reg/U303  ( .A1(w_d[288]), .A2(\w_reg/n870 ), .ZN(\w_reg/N291 )
         );
  AND2_X2 \w_reg/U302  ( .A1(w_d[289]), .A2(\w_reg/n870 ), .ZN(\w_reg/N292 )
         );
  AND2_X2 \w_reg/U301  ( .A1(w_d[290]), .A2(\w_reg/n870 ), .ZN(\w_reg/N293 )
         );
  AND2_X2 \w_reg/U300  ( .A1(w_d[291]), .A2(\w_reg/n870 ), .ZN(\w_reg/N294 )
         );
  AND2_X2 \w_reg/U299  ( .A1(w_d[292]), .A2(\w_reg/n860 ), .ZN(\w_reg/N295 )
         );
  AND2_X2 \w_reg/U298  ( .A1(w_d[293]), .A2(\w_reg/n860 ), .ZN(\w_reg/N296 )
         );
  AND2_X2 \w_reg/U297  ( .A1(w_d[294]), .A2(\w_reg/n860 ), .ZN(\w_reg/N297 )
         );
  AND2_X2 \w_reg/U296  ( .A1(w_d[295]), .A2(\w_reg/n860 ), .ZN(\w_reg/N298 )
         );
  AND2_X2 \w_reg/U295  ( .A1(w_d[296]), .A2(\w_reg/n860 ), .ZN(\w_reg/N299 )
         );
  AND2_X2 \w_reg/U292  ( .A1(w_d[297]), .A2(\w_reg/n860 ), .ZN(\w_reg/N300 )
         );
  AND2_X2 \w_reg/U291  ( .A1(w_d[298]), .A2(\w_reg/n860 ), .ZN(\w_reg/N301 )
         );
  AND2_X2 \w_reg/U290  ( .A1(w_d[299]), .A2(\w_reg/n860 ), .ZN(\w_reg/N302 )
         );
  AND2_X2 \w_reg/U289  ( .A1(w_d[300]), .A2(\w_reg/n860 ), .ZN(\w_reg/N303 )
         );
  AND2_X2 \w_reg/U288  ( .A1(w_d[301]), .A2(\w_reg/n850 ), .ZN(\w_reg/N304 )
         );
  AND2_X2 \w_reg/U287  ( .A1(w_d[302]), .A2(\w_reg/n850 ), .ZN(\w_reg/N305 )
         );
  AND2_X2 \w_reg/U286  ( .A1(w_d[303]), .A2(\w_reg/n850 ), .ZN(\w_reg/N306 )
         );
  AND2_X2 \w_reg/U285  ( .A1(w_d[304]), .A2(\w_reg/n850 ), .ZN(\w_reg/N307 )
         );
  AND2_X2 \w_reg/U284  ( .A1(w_d[305]), .A2(\w_reg/n850 ), .ZN(\w_reg/N308 )
         );
  AND2_X2 \w_reg/U283  ( .A1(w_d[306]), .A2(\w_reg/n850 ), .ZN(\w_reg/N309 )
         );
  AND2_X2 \w_reg/U281  ( .A1(w_d[307]), .A2(\w_reg/n850 ), .ZN(\w_reg/N310 )
         );
  AND2_X2 \w_reg/U280  ( .A1(w_d[308]), .A2(\w_reg/n850 ), .ZN(\w_reg/N311 )
         );
  AND2_X2 \w_reg/U279  ( .A1(w_d[309]), .A2(\w_reg/n850 ), .ZN(\w_reg/N312 )
         );
  AND2_X2 \w_reg/U278  ( .A1(w_d[310]), .A2(\w_reg/n850 ), .ZN(\w_reg/N313 )
         );
  AND2_X2 \w_reg/U277  ( .A1(w_d[311]), .A2(\w_reg/n840 ), .ZN(\w_reg/N314 )
         );
  AND2_X2 \w_reg/U276  ( .A1(w_d[312]), .A2(\w_reg/n840 ), .ZN(\w_reg/N315 )
         );
  AND2_X2 \w_reg/U275  ( .A1(w_d[313]), .A2(\w_reg/n840 ), .ZN(\w_reg/N316 )
         );
  AND2_X2 \w_reg/U274  ( .A1(w_d[314]), .A2(\w_reg/n840 ), .ZN(\w_reg/N317 )
         );
  AND2_X2 \w_reg/U273  ( .A1(w_d[315]), .A2(\w_reg/n840 ), .ZN(\w_reg/N318 )
         );
  AND2_X2 \w_reg/U272  ( .A1(w_d[316]), .A2(\w_reg/n840 ), .ZN(\w_reg/N319 )
         );
  AND2_X2 \w_reg/U270  ( .A1(w_d[317]), .A2(\w_reg/n840 ), .ZN(\w_reg/N320 )
         );
  AND2_X2 \w_reg/U269  ( .A1(w_d[318]), .A2(\w_reg/n840 ), .ZN(\w_reg/N321 )
         );
  AND2_X2 \w_reg/U268  ( .A1(w_d[319]), .A2(\w_reg/n840 ), .ZN(\w_reg/N322 )
         );
  AND2_X2 \w_reg/U267  ( .A1(w_d[320]), .A2(\w_reg/n840 ), .ZN(\w_reg/N323 )
         );
  AND2_X2 \w_reg/U266  ( .A1(w_d[321]), .A2(\w_reg/n830 ), .ZN(\w_reg/N324 )
         );
  AND2_X2 \w_reg/U265  ( .A1(w_d[322]), .A2(\w_reg/n830 ), .ZN(\w_reg/N325 )
         );
  AND2_X2 \w_reg/U264  ( .A1(w_d[323]), .A2(\w_reg/n830 ), .ZN(\w_reg/N326 )
         );
  AND2_X2 \w_reg/U263  ( .A1(w_d[324]), .A2(\w_reg/n830 ), .ZN(\w_reg/N327 )
         );
  AND2_X2 \w_reg/U262  ( .A1(w_d[325]), .A2(\w_reg/n830 ), .ZN(\w_reg/N328 )
         );
  AND2_X2 \w_reg/U261  ( .A1(w_d[326]), .A2(\w_reg/n830 ), .ZN(\w_reg/N329 )
         );
  AND2_X2 \w_reg/U259  ( .A1(w_d[327]), .A2(\w_reg/n830 ), .ZN(\w_reg/N330 )
         );
  AND2_X2 \w_reg/U258  ( .A1(w_d[328]), .A2(\w_reg/n830 ), .ZN(\w_reg/N331 )
         );
  AND2_X2 \w_reg/U257  ( .A1(w_d[329]), .A2(\w_reg/n830 ), .ZN(\w_reg/N332 )
         );
  AND2_X2 \w_reg/U256  ( .A1(w_d[330]), .A2(\w_reg/n830 ), .ZN(\w_reg/N333 )
         );
  AND2_X2 \w_reg/U255  ( .A1(w_d[331]), .A2(\w_reg/n820 ), .ZN(\w_reg/N334 )
         );
  AND2_X2 \w_reg/U254  ( .A1(w_d[332]), .A2(\w_reg/n820 ), .ZN(\w_reg/N335 )
         );
  AND2_X2 \w_reg/U253  ( .A1(w_d[333]), .A2(\w_reg/n820 ), .ZN(\w_reg/N336 )
         );
  AND2_X2 \w_reg/U252  ( .A1(w_d[334]), .A2(\w_reg/n820 ), .ZN(\w_reg/N337 )
         );
  AND2_X2 \w_reg/U251  ( .A1(w_d[335]), .A2(\w_reg/n820 ), .ZN(\w_reg/N338 )
         );
  AND2_X2 \w_reg/U250  ( .A1(w_d[336]), .A2(\w_reg/n820 ), .ZN(\w_reg/N339 )
         );
  AND2_X2 \w_reg/U248  ( .A1(w_d[337]), .A2(\w_reg/n820 ), .ZN(\w_reg/N340 )
         );
  AND2_X2 \w_reg/U247  ( .A1(w_d[338]), .A2(\w_reg/n820 ), .ZN(\w_reg/N341 )
         );
  AND2_X2 \w_reg/U246  ( .A1(w_d[339]), .A2(\w_reg/n820 ), .ZN(\w_reg/N342 )
         );
  AND2_X2 \w_reg/U245  ( .A1(w_d[340]), .A2(\w_reg/n820 ), .ZN(\w_reg/N343 )
         );
  AND2_X2 \w_reg/U244  ( .A1(w_d[341]), .A2(\w_reg/n810 ), .ZN(\w_reg/N344 )
         );
  AND2_X2 \w_reg/U243  ( .A1(w_d[342]), .A2(\w_reg/n810 ), .ZN(\w_reg/N345 )
         );
  AND2_X2 \w_reg/U242  ( .A1(w_d[343]), .A2(\w_reg/n810 ), .ZN(\w_reg/N346 )
         );
  AND2_X2 \w_reg/U241  ( .A1(w_d[344]), .A2(\w_reg/n810 ), .ZN(\w_reg/N347 )
         );
  AND2_X2 \w_reg/U240  ( .A1(w_d[345]), .A2(\w_reg/n810 ), .ZN(\w_reg/N348 )
         );
  AND2_X2 \w_reg/U239  ( .A1(w_d[346]), .A2(\w_reg/n810 ), .ZN(\w_reg/N349 )
         );
  AND2_X2 \w_reg/U238  ( .A1(w_d[32]), .A2(\w_reg/n810 ), .ZN(\w_reg/N35 ) );
  AND2_X2 \w_reg/U237  ( .A1(w_d[347]), .A2(\w_reg/n810 ), .ZN(\w_reg/N350 )
         );
  AND2_X2 \w_reg/U236  ( .A1(w_d[348]), .A2(\w_reg/n810 ), .ZN(\w_reg/N351 )
         );
  AND2_X2 \w_reg/U235  ( .A1(w_d[349]), .A2(\w_reg/n810 ), .ZN(\w_reg/N352 )
         );
  AND2_X2 \w_reg/U234  ( .A1(w_d[350]), .A2(\w_reg/n810 ), .ZN(\w_reg/N353 )
         );
  AND2_X2 \w_reg/U233  ( .A1(w_d[351]), .A2(\w_reg/n800 ), .ZN(\w_reg/N354 )
         );
  AND2_X2 \w_reg/U232  ( .A1(w_d[352]), .A2(\w_reg/n800 ), .ZN(\w_reg/N355 )
         );
  AND2_X2 \w_reg/U231  ( .A1(w_d[353]), .A2(\w_reg/n800 ), .ZN(\w_reg/N356 )
         );
  AND2_X2 \w_reg/U230  ( .A1(w_d[354]), .A2(\w_reg/n800 ), .ZN(\w_reg/N357 )
         );
  AND2_X2 \w_reg/U229  ( .A1(w_d[355]), .A2(\w_reg/n800 ), .ZN(\w_reg/N358 )
         );
  AND2_X2 \w_reg/U228  ( .A1(w_d[356]), .A2(\w_reg/n800 ), .ZN(\w_reg/N359 )
         );
  AND2_X2 \w_reg/U227  ( .A1(w_d[33]), .A2(\w_reg/n800 ), .ZN(\w_reg/N36 ) );
  AND2_X2 \w_reg/U226  ( .A1(w_d[357]), .A2(\w_reg/n800 ), .ZN(\w_reg/N360 )
         );
  AND2_X2 \w_reg/U225  ( .A1(w_d[358]), .A2(\w_reg/n800 ), .ZN(\w_reg/N361 )
         );
  AND2_X2 \w_reg/U224  ( .A1(w_d[359]), .A2(\w_reg/n800 ), .ZN(\w_reg/N362 )
         );
  AND2_X2 \w_reg/U223  ( .A1(w_d[360]), .A2(\w_reg/n800 ), .ZN(\w_reg/N363 )
         );
  AND2_X2 \w_reg/U222  ( .A1(w_d[361]), .A2(\w_reg/n790 ), .ZN(\w_reg/N364 )
         );
  AND2_X2 \w_reg/U221  ( .A1(w_d[362]), .A2(\w_reg/n790 ), .ZN(\w_reg/N365 )
         );
  AND2_X2 \w_reg/U220  ( .A1(w_d[363]), .A2(\w_reg/n790 ), .ZN(\w_reg/N366 )
         );
  AND2_X2 \w_reg/U219  ( .A1(w_d[364]), .A2(\w_reg/n790 ), .ZN(\w_reg/N367 )
         );
  AND2_X2 \w_reg/U218  ( .A1(w_d[365]), .A2(\w_reg/n790 ), .ZN(\w_reg/N368 )
         );
  AND2_X2 \w_reg/U217  ( .A1(w_d[366]), .A2(\w_reg/n790 ), .ZN(\w_reg/N369 )
         );
  AND2_X2 \w_reg/U216  ( .A1(w_d[34]), .A2(\w_reg/n790 ), .ZN(\w_reg/N37 ) );
  AND2_X2 \w_reg/U215  ( .A1(w_d[367]), .A2(\w_reg/n790 ), .ZN(\w_reg/N370 )
         );
  AND2_X2 \w_reg/U214  ( .A1(w_d[368]), .A2(\w_reg/n790 ), .ZN(\w_reg/N371 )
         );
  AND2_X2 \w_reg/U213  ( .A1(w_d[369]), .A2(\w_reg/n790 ), .ZN(\w_reg/N372 )
         );
  AND2_X2 \w_reg/U212  ( .A1(w_d[370]), .A2(\w_reg/n790 ), .ZN(\w_reg/N373 )
         );
  AND2_X2 \w_reg/U211  ( .A1(w_d[371]), .A2(\w_reg/n780 ), .ZN(\w_reg/N374 )
         );
  AND2_X2 \w_reg/U210  ( .A1(w_d[372]), .A2(\w_reg/n780 ), .ZN(\w_reg/N375 )
         );
  AND2_X2 \w_reg/U209  ( .A1(w_d[373]), .A2(\w_reg/n780 ), .ZN(\w_reg/N376 )
         );
  AND2_X2 \w_reg/U208  ( .A1(w_d[374]), .A2(\w_reg/n780 ), .ZN(\w_reg/N377 )
         );
  AND2_X2 \w_reg/U207  ( .A1(w_d[375]), .A2(\w_reg/n780 ), .ZN(\w_reg/N378 )
         );
  AND2_X2 \w_reg/U206  ( .A1(w_d[376]), .A2(\w_reg/n780 ), .ZN(\w_reg/N379 )
         );
  AND2_X2 \w_reg/U205  ( .A1(w_d[35]), .A2(\w_reg/n780 ), .ZN(\w_reg/N38 ) );
  AND2_X2 \w_reg/U204  ( .A1(w_d[377]), .A2(\w_reg/n780 ), .ZN(\w_reg/N380 )
         );
  AND2_X2 \w_reg/U203  ( .A1(w_d[378]), .A2(\w_reg/n780 ), .ZN(\w_reg/N381 )
         );
  AND2_X2 \w_reg/U202  ( .A1(w_d[379]), .A2(\w_reg/n780 ), .ZN(\w_reg/N382 )
         );
  AND2_X2 \w_reg/U201  ( .A1(w_d[380]), .A2(\w_reg/n780 ), .ZN(\w_reg/N383 )
         );
  AND2_X2 \w_reg/U200  ( .A1(w_d[381]), .A2(\w_reg/n770 ), .ZN(\w_reg/N384 )
         );
  AND2_X2 \w_reg/U199  ( .A1(w_d[382]), .A2(\w_reg/n770 ), .ZN(\w_reg/N385 )
         );
  AND2_X2 \w_reg/U198  ( .A1(w_d[383]), .A2(\w_reg/n770 ), .ZN(\w_reg/N386 )
         );
  AND2_X2 \w_reg/U197  ( .A1(w_d[384]), .A2(\w_reg/n770 ), .ZN(\w_reg/N387 )
         );
  AND2_X2 \w_reg/U196  ( .A1(w_d[385]), .A2(\w_reg/n770 ), .ZN(\w_reg/N388 )
         );
  AND2_X2 \w_reg/U195  ( .A1(w_d[386]), .A2(\w_reg/n770 ), .ZN(\w_reg/N389 )
         );
  AND2_X2 \w_reg/U194  ( .A1(w_d[36]), .A2(\w_reg/n770 ), .ZN(\w_reg/N39 ) );
  AND2_X2 \w_reg/U193  ( .A1(w_d[387]), .A2(\w_reg/n770 ), .ZN(\w_reg/N390 )
         );
  AND2_X2 \w_reg/U192  ( .A1(w_d[388]), .A2(\w_reg/n770 ), .ZN(\w_reg/N391 )
         );
  AND2_X2 \w_reg/U191  ( .A1(w_d[389]), .A2(\w_reg/n770 ), .ZN(\w_reg/N392 )
         );
  AND2_X2 \w_reg/U190  ( .A1(w_d[390]), .A2(\w_reg/n770 ), .ZN(\w_reg/N393 )
         );
  AND2_X2 \w_reg/U189  ( .A1(w_d[391]), .A2(\w_reg/n760 ), .ZN(\w_reg/N394 )
         );
  AND2_X2 \w_reg/U188  ( .A1(w_d[392]), .A2(\w_reg/n760 ), .ZN(\w_reg/N395 )
         );
  AND2_X2 \w_reg/U187  ( .A1(w_d[393]), .A2(\w_reg/n760 ), .ZN(\w_reg/N396 )
         );
  AND2_X2 \w_reg/U186  ( .A1(w_d[394]), .A2(\w_reg/n760 ), .ZN(\w_reg/N397 )
         );
  AND2_X2 \w_reg/U185  ( .A1(w_d[395]), .A2(\w_reg/n760 ), .ZN(\w_reg/N398 )
         );
  AND2_X2 \w_reg/U184  ( .A1(w_d[396]), .A2(\w_reg/n760 ), .ZN(\w_reg/N399 )
         );
  AND2_X2 \w_reg/U182  ( .A1(w_d[37]), .A2(\w_reg/n760 ), .ZN(\w_reg/N40 ) );
  AND2_X2 \w_reg/U181  ( .A1(w_d[397]), .A2(\w_reg/n760 ), .ZN(\w_reg/N400 )
         );
  AND2_X2 \w_reg/U180  ( .A1(w_d[398]), .A2(\w_reg/n760 ), .ZN(\w_reg/N401 )
         );
  AND2_X2 \w_reg/U179  ( .A1(w_d[399]), .A2(\w_reg/n760 ), .ZN(\w_reg/N402 )
         );
  AND2_X2 \w_reg/U178  ( .A1(w_d[400]), .A2(\w_reg/n750 ), .ZN(\w_reg/N403 )
         );
  AND2_X2 \w_reg/U177  ( .A1(w_d[401]), .A2(\w_reg/n750 ), .ZN(\w_reg/N404 )
         );
  AND2_X2 \w_reg/U176  ( .A1(w_d[402]), .A2(\w_reg/n750 ), .ZN(\w_reg/N405 )
         );
  AND2_X2 \w_reg/U175  ( .A1(w_d[403]), .A2(\w_reg/n750 ), .ZN(\w_reg/N406 )
         );
  AND2_X2 \w_reg/U174  ( .A1(w_d[404]), .A2(\w_reg/n750 ), .ZN(\w_reg/N407 )
         );
  AND2_X2 \w_reg/U173  ( .A1(w_d[405]), .A2(\w_reg/n750 ), .ZN(\w_reg/N408 )
         );
  AND2_X2 \w_reg/U172  ( .A1(w_d[406]), .A2(\w_reg/n750 ), .ZN(\w_reg/N409 )
         );
  AND2_X2 \w_reg/U171  ( .A1(w_d[38]), .A2(\w_reg/n750 ), .ZN(\w_reg/N41 ) );
  AND2_X2 \w_reg/U170  ( .A1(w_d[407]), .A2(\w_reg/n750 ), .ZN(\w_reg/N410 )
         );
  AND2_X2 \w_reg/U169  ( .A1(w_d[408]), .A2(\w_reg/n750 ), .ZN(\w_reg/N411 )
         );
  AND2_X2 \w_reg/U168  ( .A1(w_d[409]), .A2(\w_reg/n750 ), .ZN(\w_reg/N412 )
         );
  AND2_X2 \w_reg/U167  ( .A1(w_d[410]), .A2(\w_reg/n740 ), .ZN(\w_reg/N413 )
         );
  AND2_X2 \w_reg/U166  ( .A1(w_d[411]), .A2(\w_reg/n740 ), .ZN(\w_reg/N414 )
         );
  AND2_X2 \w_reg/U165  ( .A1(w_d[412]), .A2(\w_reg/n740 ), .ZN(\w_reg/N415 )
         );
  AND2_X2 \w_reg/U164  ( .A1(w_d[413]), .A2(\w_reg/n740 ), .ZN(\w_reg/N416 )
         );
  AND2_X2 \w_reg/U163  ( .A1(w_d[414]), .A2(\w_reg/n740 ), .ZN(\w_reg/N417 )
         );
  AND2_X2 \w_reg/U162  ( .A1(w_d[415]), .A2(\w_reg/n740 ), .ZN(\w_reg/N418 )
         );
  AND2_X2 \w_reg/U161  ( .A1(w_d[416]), .A2(\w_reg/n740 ), .ZN(\w_reg/N419 )
         );
  AND2_X2 \w_reg/U160  ( .A1(w_d[39]), .A2(\w_reg/n740 ), .ZN(\w_reg/N42 ) );
  AND2_X2 \w_reg/U159  ( .A1(w_d[417]), .A2(\w_reg/n740 ), .ZN(\w_reg/N420 )
         );
  AND2_X2 \w_reg/U158  ( .A1(w_d[418]), .A2(\w_reg/n740 ), .ZN(\w_reg/N421 )
         );
  AND2_X2 \w_reg/U157  ( .A1(w_d[419]), .A2(\w_reg/n740 ), .ZN(\w_reg/N422 )
         );
  AND2_X2 \w_reg/U156  ( .A1(w_d[420]), .A2(\w_reg/n730 ), .ZN(\w_reg/N423 )
         );
  AND2_X2 \w_reg/U155  ( .A1(w_d[421]), .A2(\w_reg/n730 ), .ZN(\w_reg/N424 )
         );
  AND2_X2 \w_reg/U154  ( .A1(w_d[422]), .A2(\w_reg/n730 ), .ZN(\w_reg/N425 )
         );
  AND2_X2 \w_reg/U153  ( .A1(w_d[423]), .A2(\w_reg/n730 ), .ZN(\w_reg/N426 )
         );
  AND2_X2 \w_reg/U152  ( .A1(w_d[424]), .A2(\w_reg/n730 ), .ZN(\w_reg/N427 )
         );
  AND2_X2 \w_reg/U151  ( .A1(w_d[425]), .A2(\w_reg/n730 ), .ZN(\w_reg/N428 )
         );
  AND2_X2 \w_reg/U150  ( .A1(w_d[426]), .A2(\w_reg/n730 ), .ZN(\w_reg/N429 )
         );
  AND2_X2 \w_reg/U149  ( .A1(w_d[40]), .A2(\w_reg/n730 ), .ZN(\w_reg/N43 ) );
  AND2_X2 \w_reg/U148  ( .A1(w_d[427]), .A2(\w_reg/n730 ), .ZN(\w_reg/N430 )
         );
  AND2_X2 \w_reg/U147  ( .A1(w_d[428]), .A2(\w_reg/n730 ), .ZN(\w_reg/N431 )
         );
  AND2_X2 \w_reg/U146  ( .A1(w_d[429]), .A2(\w_reg/n730 ), .ZN(\w_reg/N432 )
         );
  AND2_X2 \w_reg/U145  ( .A1(w_d[430]), .A2(\w_reg/n720 ), .ZN(\w_reg/N433 )
         );
  AND2_X2 \w_reg/U144  ( .A1(w_d[431]), .A2(\w_reg/n720 ), .ZN(\w_reg/N434 )
         );
  AND2_X2 \w_reg/U143  ( .A1(w_d[432]), .A2(\w_reg/n720 ), .ZN(\w_reg/N435 )
         );
  AND2_X2 \w_reg/U142  ( .A1(w_d[433]), .A2(\w_reg/n720 ), .ZN(\w_reg/N436 )
         );
  AND2_X2 \w_reg/U141  ( .A1(w_d[434]), .A2(\w_reg/n720 ), .ZN(\w_reg/N437 )
         );
  AND2_X2 \w_reg/U140  ( .A1(w_d[435]), .A2(\w_reg/n720 ), .ZN(\w_reg/N438 )
         );
  AND2_X2 \w_reg/U139  ( .A1(w_d[436]), .A2(\w_reg/n720 ), .ZN(\w_reg/N439 )
         );
  AND2_X2 \w_reg/U138  ( .A1(w_d[41]), .A2(\w_reg/n720 ), .ZN(\w_reg/N44 ) );
  AND2_X2 \w_reg/U137  ( .A1(w_d[437]), .A2(\w_reg/n720 ), .ZN(\w_reg/N440 )
         );
  AND2_X2 \w_reg/U136  ( .A1(w_d[438]), .A2(\w_reg/n720 ), .ZN(\w_reg/N441 )
         );
  AND2_X2 \w_reg/U135  ( .A1(w_d[439]), .A2(\w_reg/n720 ), .ZN(\w_reg/N442 )
         );
  AND2_X2 \w_reg/U134  ( .A1(w_d[440]), .A2(\w_reg/n710 ), .ZN(\w_reg/N443 )
         );
  AND2_X2 \w_reg/U133  ( .A1(w_d[441]), .A2(\w_reg/n710 ), .ZN(\w_reg/N444 )
         );
  AND2_X2 \w_reg/U132  ( .A1(w_d[442]), .A2(\w_reg/n710 ), .ZN(\w_reg/N445 )
         );
  AND2_X2 \w_reg/U131  ( .A1(w_d[443]), .A2(\w_reg/n710 ), .ZN(\w_reg/N446 )
         );
  AND2_X2 \w_reg/U130  ( .A1(w_d[444]), .A2(\w_reg/n710 ), .ZN(\w_reg/N447 )
         );
  AND2_X2 \w_reg/U129  ( .A1(w_d[445]), .A2(\w_reg/n710 ), .ZN(\w_reg/N448 )
         );
  AND2_X2 \w_reg/U128  ( .A1(w_d[446]), .A2(\w_reg/n710 ), .ZN(\w_reg/N449 )
         );
  AND2_X2 \w_reg/U127  ( .A1(w_d[42]), .A2(\w_reg/n710 ), .ZN(\w_reg/N45 ) );
  AND2_X2 \w_reg/U126  ( .A1(w_d[447]), .A2(\w_reg/n710 ), .ZN(\w_reg/N450 )
         );
  AND2_X2 \w_reg/U125  ( .A1(w_d[448]), .A2(\w_reg/n710 ), .ZN(\w_reg/N451 )
         );
  AND2_X2 \w_reg/U124  ( .A1(w_d[449]), .A2(\w_reg/n710 ), .ZN(\w_reg/N452 )
         );
  AND2_X2 \w_reg/U123  ( .A1(w_d[450]), .A2(\w_reg/n700 ), .ZN(\w_reg/N453 )
         );
  AND2_X2 \w_reg/U122  ( .A1(w_d[451]), .A2(\w_reg/n700 ), .ZN(\w_reg/N454 )
         );
  AND2_X2 \w_reg/U121  ( .A1(w_d[452]), .A2(\w_reg/n700 ), .ZN(\w_reg/N455 )
         );
  AND2_X2 \w_reg/U120  ( .A1(w_d[453]), .A2(\w_reg/n700 ), .ZN(\w_reg/N456 )
         );
  AND2_X2 \w_reg/U119  ( .A1(w_d[454]), .A2(\w_reg/n700 ), .ZN(\w_reg/N457 )
         );
  AND2_X2 \w_reg/U118  ( .A1(w_d[455]), .A2(\w_reg/n700 ), .ZN(\w_reg/N458 )
         );
  AND2_X2 \w_reg/U117  ( .A1(w_d[456]), .A2(\w_reg/n700 ), .ZN(\w_reg/N459 )
         );
  AND2_X2 \w_reg/U116  ( .A1(w_d[43]), .A2(\w_reg/n700 ), .ZN(\w_reg/N46 ) );
  AND2_X2 \w_reg/U115  ( .A1(w_d[457]), .A2(\w_reg/n700 ), .ZN(\w_reg/N460 )
         );
  AND2_X2 \w_reg/U114  ( .A1(w_d[458]), .A2(\w_reg/n700 ), .ZN(\w_reg/N461 )
         );
  AND2_X2 \w_reg/U113  ( .A1(w_d[459]), .A2(\w_reg/n700 ), .ZN(\w_reg/N462 )
         );
  AND2_X2 \w_reg/U112  ( .A1(w_d[460]), .A2(\w_reg/n690 ), .ZN(\w_reg/N463 )
         );
  AND2_X2 \w_reg/U111  ( .A1(w_d[461]), .A2(\w_reg/n690 ), .ZN(\w_reg/N464 )
         );
  AND2_X2 \w_reg/U110  ( .A1(w_d[462]), .A2(\w_reg/n690 ), .ZN(\w_reg/N465 )
         );
  AND2_X2 \w_reg/U109  ( .A1(w_d[463]), .A2(\w_reg/n690 ), .ZN(\w_reg/N466 )
         );
  AND2_X2 \w_reg/U108  ( .A1(w_d[464]), .A2(\w_reg/n690 ), .ZN(\w_reg/N467 )
         );
  AND2_X2 \w_reg/U107  ( .A1(w_d[465]), .A2(\w_reg/n690 ), .ZN(\w_reg/N468 )
         );
  AND2_X2 \w_reg/U106  ( .A1(w_d[466]), .A2(\w_reg/n690 ), .ZN(\w_reg/N469 )
         );
  AND2_X2 \w_reg/U105  ( .A1(w_d[44]), .A2(\w_reg/n690 ), .ZN(\w_reg/N47 ) );
  AND2_X2 \w_reg/U104  ( .A1(w_d[467]), .A2(\w_reg/n690 ), .ZN(\w_reg/N470 )
         );
  AND2_X2 \w_reg/U103  ( .A1(w_d[468]), .A2(\w_reg/n690 ), .ZN(\w_reg/N471 )
         );
  AND2_X2 \w_reg/U102  ( .A1(w_d[469]), .A2(\w_reg/n690 ), .ZN(\w_reg/N472 )
         );
  AND2_X2 \w_reg/U101  ( .A1(w_d[470]), .A2(\w_reg/n680 ), .ZN(\w_reg/N473 )
         );
  AND2_X2 \w_reg/U100  ( .A1(w_d[471]), .A2(\w_reg/n680 ), .ZN(\w_reg/N474 )
         );
  AND2_X2 \w_reg/U99  ( .A1(w_d[472]), .A2(\w_reg/n680 ), .ZN(\w_reg/N475 ) );
  AND2_X2 \w_reg/U98  ( .A1(w_d[473]), .A2(\w_reg/n680 ), .ZN(\w_reg/N476 ) );
  AND2_X2 \w_reg/U97  ( .A1(w_d[474]), .A2(\w_reg/n680 ), .ZN(\w_reg/N477 ) );
  AND2_X2 \w_reg/U96  ( .A1(w_d[475]), .A2(\w_reg/n680 ), .ZN(\w_reg/N478 ) );
  AND2_X2 \w_reg/U95  ( .A1(w_d[476]), .A2(\w_reg/n680 ), .ZN(\w_reg/N479 ) );
  AND2_X2 \w_reg/U94  ( .A1(w_d[45]), .A2(\w_reg/n680 ), .ZN(\w_reg/N48 ) );
  AND2_X2 \w_reg/U93  ( .A1(w_d[477]), .A2(\w_reg/n680 ), .ZN(\w_reg/N480 ) );
  AND2_X2 \w_reg/U92  ( .A1(w_d[478]), .A2(\w_reg/n680 ), .ZN(\w_reg/N481 ) );
  AND2_X2 \w_reg/U91  ( .A1(w_d[479]), .A2(\w_reg/n680 ), .ZN(\w_reg/N482 ) );
  AND2_X2 \w_reg/U83  ( .A1(w_d[46]), .A2(\w_reg/n670 ), .ZN(\w_reg/N49 ) );
  AND2_X2 \w_reg/U71  ( .A1(w_d[47]), .A2(\w_reg/n670 ), .ZN(\w_reg/N50 ) );
  AND2_X2 \w_reg/U69  ( .A1(w_d[498]), .A2(\w_reg/n670 ), .ZN(\w_reg/N501 ) );
  AND2_X2 \w_reg/U68  ( .A1(w_d[499]), .A2(\w_reg/n670 ), .ZN(\w_reg/N502 ) );
  AND2_X2 \w_reg/U67  ( .A1(w_d[500]), .A2(\w_reg/n670 ), .ZN(\w_reg/N503 ) );
  AND2_X2 \w_reg/U66  ( .A1(w_d[501]), .A2(\w_reg/n670 ), .ZN(\w_reg/N504 ) );
  AND2_X2 \w_reg/U65  ( .A1(w_d[502]), .A2(\w_reg/n670 ), .ZN(\w_reg/N505 ) );
  AND2_X2 \w_reg/U64  ( .A1(w_d[503]), .A2(\w_reg/n670 ), .ZN(\w_reg/N506 ) );
  AND2_X2 \w_reg/U63  ( .A1(w_d[504]), .A2(\w_reg/n670 ), .ZN(\w_reg/N507 ) );
  AND2_X2 \w_reg/U62  ( .A1(w_d[505]), .A2(\w_reg/n670 ), .ZN(\w_reg/N508 ) );
  AND2_X2 \w_reg/U61  ( .A1(w_d[506]), .A2(\w_reg/n660 ), .ZN(\w_reg/N509 ) );
  AND2_X2 \w_reg/U60  ( .A1(w_d[48]), .A2(\w_reg/n660 ), .ZN(\w_reg/N51 ) );
  AND2_X2 \w_reg/U59  ( .A1(w_d[507]), .A2(\w_reg/n660 ), .ZN(\w_reg/N510 ) );
  AND2_X2 \w_reg/U58  ( .A1(w_d[508]), .A2(\w_reg/n660 ), .ZN(\w_reg/N511 ) );
  AND2_X2 \w_reg/U57  ( .A1(w_d[509]), .A2(\w_reg/n660 ), .ZN(\w_reg/N512 ) );
  AND2_X2 \w_reg/U56  ( .A1(w_d[510]), .A2(\w_reg/n660 ), .ZN(\w_reg/N513 ) );
  AND2_X2 \w_reg/U55  ( .A1(w_d[511]), .A2(\w_reg/n660 ), .ZN(\w_reg/N514 ) );
  AND2_X2 \w_reg/U54  ( .A1(w_d[49]), .A2(\w_reg/n660 ), .ZN(\w_reg/N52 ) );
  AND2_X2 \w_reg/U53  ( .A1(w_d[50]), .A2(\w_reg/n660 ), .ZN(\w_reg/N53 ) );
  AND2_X2 \w_reg/U52  ( .A1(w_d[51]), .A2(\w_reg/n660 ), .ZN(\w_reg/N54 ) );
  AND2_X2 \w_reg/U51  ( .A1(w_d[52]), .A2(\w_reg/n660 ), .ZN(\w_reg/N55 ) );
  AND2_X2 \w_reg/U50  ( .A1(w_d[53]), .A2(\w_reg/n650 ), .ZN(\w_reg/N56 ) );
  AND2_X2 \w_reg/U49  ( .A1(w_d[54]), .A2(\w_reg/n650 ), .ZN(\w_reg/N57 ) );
  AND2_X2 \w_reg/U48  ( .A1(w_d[55]), .A2(\w_reg/n650 ), .ZN(\w_reg/N58 ) );
  AND2_X2 \w_reg/U47  ( .A1(w_d[56]), .A2(\w_reg/n650 ), .ZN(\w_reg/N59 ) );
  AND2_X2 \w_reg/U45  ( .A1(w_d[57]), .A2(\w_reg/n650 ), .ZN(\w_reg/N60 ) );
  AND2_X2 \w_reg/U44  ( .A1(w_d[58]), .A2(\w_reg/n650 ), .ZN(\w_reg/N61 ) );
  AND2_X2 \w_reg/U43  ( .A1(w_d[59]), .A2(\w_reg/n650 ), .ZN(\w_reg/N62 ) );
  AND2_X2 \w_reg/U42  ( .A1(w_d[60]), .A2(\w_reg/n650 ), .ZN(\w_reg/N63 ) );
  AND2_X2 \w_reg/U41  ( .A1(w_d[61]), .A2(\w_reg/n650 ), .ZN(\w_reg/N64 ) );
  AND2_X2 \w_reg/U40  ( .A1(w_d[62]), .A2(\w_reg/n650 ), .ZN(\w_reg/N65 ) );
  AND2_X2 \w_reg/U39  ( .A1(w_d[63]), .A2(\w_reg/n640 ), .ZN(\w_reg/N66 ) );
  AND2_X2 \w_reg/U38  ( .A1(w_d[64]), .A2(\w_reg/n640 ), .ZN(\w_reg/N67 ) );
  AND2_X2 \w_reg/U37  ( .A1(w_d[65]), .A2(\w_reg/n640 ), .ZN(\w_reg/N68 ) );
  AND2_X2 \w_reg/U36  ( .A1(w_d[66]), .A2(\w_reg/n640 ), .ZN(\w_reg/N69 ) );
  AND2_X2 \w_reg/U34  ( .A1(w_d[67]), .A2(\w_reg/n640 ), .ZN(\w_reg/N70 ) );
  AND2_X2 \w_reg/U33  ( .A1(w_d[68]), .A2(\w_reg/n640 ), .ZN(\w_reg/N71 ) );
  AND2_X2 \w_reg/U32  ( .A1(w_d[69]), .A2(\w_reg/n640 ), .ZN(\w_reg/N72 ) );
  AND2_X2 \w_reg/U31  ( .A1(w_d[70]), .A2(\w_reg/n640 ), .ZN(\w_reg/N73 ) );
  AND2_X2 \w_reg/U30  ( .A1(w_d[71]), .A2(\w_reg/n640 ), .ZN(\w_reg/N74 ) );
  AND2_X2 \w_reg/U29  ( .A1(w_d[72]), .A2(\w_reg/n640 ), .ZN(\w_reg/N75 ) );
  AND2_X2 \w_reg/U28  ( .A1(w_d[73]), .A2(\w_reg/n630 ), .ZN(\w_reg/N76 ) );
  AND2_X2 \w_reg/U27  ( .A1(w_d[74]), .A2(\w_reg/n630 ), .ZN(\w_reg/N77 ) );
  AND2_X2 \w_reg/U26  ( .A1(w_d[75]), .A2(\w_reg/n630 ), .ZN(\w_reg/N78 ) );
  AND2_X2 \w_reg/U25  ( .A1(w_d[76]), .A2(\w_reg/n630 ), .ZN(\w_reg/N79 ) );
  AND2_X2 \w_reg/U23  ( .A1(w_d[77]), .A2(\w_reg/n630 ), .ZN(\w_reg/N80 ) );
  AND2_X2 \w_reg/U22  ( .A1(w_d[78]), .A2(\w_reg/n630 ), .ZN(\w_reg/N81 ) );
  AND2_X2 \w_reg/U21  ( .A1(w_d[79]), .A2(\w_reg/n630 ), .ZN(\w_reg/N82 ) );
  AND2_X2 \w_reg/U20  ( .A1(w_d[80]), .A2(\w_reg/n630 ), .ZN(\w_reg/N83 ) );
  AND2_X2 \w_reg/U19  ( .A1(w_d[81]), .A2(\w_reg/n630 ), .ZN(\w_reg/N84 ) );
  AND2_X2 \w_reg/U18  ( .A1(w_d[82]), .A2(\w_reg/n630 ), .ZN(\w_reg/N85 ) );
  AND2_X2 \w_reg/U17  ( .A1(w_d[83]), .A2(\w_reg/n620 ), .ZN(\w_reg/N86 ) );
  AND2_X2 \w_reg/U16  ( .A1(w_d[84]), .A2(\w_reg/n620 ), .ZN(\w_reg/N87 ) );
  AND2_X2 \w_reg/U15  ( .A1(w_d[85]), .A2(\w_reg/n620 ), .ZN(\w_reg/N88 ) );
  AND2_X2 \w_reg/U14  ( .A1(w_d[86]), .A2(\w_reg/n620 ), .ZN(\w_reg/N89 ) );
  AND2_X2 \w_reg/U12  ( .A1(w_d[87]), .A2(\w_reg/n620 ), .ZN(\w_reg/N90 ) );
  AND2_X2 \w_reg/U11  ( .A1(w_d[88]), .A2(\w_reg/n620 ), .ZN(\w_reg/N91 ) );
  AND2_X2 \w_reg/U10  ( .A1(w_d[89]), .A2(\w_reg/n620 ), .ZN(\w_reg/N92 ) );
  AND2_X2 \w_reg/U9  ( .A1(w_d[90]), .A2(\w_reg/n620 ), .ZN(\w_reg/N93 ) );
  AND2_X2 \w_reg/U8  ( .A1(w_d[91]), .A2(\w_reg/n620 ), .ZN(\w_reg/N94 ) );
  AND2_X2 \w_reg/U7  ( .A1(w_d[92]), .A2(\w_reg/n620 ), .ZN(\w_reg/N95 ) );
  AND2_X2 \w_reg/U6  ( .A1(w_d[93]), .A2(\w_reg/n610 ), .ZN(\w_reg/N96 ) );
  AND2_X2 \w_reg/U5  ( .A1(w_d[94]), .A2(\w_reg/n610 ), .ZN(\w_reg/N97 ) );
  AND2_X2 \w_reg/U4  ( .A1(w_d[95]), .A2(\w_reg/n610 ), .ZN(\w_reg/N98 ) );
  AND2_X2 \w_reg/U3  ( .A1(w_d[96]), .A2(\w_reg/n610 ), .ZN(\w_reg/N99 ) );
  DFF_X2 \w_reg/q_reg_0_  ( .D(\w_reg/N3 ), .CK(clk), .Q(w_q[0]), .QN() );
  DFF_X2 \w_reg/q_reg_1_  ( .D(\w_reg/N4 ), .CK(clk), .Q(w_q[1]), .QN() );
  DFF_X2 \w_reg/q_reg_2_  ( .D(\w_reg/N5 ), .CK(clk), .Q(w_q[2]), .QN() );
  DFF_X2 \w_reg/q_reg_3_  ( .D(\w_reg/N6 ), .CK(clk), .Q(w_q[3]), .QN() );
  DFF_X2 \w_reg/q_reg_4_  ( .D(\w_reg/N7 ), .CK(clk), .Q(w_q[4]), .QN() );
  DFF_X2 \w_reg/q_reg_5_  ( .D(\w_reg/N8 ), .CK(clk), .Q(w_q[5]), .QN() );
  DFF_X2 \w_reg/q_reg_6_  ( .D(\w_reg/N9 ), .CK(clk), .Q(w_q[6]), .QN() );
  DFF_X2 \w_reg/q_reg_7_  ( .D(\w_reg/N10 ), .CK(clk), .Q(w_q[7]), .QN() );
  DFF_X2 \w_reg/q_reg_8_  ( .D(\w_reg/N11 ), .CK(clk), .Q(w_q[8]), .QN() );
  DFF_X2 \w_reg/q_reg_9_  ( .D(\w_reg/N12 ), .CK(clk), .Q(w_q[9]), .QN() );
  DFF_X2 \w_reg/q_reg_10_  ( .D(\w_reg/N13 ), .CK(clk), .Q(w_q[10]), .QN() );
  DFF_X2 \w_reg/q_reg_11_  ( .D(\w_reg/N14 ), .CK(clk), .Q(w_q[11]), .QN() );
  DFF_X2 \w_reg/q_reg_12_  ( .D(\w_reg/N15 ), .CK(clk), .Q(w_q[12]), .QN() );
  DFF_X2 \w_reg/q_reg_13_  ( .D(\w_reg/N16 ), .CK(clk), .Q(w_q[13]), .QN() );
  DFF_X2 \w_reg/q_reg_14_  ( .D(\w_reg/N17 ), .CK(clk), .Q(w_q[14]), .QN() );
  DFF_X2 \w_reg/q_reg_15_  ( .D(\w_reg/N18 ), .CK(clk), .Q(w_q[15]), .QN() );
  DFF_X2 \w_reg/q_reg_16_  ( .D(\w_reg/N19 ), .CK(clk), .Q(w_q[16]), .QN() );
  DFF_X2 \w_reg/q_reg_17_  ( .D(\w_reg/N20 ), .CK(clk), .Q(w_q[17]), .QN() );
  DFF_X2 \w_reg/q_reg_18_  ( .D(\w_reg/N21 ), .CK(clk), .Q(w_q[18]), .QN() );
  DFF_X2 \w_reg/q_reg_19_  ( .D(\w_reg/N22 ), .CK(clk), .Q(w_q[19]), .QN() );
  DFF_X2 \w_reg/q_reg_20_  ( .D(\w_reg/N23 ), .CK(clk), .Q(w_q[20]), .QN() );
  DFF_X2 \w_reg/q_reg_21_  ( .D(\w_reg/N24 ), .CK(clk), .Q(w_q[21]), .QN() );
  DFF_X2 \w_reg/q_reg_22_  ( .D(\w_reg/N25 ), .CK(clk), .Q(w_q[22]), .QN() );
  DFF_X2 \w_reg/q_reg_23_  ( .D(\w_reg/N26 ), .CK(clk), .Q(w_q[23]), .QN() );
  DFF_X2 \w_reg/q_reg_24_  ( .D(\w_reg/N27 ), .CK(clk), .Q(w_q[24]), .QN() );
  DFF_X2 \w_reg/q_reg_25_  ( .D(\w_reg/N28 ), .CK(clk), .Q(w_q[25]), .QN() );
  DFF_X2 \w_reg/q_reg_26_  ( .D(\w_reg/N29 ), .CK(clk), .Q(w_q[26]), .QN() );
  DFF_X2 \w_reg/q_reg_27_  ( .D(\w_reg/N30 ), .CK(clk), .Q(w_q[27]), .QN() );
  DFF_X2 \w_reg/q_reg_28_  ( .D(\w_reg/N31 ), .CK(clk), .Q(w_q[28]), .QN() );
  DFF_X2 \w_reg/q_reg_29_  ( .D(\w_reg/N32 ), .CK(clk), .Q(w_q[29]), .QN() );
  DFF_X2 \w_reg/q_reg_30_  ( .D(\w_reg/N33 ), .CK(clk), .Q(w_q[30]), .QN() );
  DFF_X2 \w_reg/q_reg_31_  ( .D(\w_reg/N34 ), .CK(clk), .Q(w_q[31]), .QN() );
  DFF_X2 \w_reg/q_reg_32_  ( .D(\w_reg/N35 ), .CK(clk), .Q(w_q[32]), .QN() );
  DFF_X2 \w_reg/q_reg_33_  ( .D(\w_reg/N36 ), .CK(clk), .Q(w_q[33]), .QN() );
  DFF_X2 \w_reg/q_reg_34_  ( .D(\w_reg/N37 ), .CK(clk), .Q(w_q[34]), .QN() );
  DFF_X2 \w_reg/q_reg_35_  ( .D(\w_reg/N38 ), .CK(clk), .Q(w_q[35]), .QN() );
  DFF_X2 \w_reg/q_reg_36_  ( .D(\w_reg/N39 ), .CK(clk), .Q(w_q[36]), .QN() );
  DFF_X2 \w_reg/q_reg_37_  ( .D(\w_reg/N40 ), .CK(clk), .Q(w_q[37]), .QN() );
  DFF_X2 \w_reg/q_reg_38_  ( .D(\w_reg/N41 ), .CK(clk), .Q(w_q[38]), .QN() );
  DFF_X2 \w_reg/q_reg_39_  ( .D(\w_reg/N42 ), .CK(clk), .Q(w_q[39]), .QN() );
  DFF_X2 \w_reg/q_reg_40_  ( .D(\w_reg/N43 ), .CK(clk), .Q(w_q[40]), .QN() );
  DFF_X2 \w_reg/q_reg_41_  ( .D(\w_reg/N44 ), .CK(clk), .Q(w_q[41]), .QN() );
  DFF_X2 \w_reg/q_reg_42_  ( .D(\w_reg/N45 ), .CK(clk), .Q(w_q[42]), .QN() );
  DFF_X2 \w_reg/q_reg_43_  ( .D(\w_reg/N46 ), .CK(clk), .Q(w_q[43]), .QN() );
  DFF_X2 \w_reg/q_reg_44_  ( .D(\w_reg/N47 ), .CK(clk), .Q(w_q[44]), .QN() );
  DFF_X2 \w_reg/q_reg_45_  ( .D(\w_reg/N48 ), .CK(clk), .Q(w_q[45]), .QN() );
  DFF_X2 \w_reg/q_reg_46_  ( .D(\w_reg/N49 ), .CK(clk), .Q(w_q[46]), .QN() );
  DFF_X2 \w_reg/q_reg_47_  ( .D(\w_reg/N50 ), .CK(clk), .Q(w_q[47]), .QN() );
  DFF_X2 \w_reg/q_reg_48_  ( .D(\w_reg/N51 ), .CK(clk), .Q(w_q[48]), .QN() );
  DFF_X2 \w_reg/q_reg_49_  ( .D(\w_reg/N52 ), .CK(clk), .Q(w_q[49]), .QN() );
  DFF_X2 \w_reg/q_reg_50_  ( .D(\w_reg/N53 ), .CK(clk), .Q(w_q[50]), .QN() );
  DFF_X2 \w_reg/q_reg_51_  ( .D(\w_reg/N54 ), .CK(clk), .Q(w_q[51]), .QN() );
  DFF_X2 \w_reg/q_reg_52_  ( .D(\w_reg/N55 ), .CK(clk), .Q(w_q[52]), .QN() );
  DFF_X2 \w_reg/q_reg_53_  ( .D(\w_reg/N56 ), .CK(clk), .Q(w_q[53]), .QN() );
  DFF_X2 \w_reg/q_reg_54_  ( .D(\w_reg/N57 ), .CK(clk), .Q(w_q[54]), .QN() );
  DFF_X2 \w_reg/q_reg_55_  ( .D(\w_reg/N58 ), .CK(clk), .Q(w_q[55]), .QN() );
  DFF_X2 \w_reg/q_reg_56_  ( .D(\w_reg/N59 ), .CK(clk), .Q(w_q[56]), .QN() );
  DFF_X2 \w_reg/q_reg_57_  ( .D(\w_reg/N60 ), .CK(clk), .Q(w_q[57]), .QN() );
  DFF_X2 \w_reg/q_reg_58_  ( .D(\w_reg/N61 ), .CK(clk), .Q(w_q[58]), .QN() );
  DFF_X2 \w_reg/q_reg_59_  ( .D(\w_reg/N62 ), .CK(clk), .Q(w_q[59]), .QN() );
  DFF_X2 \w_reg/q_reg_60_  ( .D(\w_reg/N63 ), .CK(clk), .Q(w_q[60]), .QN() );
  DFF_X2 \w_reg/q_reg_61_  ( .D(\w_reg/N64 ), .CK(clk), .Q(w_q[61]), .QN() );
  DFF_X2 \w_reg/q_reg_62_  ( .D(\w_reg/N65 ), .CK(clk), .Q(w_q[62]), .QN() );
  DFF_X2 \w_reg/q_reg_63_  ( .D(\w_reg/N66 ), .CK(clk), .Q(w_q[63]), .QN() );
  DFF_X2 \w_reg/q_reg_64_  ( .D(\w_reg/N67 ), .CK(clk), .Q(w_q[64]), .QN() );
  DFF_X2 \w_reg/q_reg_65_  ( .D(\w_reg/N68 ), .CK(clk), .Q(w_q[65]), .QN() );
  DFF_X2 \w_reg/q_reg_66_  ( .D(\w_reg/N69 ), .CK(clk), .Q(w_q[66]), .QN() );
  DFF_X2 \w_reg/q_reg_67_  ( .D(\w_reg/N70 ), .CK(clk), .Q(w_q[67]), .QN() );
  DFF_X2 \w_reg/q_reg_68_  ( .D(\w_reg/N71 ), .CK(clk), .Q(w_q[68]), .QN() );
  DFF_X2 \w_reg/q_reg_69_  ( .D(\w_reg/N72 ), .CK(clk), .Q(w_q[69]), .QN() );
  DFF_X2 \w_reg/q_reg_70_  ( .D(\w_reg/N73 ), .CK(clk), .Q(w_q[70]), .QN() );
  DFF_X2 \w_reg/q_reg_71_  ( .D(\w_reg/N74 ), .CK(clk), .Q(w_q[71]), .QN() );
  DFF_X2 \w_reg/q_reg_72_  ( .D(\w_reg/N75 ), .CK(clk), .Q(w_q[72]), .QN() );
  DFF_X2 \w_reg/q_reg_73_  ( .D(\w_reg/N76 ), .CK(clk), .Q(w_q[73]), .QN() );
  DFF_X2 \w_reg/q_reg_74_  ( .D(\w_reg/N77 ), .CK(clk), .Q(w_q[74]), .QN() );
  DFF_X2 \w_reg/q_reg_75_  ( .D(\w_reg/N78 ), .CK(clk), .Q(w_q[75]), .QN() );
  DFF_X2 \w_reg/q_reg_76_  ( .D(\w_reg/N79 ), .CK(clk), .Q(w_q[76]), .QN() );
  DFF_X2 \w_reg/q_reg_77_  ( .D(\w_reg/N80 ), .CK(clk), .Q(w_q[77]), .QN() );
  DFF_X2 \w_reg/q_reg_78_  ( .D(\w_reg/N81 ), .CK(clk), .Q(w_q[78]), .QN() );
  DFF_X2 \w_reg/q_reg_79_  ( .D(\w_reg/N82 ), .CK(clk), .Q(w_q[79]), .QN() );
  DFF_X2 \w_reg/q_reg_80_  ( .D(\w_reg/N83 ), .CK(clk), .Q(w_q[80]), .QN() );
  DFF_X2 \w_reg/q_reg_81_  ( .D(\w_reg/N84 ), .CK(clk), .Q(w_q[81]), .QN() );
  DFF_X2 \w_reg/q_reg_82_  ( .D(\w_reg/N85 ), .CK(clk), .Q(w_q[82]), .QN() );
  DFF_X2 \w_reg/q_reg_83_  ( .D(\w_reg/N86 ), .CK(clk), .Q(w_q[83]), .QN() );
  DFF_X2 \w_reg/q_reg_84_  ( .D(\w_reg/N87 ), .CK(clk), .Q(w_q[84]), .QN() );
  DFF_X2 \w_reg/q_reg_85_  ( .D(\w_reg/N88 ), .CK(clk), .Q(w_q[85]), .QN() );
  DFF_X2 \w_reg/q_reg_86_  ( .D(\w_reg/N89 ), .CK(clk), .Q(w_q[86]), .QN() );
  DFF_X2 \w_reg/q_reg_87_  ( .D(\w_reg/N90 ), .CK(clk), .Q(w_q[87]), .QN() );
  DFF_X2 \w_reg/q_reg_88_  ( .D(\w_reg/N91 ), .CK(clk), .Q(w_q[88]), .QN() );
  DFF_X2 \w_reg/q_reg_89_  ( .D(\w_reg/N92 ), .CK(clk), .Q(w_q[89]), .QN() );
  DFF_X2 \w_reg/q_reg_90_  ( .D(\w_reg/N93 ), .CK(clk), .Q(w_q[90]), .QN() );
  DFF_X2 \w_reg/q_reg_91_  ( .D(\w_reg/N94 ), .CK(clk), .Q(w_q[91]), .QN() );
  DFF_X2 \w_reg/q_reg_92_  ( .D(\w_reg/N95 ), .CK(clk), .Q(w_q[92]), .QN() );
  DFF_X2 \w_reg/q_reg_93_  ( .D(\w_reg/N96 ), .CK(clk), .Q(w_q[93]), .QN() );
  DFF_X2 \w_reg/q_reg_94_  ( .D(\w_reg/N97 ), .CK(clk), .Q(w_q[94]), .QN() );
  DFF_X2 \w_reg/q_reg_95_  ( .D(\w_reg/N98 ), .CK(clk), .Q(w_q[95]), .QN() );
  DFF_X2 \w_reg/q_reg_96_  ( .D(\w_reg/N99 ), .CK(clk), .Q(w_q[96]), .QN() );
  DFF_X2 \w_reg/q_reg_97_  ( .D(\w_reg/N100 ), .CK(clk), .Q(w_q[97]), .QN() );
  DFF_X2 \w_reg/q_reg_98_  ( .D(\w_reg/N101 ), .CK(clk), .Q(w_q[98]), .QN() );
  DFF_X2 \w_reg/q_reg_99_  ( .D(\w_reg/N102 ), .CK(clk), .Q(w_q[99]), .QN() );
  DFF_X2 \w_reg/q_reg_100_  ( .D(\w_reg/N103 ), .CK(clk), .Q(w_q[100]), .QN()
         );
  DFF_X2 \w_reg/q_reg_101_  ( .D(\w_reg/N104 ), .CK(clk), .Q(w_q[101]), .QN()
         );
  DFF_X2 \w_reg/q_reg_102_  ( .D(\w_reg/N105 ), .CK(clk), .Q(w_q[102]), .QN()
         );
  DFF_X2 \w_reg/q_reg_103_  ( .D(\w_reg/N106 ), .CK(clk), .Q(w_q[103]), .QN()
         );
  DFF_X2 \w_reg/q_reg_104_  ( .D(\w_reg/N107 ), .CK(clk), .Q(w_q[104]), .QN()
         );
  DFF_X2 \w_reg/q_reg_105_  ( .D(\w_reg/N108 ), .CK(clk), .Q(w_q[105]), .QN()
         );
  DFF_X2 \w_reg/q_reg_106_  ( .D(\w_reg/N109 ), .CK(clk), .Q(w_q[106]), .QN()
         );
  DFF_X2 \w_reg/q_reg_107_  ( .D(\w_reg/N110 ), .CK(clk), .Q(w_q[107]), .QN()
         );
  DFF_X2 \w_reg/q_reg_108_  ( .D(\w_reg/N111 ), .CK(clk), .Q(w_q[108]), .QN()
         );
  DFF_X2 \w_reg/q_reg_109_  ( .D(\w_reg/N112 ), .CK(clk), .Q(w_q[109]), .QN()
         );
  DFF_X2 \w_reg/q_reg_110_  ( .D(\w_reg/N113 ), .CK(clk), .Q(w_q[110]), .QN()
         );
  DFF_X2 \w_reg/q_reg_111_  ( .D(\w_reg/N114 ), .CK(clk), .Q(w_q[111]), .QN()
         );
  DFF_X2 \w_reg/q_reg_112_  ( .D(\w_reg/N115 ), .CK(clk), .Q(w_q[112]), .QN()
         );
  DFF_X2 \w_reg/q_reg_113_  ( .D(\w_reg/N116 ), .CK(clk), .Q(w_q[113]), .QN()
         );
  DFF_X2 \w_reg/q_reg_114_  ( .D(\w_reg/N117 ), .CK(clk), .Q(w_q[114]), .QN()
         );
  DFF_X2 \w_reg/q_reg_115_  ( .D(\w_reg/N118 ), .CK(clk), .Q(w_q[115]), .QN()
         );
  DFF_X2 \w_reg/q_reg_116_  ( .D(\w_reg/N119 ), .CK(clk), .Q(w_q[116]), .QN()
         );
  DFF_X2 \w_reg/q_reg_117_  ( .D(\w_reg/N120 ), .CK(clk), .Q(w_q[117]), .QN()
         );
  DFF_X2 \w_reg/q_reg_118_  ( .D(\w_reg/N121 ), .CK(clk), .Q(w_q[118]), .QN()
         );
  DFF_X2 \w_reg/q_reg_119_  ( .D(\w_reg/N122 ), .CK(clk), .Q(w_q[119]), .QN()
         );
  DFF_X2 \w_reg/q_reg_120_  ( .D(\w_reg/N123 ), .CK(clk), .Q(w_q[120]), .QN()
         );
  DFF_X2 \w_reg/q_reg_121_  ( .D(\w_reg/N124 ), .CK(clk), .Q(w_q[121]), .QN()
         );
  DFF_X2 \w_reg/q_reg_122_  ( .D(\w_reg/N125 ), .CK(clk), .Q(w_q[122]), .QN()
         );
  DFF_X2 \w_reg/q_reg_123_  ( .D(\w_reg/N126 ), .CK(clk), .Q(w_q[123]), .QN()
         );
  DFF_X2 \w_reg/q_reg_124_  ( .D(\w_reg/N127 ), .CK(clk), .Q(w_q[124]), .QN()
         );
  DFF_X2 \w_reg/q_reg_125_  ( .D(\w_reg/N128 ), .CK(clk), .Q(w_q[125]), .QN()
         );
  DFF_X2 \w_reg/q_reg_126_  ( .D(\w_reg/N129 ), .CK(clk), .Q(w_q[126]), .QN()
         );
  DFF_X2 \w_reg/q_reg_127_  ( .D(\w_reg/N130 ), .CK(clk), .Q(w_q[127]), .QN()
         );
  DFF_X2 \w_reg/q_reg_128_  ( .D(\w_reg/N131 ), .CK(clk), .Q(w_q[128]), .QN()
         );
  DFF_X2 \w_reg/q_reg_129_  ( .D(\w_reg/N132 ), .CK(clk), .Q(w_q[129]), .QN()
         );
  DFF_X2 \w_reg/q_reg_130_  ( .D(\w_reg/N133 ), .CK(clk), .Q(w_q[130]), .QN()
         );
  DFF_X2 \w_reg/q_reg_131_  ( .D(\w_reg/N134 ), .CK(clk), .Q(w_q[131]), .QN()
         );
  DFF_X2 \w_reg/q_reg_132_  ( .D(\w_reg/N135 ), .CK(clk), .Q(w_q[132]), .QN()
         );
  DFF_X2 \w_reg/q_reg_133_  ( .D(\w_reg/N136 ), .CK(clk), .Q(w_q[133]), .QN()
         );
  DFF_X2 \w_reg/q_reg_134_  ( .D(\w_reg/N137 ), .CK(clk), .Q(w_q[134]), .QN()
         );
  DFF_X2 \w_reg/q_reg_135_  ( .D(\w_reg/N138 ), .CK(clk), .Q(w_q[135]), .QN()
         );
  DFF_X2 \w_reg/q_reg_136_  ( .D(\w_reg/N139 ), .CK(clk), .Q(w_q[136]), .QN()
         );
  DFF_X2 \w_reg/q_reg_137_  ( .D(\w_reg/N140 ), .CK(clk), .Q(w_q[137]), .QN()
         );
  DFF_X2 \w_reg/q_reg_138_  ( .D(\w_reg/N141 ), .CK(clk), .Q(w_q[138]), .QN()
         );
  DFF_X2 \w_reg/q_reg_139_  ( .D(\w_reg/N142 ), .CK(clk), .Q(w_q[139]), .QN()
         );
  DFF_X2 \w_reg/q_reg_140_  ( .D(\w_reg/N143 ), .CK(clk), .Q(w_q[140]), .QN()
         );
  DFF_X2 \w_reg/q_reg_141_  ( .D(\w_reg/N144 ), .CK(clk), .Q(w_q[141]), .QN()
         );
  DFF_X2 \w_reg/q_reg_142_  ( .D(\w_reg/N145 ), .CK(clk), .Q(w_q[142]), .QN()
         );
  DFF_X2 \w_reg/q_reg_143_  ( .D(\w_reg/N146 ), .CK(clk), .Q(w_q[143]), .QN()
         );
  DFF_X2 \w_reg/q_reg_144_  ( .D(\w_reg/N147 ), .CK(clk), .Q(w_q[144]), .QN()
         );
  DFF_X2 \w_reg/q_reg_145_  ( .D(\w_reg/N148 ), .CK(clk), .Q(w_q[145]), .QN()
         );
  DFF_X2 \w_reg/q_reg_146_  ( .D(\w_reg/N149 ), .CK(clk), .Q(w_q[146]), .QN()
         );
  DFF_X2 \w_reg/q_reg_147_  ( .D(\w_reg/N150 ), .CK(clk), .Q(w_q[147]), .QN()
         );
  DFF_X2 \w_reg/q_reg_148_  ( .D(\w_reg/N151 ), .CK(clk), .Q(w_q[148]), .QN()
         );
  DFF_X2 \w_reg/q_reg_149_  ( .D(\w_reg/N152 ), .CK(clk), .Q(w_q[149]), .QN()
         );
  DFF_X2 \w_reg/q_reg_150_  ( .D(\w_reg/N153 ), .CK(clk), .Q(w_q[150]), .QN()
         );
  DFF_X2 \w_reg/q_reg_151_  ( .D(\w_reg/N154 ), .CK(clk), .Q(w_q[151]), .QN()
         );
  DFF_X2 \w_reg/q_reg_152_  ( .D(\w_reg/N155 ), .CK(clk), .Q(w_q[152]), .QN()
         );
  DFF_X2 \w_reg/q_reg_153_  ( .D(\w_reg/N156 ), .CK(clk), .Q(w_q[153]), .QN()
         );
  DFF_X2 \w_reg/q_reg_154_  ( .D(\w_reg/N157 ), .CK(clk), .Q(w_q[154]), .QN()
         );
  DFF_X2 \w_reg/q_reg_155_  ( .D(\w_reg/N158 ), .CK(clk), .Q(w_q[155]), .QN()
         );
  DFF_X2 \w_reg/q_reg_156_  ( .D(\w_reg/N159 ), .CK(clk), .Q(w_q[156]), .QN()
         );
  DFF_X2 \w_reg/q_reg_157_  ( .D(\w_reg/N160 ), .CK(clk), .Q(w_q[157]), .QN()
         );
  DFF_X2 \w_reg/q_reg_158_  ( .D(\w_reg/N161 ), .CK(clk), .Q(w_q[158]), .QN()
         );
  DFF_X2 \w_reg/q_reg_159_  ( .D(\w_reg/N162 ), .CK(clk), .Q(w_q[159]), .QN()
         );
  DFF_X2 \w_reg/q_reg_160_  ( .D(\w_reg/N163 ), .CK(clk), .Q(w_q[160]), .QN()
         );
  DFF_X2 \w_reg/q_reg_161_  ( .D(\w_reg/N164 ), .CK(clk), .Q(w_q[161]), .QN()
         );
  DFF_X2 \w_reg/q_reg_162_  ( .D(\w_reg/N165 ), .CK(clk), .Q(w_q[162]), .QN()
         );
  DFF_X2 \w_reg/q_reg_163_  ( .D(\w_reg/N166 ), .CK(clk), .Q(w_q[163]), .QN()
         );
  DFF_X2 \w_reg/q_reg_164_  ( .D(\w_reg/N167 ), .CK(clk), .Q(w_q[164]), .QN()
         );
  DFF_X2 \w_reg/q_reg_165_  ( .D(\w_reg/N168 ), .CK(clk), .Q(w_q[165]), .QN()
         );
  DFF_X2 \w_reg/q_reg_166_  ( .D(\w_reg/N169 ), .CK(clk), .Q(w_q[166]), .QN()
         );
  DFF_X2 \w_reg/q_reg_167_  ( .D(\w_reg/N170 ), .CK(clk), .Q(w_q[167]), .QN()
         );
  DFF_X2 \w_reg/q_reg_168_  ( .D(\w_reg/N171 ), .CK(clk), .Q(w_q[168]), .QN()
         );
  DFF_X2 \w_reg/q_reg_169_  ( .D(\w_reg/N172 ), .CK(clk), .Q(w_q[169]), .QN()
         );
  DFF_X2 \w_reg/q_reg_170_  ( .D(\w_reg/N173 ), .CK(clk), .Q(w_q[170]), .QN()
         );
  DFF_X2 \w_reg/q_reg_171_  ( .D(\w_reg/N174 ), .CK(clk), .Q(w_q[171]), .QN()
         );
  DFF_X2 \w_reg/q_reg_172_  ( .D(\w_reg/N175 ), .CK(clk), .Q(w_q[172]), .QN()
         );
  DFF_X2 \w_reg/q_reg_173_  ( .D(\w_reg/N176 ), .CK(clk), .Q(w_q[173]), .QN()
         );
  DFF_X2 \w_reg/q_reg_174_  ( .D(\w_reg/N177 ), .CK(clk), .Q(w_q[174]), .QN()
         );
  DFF_X2 \w_reg/q_reg_175_  ( .D(\w_reg/N178 ), .CK(clk), .Q(w_q[175]), .QN()
         );
  DFF_X2 \w_reg/q_reg_176_  ( .D(\w_reg/N179 ), .CK(clk), .Q(w_q[176]), .QN()
         );
  DFF_X2 \w_reg/q_reg_177_  ( .D(\w_reg/N180 ), .CK(clk), .Q(w_q[177]), .QN()
         );
  DFF_X2 \w_reg/q_reg_178_  ( .D(\w_reg/N181 ), .CK(clk), .Q(w_q[178]), .QN()
         );
  DFF_X2 \w_reg/q_reg_179_  ( .D(\w_reg/N182 ), .CK(clk), .Q(w_q[179]), .QN()
         );
  DFF_X2 \w_reg/q_reg_180_  ( .D(\w_reg/N183 ), .CK(clk), .Q(w_q[180]), .QN()
         );
  DFF_X2 \w_reg/q_reg_181_  ( .D(\w_reg/N184 ), .CK(clk), .Q(w_q[181]), .QN()
         );
  DFF_X2 \w_reg/q_reg_182_  ( .D(\w_reg/N185 ), .CK(clk), .Q(w_q[182]), .QN()
         );
  DFF_X2 \w_reg/q_reg_183_  ( .D(\w_reg/N186 ), .CK(clk), .Q(w_q[183]), .QN()
         );
  DFF_X2 \w_reg/q_reg_184_  ( .D(\w_reg/N187 ), .CK(clk), .Q(w_q[184]), .QN()
         );
  DFF_X2 \w_reg/q_reg_185_  ( .D(\w_reg/N188 ), .CK(clk), .Q(w_q[185]), .QN()
         );
  DFF_X2 \w_reg/q_reg_186_  ( .D(\w_reg/N189 ), .CK(clk), .Q(w_q[186]), .QN()
         );
  DFF_X2 \w_reg/q_reg_187_  ( .D(\w_reg/N190 ), .CK(clk), .Q(w_q[187]), .QN()
         );
  DFF_X2 \w_reg/q_reg_188_  ( .D(\w_reg/N191 ), .CK(clk), .Q(w_q[188]), .QN()
         );
  DFF_X2 \w_reg/q_reg_189_  ( .D(\w_reg/N192 ), .CK(clk), .Q(w_q[189]), .QN()
         );
  DFF_X2 \w_reg/q_reg_190_  ( .D(\w_reg/N193 ), .CK(clk), .Q(w_q[190]), .QN()
         );
  DFF_X2 \w_reg/q_reg_191_  ( .D(\w_reg/N194 ), .CK(clk), .Q(w_q[191]), .QN()
         );
  DFF_X2 \w_reg/q_reg_192_  ( .D(\w_reg/N195 ), .CK(clk), .Q(w_q[192]), .QN()
         );
  DFF_X2 \w_reg/q_reg_193_  ( .D(\w_reg/N196 ), .CK(clk), .Q(w_q[193]), .QN()
         );
  DFF_X2 \w_reg/q_reg_194_  ( .D(\w_reg/N197 ), .CK(clk), .Q(w_q[194]), .QN()
         );
  DFF_X2 \w_reg/q_reg_195_  ( .D(\w_reg/N198 ), .CK(clk), .Q(w_q[195]), .QN()
         );
  DFF_X2 \w_reg/q_reg_196_  ( .D(\w_reg/N199 ), .CK(clk), .Q(w_q[196]), .QN()
         );
  DFF_X2 \w_reg/q_reg_197_  ( .D(\w_reg/N200 ), .CK(clk), .Q(w_q[197]), .QN()
         );
  DFF_X2 \w_reg/q_reg_198_  ( .D(\w_reg/N201 ), .CK(clk), .Q(w_q[198]), .QN()
         );
  DFF_X2 \w_reg/q_reg_199_  ( .D(\w_reg/N202 ), .CK(clk), .Q(w_q[199]), .QN()
         );
  DFF_X2 \w_reg/q_reg_200_  ( .D(\w_reg/N203 ), .CK(clk), .Q(w_q[200]), .QN()
         );
  DFF_X2 \w_reg/q_reg_201_  ( .D(\w_reg/N204 ), .CK(clk), .Q(w_q[201]), .QN()
         );
  DFF_X2 \w_reg/q_reg_202_  ( .D(\w_reg/N205 ), .CK(clk), .Q(w_q[202]), .QN()
         );
  DFF_X2 \w_reg/q_reg_203_  ( .D(\w_reg/N206 ), .CK(clk), .Q(w_q[203]), .QN()
         );
  DFF_X2 \w_reg/q_reg_204_  ( .D(\w_reg/N207 ), .CK(clk), .Q(w_q[204]), .QN()
         );
  DFF_X2 \w_reg/q_reg_205_  ( .D(\w_reg/N208 ), .CK(clk), .Q(w_q[205]), .QN()
         );
  DFF_X2 \w_reg/q_reg_206_  ( .D(\w_reg/N209 ), .CK(clk), .Q(w_q[206]), .QN()
         );
  DFF_X2 \w_reg/q_reg_207_  ( .D(\w_reg/N210 ), .CK(clk), .Q(w_q[207]), .QN()
         );
  DFF_X2 \w_reg/q_reg_208_  ( .D(\w_reg/N211 ), .CK(clk), .Q(w_q[208]), .QN()
         );
  DFF_X2 \w_reg/q_reg_209_  ( .D(\w_reg/N212 ), .CK(clk), .Q(w_q[209]), .QN()
         );
  DFF_X2 \w_reg/q_reg_210_  ( .D(\w_reg/N213 ), .CK(clk), .Q(w_q[210]), .QN()
         );
  DFF_X2 \w_reg/q_reg_211_  ( .D(\w_reg/N214 ), .CK(clk), .Q(w_q[211]), .QN()
         );
  DFF_X2 \w_reg/q_reg_212_  ( .D(\w_reg/N215 ), .CK(clk), .Q(w_q[212]), .QN()
         );
  DFF_X2 \w_reg/q_reg_213_  ( .D(\w_reg/N216 ), .CK(clk), .Q(w_q[213]), .QN()
         );
  DFF_X2 \w_reg/q_reg_214_  ( .D(\w_reg/N217 ), .CK(clk), .Q(w_q[214]), .QN()
         );
  DFF_X2 \w_reg/q_reg_215_  ( .D(\w_reg/N218 ), .CK(clk), .Q(w_q[215]), .QN()
         );
  DFF_X2 \w_reg/q_reg_216_  ( .D(\w_reg/N219 ), .CK(clk), .Q(w_q[216]), .QN()
         );
  DFF_X2 \w_reg/q_reg_217_  ( .D(\w_reg/N220 ), .CK(clk), .Q(w_q[217]), .QN()
         );
  DFF_X2 \w_reg/q_reg_218_  ( .D(\w_reg/N221 ), .CK(clk), .Q(w_q[218]), .QN()
         );
  DFF_X2 \w_reg/q_reg_219_  ( .D(\w_reg/N222 ), .CK(clk), .Q(w_q[219]), .QN()
         );
  DFF_X2 \w_reg/q_reg_220_  ( .D(\w_reg/N223 ), .CK(clk), .Q(w_q[220]), .QN()
         );
  DFF_X2 \w_reg/q_reg_221_  ( .D(\w_reg/N224 ), .CK(clk), .Q(w_q[221]), .QN()
         );
  DFF_X2 \w_reg/q_reg_222_  ( .D(\w_reg/N225 ), .CK(clk), .Q(w_q[222]), .QN()
         );
  DFF_X2 \w_reg/q_reg_223_  ( .D(\w_reg/N226 ), .CK(clk), .Q(w_q[223]), .QN()
         );
  DFF_X2 \w_reg/q_reg_224_  ( .D(\w_reg/N227 ), .CK(clk), .Q(w_q[224]), .QN()
         );
  DFF_X2 \w_reg/q_reg_225_  ( .D(\w_reg/N228 ), .CK(clk), .Q(w_q[225]), .QN()
         );
  DFF_X2 \w_reg/q_reg_226_  ( .D(\w_reg/N229 ), .CK(clk), .Q(w_q[226]), .QN()
         );
  DFF_X2 \w_reg/q_reg_227_  ( .D(\w_reg/N230 ), .CK(clk), .Q(w_q[227]), .QN()
         );
  DFF_X2 \w_reg/q_reg_228_  ( .D(\w_reg/N231 ), .CK(clk), .Q(w_q[228]), .QN()
         );
  DFF_X2 \w_reg/q_reg_229_  ( .D(\w_reg/N232 ), .CK(clk), .Q(w_q[229]), .QN()
         );
  DFF_X2 \w_reg/q_reg_230_  ( .D(\w_reg/N233 ), .CK(clk), .Q(w_q[230]), .QN()
         );
  DFF_X2 \w_reg/q_reg_231_  ( .D(\w_reg/N234 ), .CK(clk), .Q(w_q[231]), .QN()
         );
  DFF_X2 \w_reg/q_reg_232_  ( .D(\w_reg/N235 ), .CK(clk), .Q(w_q[232]), .QN()
         );
  DFF_X2 \w_reg/q_reg_233_  ( .D(\w_reg/N236 ), .CK(clk), .Q(w_q[233]), .QN()
         );
  DFF_X2 \w_reg/q_reg_234_  ( .D(\w_reg/N237 ), .CK(clk), .Q(w_q[234]), .QN()
         );
  DFF_X2 \w_reg/q_reg_235_  ( .D(\w_reg/N238 ), .CK(clk), .Q(w_q[235]), .QN()
         );
  DFF_X2 \w_reg/q_reg_236_  ( .D(\w_reg/N239 ), .CK(clk), .Q(w_q[236]), .QN()
         );
  DFF_X2 \w_reg/q_reg_237_  ( .D(\w_reg/N240 ), .CK(clk), .Q(w_q[237]), .QN()
         );
  DFF_X2 \w_reg/q_reg_238_  ( .D(\w_reg/N241 ), .CK(clk), .Q(w_q[238]), .QN()
         );
  DFF_X2 \w_reg/q_reg_239_  ( .D(\w_reg/N242 ), .CK(clk), .Q(w_q[239]), .QN()
         );
  DFF_X2 \w_reg/q_reg_240_  ( .D(\w_reg/N243 ), .CK(clk), .Q(w_q[240]), .QN()
         );
  DFF_X2 \w_reg/q_reg_241_  ( .D(\w_reg/N244 ), .CK(clk), .Q(w_q[241]), .QN()
         );
  DFF_X2 \w_reg/q_reg_242_  ( .D(\w_reg/N245 ), .CK(clk), .Q(w_q[242]), .QN()
         );
  DFF_X2 \w_reg/q_reg_243_  ( .D(\w_reg/N246 ), .CK(clk), .Q(w_q[243]), .QN()
         );
  DFF_X2 \w_reg/q_reg_244_  ( .D(\w_reg/N247 ), .CK(clk), .Q(w_q[244]), .QN()
         );
  DFF_X2 \w_reg/q_reg_245_  ( .D(\w_reg/N248 ), .CK(clk), .Q(w_q[245]), .QN()
         );
  DFF_X2 \w_reg/q_reg_246_  ( .D(\w_reg/N249 ), .CK(clk), .Q(w_q[246]), .QN()
         );
  DFF_X2 \w_reg/q_reg_247_  ( .D(\w_reg/N250 ), .CK(clk), .Q(w_q[247]), .QN()
         );
  DFF_X2 \w_reg/q_reg_248_  ( .D(\w_reg/N251 ), .CK(clk), .Q(w_q[248]), .QN()
         );
  DFF_X2 \w_reg/q_reg_249_  ( .D(\w_reg/N252 ), .CK(clk), .Q(w_q[249]), .QN()
         );
  DFF_X2 \w_reg/q_reg_250_  ( .D(\w_reg/N253 ), .CK(clk), .Q(w_q[250]), .QN()
         );
  DFF_X2 \w_reg/q_reg_251_  ( .D(\w_reg/N254 ), .CK(clk), .Q(w_q[251]), .QN()
         );
  DFF_X2 \w_reg/q_reg_252_  ( .D(\w_reg/N255 ), .CK(clk), .Q(w_q[252]), .QN()
         );
  DFF_X2 \w_reg/q_reg_253_  ( .D(\w_reg/N256 ), .CK(clk), .Q(w_q[253]), .QN()
         );
  DFF_X2 \w_reg/q_reg_254_  ( .D(\w_reg/N257 ), .CK(clk), .Q(w_q[254]), .QN()
         );
  DFF_X2 \w_reg/q_reg_255_  ( .D(\w_reg/N258 ), .CK(clk), .Q(w_q[255]), .QN()
         );
  DFF_X2 \w_reg/q_reg_256_  ( .D(\w_reg/N259 ), .CK(clk), .Q(w_q[256]), .QN()
         );
  DFF_X2 \w_reg/q_reg_257_  ( .D(\w_reg/N260 ), .CK(clk), .Q(w_q[257]), .QN()
         );
  DFF_X2 \w_reg/q_reg_258_  ( .D(\w_reg/N261 ), .CK(clk), .Q(w_q[258]), .QN()
         );
  DFF_X2 \w_reg/q_reg_259_  ( .D(\w_reg/N262 ), .CK(clk), .Q(w_q[259]), .QN()
         );
  DFF_X2 \w_reg/q_reg_260_  ( .D(\w_reg/N263 ), .CK(clk), .Q(w_q[260]), .QN()
         );
  DFF_X2 \w_reg/q_reg_261_  ( .D(\w_reg/N264 ), .CK(clk), .Q(w_q[261]), .QN()
         );
  DFF_X2 \w_reg/q_reg_262_  ( .D(\w_reg/N265 ), .CK(clk), .Q(w_q[262]), .QN()
         );
  DFF_X2 \w_reg/q_reg_263_  ( .D(\w_reg/N266 ), .CK(clk), .Q(w_q[263]), .QN()
         );
  DFF_X2 \w_reg/q_reg_264_  ( .D(\w_reg/N267 ), .CK(clk), .Q(w_q[264]), .QN()
         );
  DFF_X2 \w_reg/q_reg_265_  ( .D(\w_reg/N268 ), .CK(clk), .Q(w_q[265]), .QN()
         );
  DFF_X2 \w_reg/q_reg_266_  ( .D(\w_reg/N269 ), .CK(clk), .Q(w_q[266]), .QN()
         );
  DFF_X2 \w_reg/q_reg_267_  ( .D(\w_reg/N270 ), .CK(clk), .Q(w_q[267]), .QN()
         );
  DFF_X2 \w_reg/q_reg_268_  ( .D(\w_reg/N271 ), .CK(clk), .Q(w_q[268]), .QN()
         );
  DFF_X2 \w_reg/q_reg_269_  ( .D(\w_reg/N272 ), .CK(clk), .Q(w_q[269]), .QN()
         );
  DFF_X2 \w_reg/q_reg_270_  ( .D(\w_reg/N273 ), .CK(clk), .Q(w_q[270]), .QN()
         );
  DFF_X2 \w_reg/q_reg_271_  ( .D(\w_reg/N274 ), .CK(clk), .Q(w_q[271]), .QN()
         );
  DFF_X2 \w_reg/q_reg_272_  ( .D(\w_reg/N275 ), .CK(clk), .Q(w_q[272]), .QN()
         );
  DFF_X2 \w_reg/q_reg_273_  ( .D(\w_reg/N276 ), .CK(clk), .Q(w_q[273]), .QN()
         );
  DFF_X2 \w_reg/q_reg_274_  ( .D(\w_reg/N277 ), .CK(clk), .Q(w_q[274]), .QN()
         );
  DFF_X2 \w_reg/q_reg_275_  ( .D(\w_reg/N278 ), .CK(clk), .Q(w_q[275]), .QN()
         );
  DFF_X2 \w_reg/q_reg_276_  ( .D(\w_reg/N279 ), .CK(clk), .Q(w_q[276]), .QN()
         );
  DFF_X2 \w_reg/q_reg_277_  ( .D(\w_reg/N280 ), .CK(clk), .Q(w_q[277]), .QN()
         );
  DFF_X2 \w_reg/q_reg_278_  ( .D(\w_reg/N281 ), .CK(clk), .Q(w_q[278]), .QN()
         );
  DFF_X2 \w_reg/q_reg_279_  ( .D(\w_reg/N282 ), .CK(clk), .Q(w_q[279]), .QN()
         );
  DFF_X2 \w_reg/q_reg_280_  ( .D(\w_reg/N283 ), .CK(clk), .Q(w_q[280]), .QN()
         );
  DFF_X2 \w_reg/q_reg_281_  ( .D(\w_reg/N284 ), .CK(clk), .Q(w_q[281]), .QN()
         );
  DFF_X2 \w_reg/q_reg_282_  ( .D(\w_reg/N285 ), .CK(clk), .Q(w_q[282]), .QN()
         );
  DFF_X2 \w_reg/q_reg_283_  ( .D(\w_reg/N286 ), .CK(clk), .Q(w_q[283]), .QN()
         );
  DFF_X2 \w_reg/q_reg_284_  ( .D(\w_reg/N287 ), .CK(clk), .Q(w_q[284]), .QN()
         );
  DFF_X2 \w_reg/q_reg_285_  ( .D(\w_reg/N288 ), .CK(clk), .Q(w_q[285]), .QN()
         );
  DFF_X2 \w_reg/q_reg_286_  ( .D(\w_reg/N289 ), .CK(clk), .Q(w_q[286]), .QN()
         );
  DFF_X2 \w_reg/q_reg_287_  ( .D(\w_reg/N290 ), .CK(clk), .Q(w_q[287]), .QN()
         );
  DFF_X2 \w_reg/q_reg_288_  ( .D(\w_reg/N291 ), .CK(clk), .Q(w_q[288]), .QN()
         );
  DFF_X2 \w_reg/q_reg_289_  ( .D(\w_reg/N292 ), .CK(clk), .Q(w_q[289]), .QN()
         );
  DFF_X2 \w_reg/q_reg_290_  ( .D(\w_reg/N293 ), .CK(clk), .Q(w_q[290]), .QN()
         );
  DFF_X2 \w_reg/q_reg_291_  ( .D(\w_reg/N294 ), .CK(clk), .Q(w_q[291]), .QN()
         );
  DFF_X2 \w_reg/q_reg_292_  ( .D(\w_reg/N295 ), .CK(clk), .Q(w_q[292]), .QN()
         );
  DFF_X2 \w_reg/q_reg_293_  ( .D(\w_reg/N296 ), .CK(clk), .Q(w_q[293]), .QN()
         );
  DFF_X2 \w_reg/q_reg_294_  ( .D(\w_reg/N297 ), .CK(clk), .Q(w_q[294]), .QN()
         );
  DFF_X2 \w_reg/q_reg_295_  ( .D(\w_reg/N298 ), .CK(clk), .Q(w_q[295]), .QN()
         );
  DFF_X2 \w_reg/q_reg_296_  ( .D(\w_reg/N299 ), .CK(clk), .Q(w_q[296]), .QN()
         );
  DFF_X2 \w_reg/q_reg_297_  ( .D(\w_reg/N300 ), .CK(clk), .Q(w_q[297]), .QN()
         );
  DFF_X2 \w_reg/q_reg_298_  ( .D(\w_reg/N301 ), .CK(clk), .Q(w_q[298]), .QN()
         );
  DFF_X2 \w_reg/q_reg_299_  ( .D(\w_reg/N302 ), .CK(clk), .Q(w_q[299]), .QN()
         );
  DFF_X2 \w_reg/q_reg_300_  ( .D(\w_reg/N303 ), .CK(clk), .Q(w_q[300]), .QN()
         );
  DFF_X2 \w_reg/q_reg_301_  ( .D(\w_reg/N304 ), .CK(clk), .Q(w_q[301]), .QN()
         );
  DFF_X2 \w_reg/q_reg_302_  ( .D(\w_reg/N305 ), .CK(clk), .Q(w_q[302]), .QN()
         );
  DFF_X2 \w_reg/q_reg_303_  ( .D(\w_reg/N306 ), .CK(clk), .Q(w_q[303]), .QN()
         );
  DFF_X2 \w_reg/q_reg_304_  ( .D(\w_reg/N307 ), .CK(clk), .Q(w_q[304]), .QN()
         );
  DFF_X2 \w_reg/q_reg_305_  ( .D(\w_reg/N308 ), .CK(clk), .Q(w_q[305]), .QN()
         );
  DFF_X2 \w_reg/q_reg_306_  ( .D(\w_reg/N309 ), .CK(clk), .Q(w_q[306]), .QN()
         );
  DFF_X2 \w_reg/q_reg_307_  ( .D(\w_reg/N310 ), .CK(clk), .Q(w_q[307]), .QN()
         );
  DFF_X2 \w_reg/q_reg_308_  ( .D(\w_reg/N311 ), .CK(clk), .Q(w_q[308]), .QN()
         );
  DFF_X2 \w_reg/q_reg_309_  ( .D(\w_reg/N312 ), .CK(clk), .Q(w_q[309]), .QN()
         );
  DFF_X2 \w_reg/q_reg_310_  ( .D(\w_reg/N313 ), .CK(clk), .Q(w_q[310]), .QN()
         );
  DFF_X2 \w_reg/q_reg_311_  ( .D(\w_reg/N314 ), .CK(clk), .Q(w_q[311]), .QN()
         );
  DFF_X2 \w_reg/q_reg_312_  ( .D(\w_reg/N315 ), .CK(clk), .Q(w_q[312]), .QN()
         );
  DFF_X2 \w_reg/q_reg_313_  ( .D(\w_reg/N316 ), .CK(clk), .Q(w_q[313]), .QN()
         );
  DFF_X2 \w_reg/q_reg_314_  ( .D(\w_reg/N317 ), .CK(clk), .Q(w_q[314]), .QN()
         );
  DFF_X2 \w_reg/q_reg_315_  ( .D(\w_reg/N318 ), .CK(clk), .Q(w_q[315]), .QN()
         );
  DFF_X2 \w_reg/q_reg_316_  ( .D(\w_reg/N319 ), .CK(clk), .Q(w_q[316]), .QN()
         );
  DFF_X2 \w_reg/q_reg_317_  ( .D(\w_reg/N320 ), .CK(clk), .Q(w_q[317]), .QN()
         );
  DFF_X2 \w_reg/q_reg_318_  ( .D(\w_reg/N321 ), .CK(clk), .Q(w_q[318]), .QN()
         );
  DFF_X2 \w_reg/q_reg_319_  ( .D(\w_reg/N322 ), .CK(clk), .Q(w_q[319]), .QN()
         );
  DFF_X2 \w_reg/q_reg_320_  ( .D(\w_reg/N323 ), .CK(clk), .Q(w_q[320]), .QN()
         );
  DFF_X2 \w_reg/q_reg_321_  ( .D(\w_reg/N324 ), .CK(clk), .Q(w_q[321]), .QN()
         );
  DFF_X2 \w_reg/q_reg_322_  ( .D(\w_reg/N325 ), .CK(clk), .Q(w_q[322]), .QN()
         );
  DFF_X2 \w_reg/q_reg_323_  ( .D(\w_reg/N326 ), .CK(clk), .Q(w_q[323]), .QN()
         );
  DFF_X2 \w_reg/q_reg_324_  ( .D(\w_reg/N327 ), .CK(clk), .Q(w_q[324]), .QN()
         );
  DFF_X2 \w_reg/q_reg_325_  ( .D(\w_reg/N328 ), .CK(clk), .Q(w_q[325]), .QN()
         );
  DFF_X2 \w_reg/q_reg_326_  ( .D(\w_reg/N329 ), .CK(clk), .Q(w_q[326]), .QN()
         );
  DFF_X2 \w_reg/q_reg_327_  ( .D(\w_reg/N330 ), .CK(clk), .Q(w_q[327]), .QN()
         );
  DFF_X2 \w_reg/q_reg_328_  ( .D(\w_reg/N331 ), .CK(clk), .Q(w_q[328]), .QN()
         );
  DFF_X2 \w_reg/q_reg_329_  ( .D(\w_reg/N332 ), .CK(clk), .Q(w_q[329]), .QN()
         );
  DFF_X2 \w_reg/q_reg_330_  ( .D(\w_reg/N333 ), .CK(clk), .Q(w_q[330]), .QN()
         );
  DFF_X2 \w_reg/q_reg_331_  ( .D(\w_reg/N334 ), .CK(clk), .Q(w_q[331]), .QN()
         );
  DFF_X2 \w_reg/q_reg_332_  ( .D(\w_reg/N335 ), .CK(clk), .Q(w_q[332]), .QN()
         );
  DFF_X2 \w_reg/q_reg_333_  ( .D(\w_reg/N336 ), .CK(clk), .Q(w_q[333]), .QN()
         );
  DFF_X2 \w_reg/q_reg_334_  ( .D(\w_reg/N337 ), .CK(clk), .Q(w_q[334]), .QN()
         );
  DFF_X2 \w_reg/q_reg_335_  ( .D(\w_reg/N338 ), .CK(clk), .Q(w_q[335]), .QN()
         );
  DFF_X2 \w_reg/q_reg_336_  ( .D(\w_reg/N339 ), .CK(clk), .Q(w_q[336]), .QN()
         );
  DFF_X2 \w_reg/q_reg_337_  ( .D(\w_reg/N340 ), .CK(clk), .Q(w_q[337]), .QN()
         );
  DFF_X2 \w_reg/q_reg_338_  ( .D(\w_reg/N341 ), .CK(clk), .Q(w_q[338]), .QN()
         );
  DFF_X2 \w_reg/q_reg_339_  ( .D(\w_reg/N342 ), .CK(clk), .Q(w_q[339]), .QN()
         );
  DFF_X2 \w_reg/q_reg_340_  ( .D(\w_reg/N343 ), .CK(clk), .Q(w_q[340]), .QN()
         );
  DFF_X2 \w_reg/q_reg_341_  ( .D(\w_reg/N344 ), .CK(clk), .Q(w_q[341]), .QN()
         );
  DFF_X2 \w_reg/q_reg_342_  ( .D(\w_reg/N345 ), .CK(clk), .Q(w_q[342]), .QN()
         );
  DFF_X2 \w_reg/q_reg_343_  ( .D(\w_reg/N346 ), .CK(clk), .Q(w_q[343]), .QN()
         );
  DFF_X2 \w_reg/q_reg_344_  ( .D(\w_reg/N347 ), .CK(clk), .Q(w_q[344]), .QN()
         );
  DFF_X2 \w_reg/q_reg_345_  ( .D(\w_reg/N348 ), .CK(clk), .Q(w_q[345]), .QN()
         );
  DFF_X2 \w_reg/q_reg_346_  ( .D(\w_reg/N349 ), .CK(clk), .Q(w_q[346]), .QN()
         );
  DFF_X2 \w_reg/q_reg_347_  ( .D(\w_reg/N350 ), .CK(clk), .Q(w_q[347]), .QN()
         );
  DFF_X2 \w_reg/q_reg_348_  ( .D(\w_reg/N351 ), .CK(clk), .Q(w_q[348]), .QN()
         );
  DFF_X2 \w_reg/q_reg_349_  ( .D(\w_reg/N352 ), .CK(clk), .Q(w_q[349]), .QN()
         );
  DFF_X2 \w_reg/q_reg_350_  ( .D(\w_reg/N353 ), .CK(clk), .Q(w_q[350]), .QN()
         );
  DFF_X2 \w_reg/q_reg_351_  ( .D(\w_reg/N354 ), .CK(clk), .Q(w_q[351]), .QN()
         );
  DFF_X2 \w_reg/q_reg_352_  ( .D(\w_reg/N355 ), .CK(clk), .Q(w_q[352]), .QN()
         );
  DFF_X2 \w_reg/q_reg_353_  ( .D(\w_reg/N356 ), .CK(clk), .Q(w_q[353]), .QN()
         );
  DFF_X2 \w_reg/q_reg_354_  ( .D(\w_reg/N357 ), .CK(clk), .Q(w_q[354]), .QN()
         );
  DFF_X2 \w_reg/q_reg_355_  ( .D(\w_reg/N358 ), .CK(clk), .Q(w_q[355]), .QN()
         );
  DFF_X2 \w_reg/q_reg_356_  ( .D(\w_reg/N359 ), .CK(clk), .Q(w_q[356]), .QN()
         );
  DFF_X2 \w_reg/q_reg_357_  ( .D(\w_reg/N360 ), .CK(clk), .Q(w_q[357]), .QN()
         );
  DFF_X2 \w_reg/q_reg_358_  ( .D(\w_reg/N361 ), .CK(clk), .Q(w_q[358]), .QN()
         );
  DFF_X2 \w_reg/q_reg_359_  ( .D(\w_reg/N362 ), .CK(clk), .Q(w_q[359]), .QN()
         );
  DFF_X2 \w_reg/q_reg_360_  ( .D(\w_reg/N363 ), .CK(clk), .Q(w_q[360]), .QN()
         );
  DFF_X2 \w_reg/q_reg_361_  ( .D(\w_reg/N364 ), .CK(clk), .Q(w_q[361]), .QN()
         );
  DFF_X2 \w_reg/q_reg_362_  ( .D(\w_reg/N365 ), .CK(clk), .Q(w_q[362]), .QN()
         );
  DFF_X2 \w_reg/q_reg_363_  ( .D(\w_reg/N366 ), .CK(clk), .Q(w_q[363]), .QN()
         );
  DFF_X2 \w_reg/q_reg_364_  ( .D(\w_reg/N367 ), .CK(clk), .Q(w_q[364]), .QN()
         );
  DFF_X2 \w_reg/q_reg_365_  ( .D(\w_reg/N368 ), .CK(clk), .Q(w_q[365]), .QN()
         );
  DFF_X2 \w_reg/q_reg_366_  ( .D(\w_reg/N369 ), .CK(clk), .Q(w_q[366]), .QN()
         );
  DFF_X2 \w_reg/q_reg_367_  ( .D(\w_reg/N370 ), .CK(clk), .Q(w_q[367]), .QN()
         );
  DFF_X2 \w_reg/q_reg_368_  ( .D(\w_reg/N371 ), .CK(clk), .Q(w_q[368]), .QN()
         );
  DFF_X2 \w_reg/q_reg_369_  ( .D(\w_reg/N372 ), .CK(clk), .Q(w_q[369]), .QN()
         );
  DFF_X2 \w_reg/q_reg_370_  ( .D(\w_reg/N373 ), .CK(clk), .Q(w_q[370]), .QN()
         );
  DFF_X2 \w_reg/q_reg_371_  ( .D(\w_reg/N374 ), .CK(clk), .Q(w_q[371]), .QN()
         );
  DFF_X2 \w_reg/q_reg_372_  ( .D(\w_reg/N375 ), .CK(clk), .Q(w_q[372]), .QN()
         );
  DFF_X2 \w_reg/q_reg_373_  ( .D(\w_reg/N376 ), .CK(clk), .Q(w_q[373]), .QN()
         );
  DFF_X2 \w_reg/q_reg_374_  ( .D(\w_reg/N377 ), .CK(clk), .Q(w_q[374]), .QN()
         );
  DFF_X2 \w_reg/q_reg_375_  ( .D(\w_reg/N378 ), .CK(clk), .Q(w_q[375]), .QN()
         );
  DFF_X2 \w_reg/q_reg_376_  ( .D(\w_reg/N379 ), .CK(clk), .Q(w_q[376]), .QN()
         );
  DFF_X2 \w_reg/q_reg_377_  ( .D(\w_reg/N380 ), .CK(clk), .Q(w_q[377]), .QN()
         );
  DFF_X2 \w_reg/q_reg_378_  ( .D(\w_reg/N381 ), .CK(clk), .Q(w_q[378]), .QN()
         );
  DFF_X2 \w_reg/q_reg_379_  ( .D(\w_reg/N382 ), .CK(clk), .Q(w_q[379]), .QN()
         );
  DFF_X2 \w_reg/q_reg_380_  ( .D(\w_reg/N383 ), .CK(clk), .Q(w_q[380]), .QN()
         );
  DFF_X2 \w_reg/q_reg_381_  ( .D(\w_reg/N384 ), .CK(clk), .Q(w_q[381]), .QN()
         );
  DFF_X2 \w_reg/q_reg_382_  ( .D(\w_reg/N385 ), .CK(clk), .Q(w_q[382]), .QN()
         );
  DFF_X2 \w_reg/q_reg_383_  ( .D(\w_reg/N386 ), .CK(clk), .Q(w_q[383]), .QN()
         );
  DFF_X2 \w_reg/q_reg_384_  ( .D(\w_reg/N387 ), .CK(clk), .Q(w_q[384]), .QN()
         );
  DFF_X2 \w_reg/q_reg_385_  ( .D(\w_reg/N388 ), .CK(clk), .Q(w_q[385]), .QN()
         );
  DFF_X2 \w_reg/q_reg_386_  ( .D(\w_reg/N389 ), .CK(clk), .Q(w_q[386]), .QN()
         );
  DFF_X2 \w_reg/q_reg_387_  ( .D(\w_reg/N390 ), .CK(clk), .Q(w_q[387]), .QN()
         );
  DFF_X2 \w_reg/q_reg_388_  ( .D(\w_reg/N391 ), .CK(clk), .Q(w_q[388]), .QN()
         );
  DFF_X2 \w_reg/q_reg_389_  ( .D(\w_reg/N392 ), .CK(clk), .Q(w_q[389]), .QN()
         );
  DFF_X2 \w_reg/q_reg_390_  ( .D(\w_reg/N393 ), .CK(clk), .Q(w_q[390]), .QN()
         );
  DFF_X2 \w_reg/q_reg_391_  ( .D(\w_reg/N394 ), .CK(clk), .Q(w_q[391]), .QN()
         );
  DFF_X2 \w_reg/q_reg_392_  ( .D(\w_reg/N395 ), .CK(clk), .Q(w_q[392]), .QN()
         );
  DFF_X2 \w_reg/q_reg_393_  ( .D(\w_reg/N396 ), .CK(clk), .Q(w_q[393]), .QN()
         );
  DFF_X2 \w_reg/q_reg_394_  ( .D(\w_reg/N397 ), .CK(clk), .Q(w_q[394]), .QN()
         );
  DFF_X2 \w_reg/q_reg_395_  ( .D(\w_reg/N398 ), .CK(clk), .Q(w_q[395]), .QN()
         );
  DFF_X2 \w_reg/q_reg_396_  ( .D(\w_reg/N399 ), .CK(clk), .Q(w_q[396]), .QN()
         );
  DFF_X2 \w_reg/q_reg_397_  ( .D(\w_reg/N400 ), .CK(clk), .Q(w_q[397]), .QN()
         );
  DFF_X2 \w_reg/q_reg_398_  ( .D(\w_reg/N401 ), .CK(clk), .Q(w_q[398]), .QN()
         );
  DFF_X2 \w_reg/q_reg_399_  ( .D(\w_reg/N402 ), .CK(clk), .Q(w_q[399]), .QN()
         );
  DFF_X2 \w_reg/q_reg_400_  ( .D(\w_reg/N403 ), .CK(clk), .Q(w_q[400]), .QN()
         );
  DFF_X2 \w_reg/q_reg_401_  ( .D(\w_reg/N404 ), .CK(clk), .Q(w_q[401]), .QN()
         );
  DFF_X2 \w_reg/q_reg_402_  ( .D(\w_reg/N405 ), .CK(clk), .Q(w_q[402]), .QN()
         );
  DFF_X2 \w_reg/q_reg_403_  ( .D(\w_reg/N406 ), .CK(clk), .Q(w_q[403]), .QN()
         );
  DFF_X2 \w_reg/q_reg_404_  ( .D(\w_reg/N407 ), .CK(clk), .Q(w_q[404]), .QN()
         );
  DFF_X2 \w_reg/q_reg_405_  ( .D(\w_reg/N408 ), .CK(clk), .Q(w_q[405]), .QN()
         );
  DFF_X2 \w_reg/q_reg_406_  ( .D(\w_reg/N409 ), .CK(clk), .Q(w_q[406]), .QN()
         );
  DFF_X2 \w_reg/q_reg_407_  ( .D(\w_reg/N410 ), .CK(clk), .Q(w_q[407]), .QN()
         );
  DFF_X2 \w_reg/q_reg_408_  ( .D(\w_reg/N411 ), .CK(clk), .Q(w_q[408]), .QN()
         );
  DFF_X2 \w_reg/q_reg_409_  ( .D(\w_reg/N412 ), .CK(clk), .Q(w_q[409]), .QN()
         );
  DFF_X2 \w_reg/q_reg_410_  ( .D(\w_reg/N413 ), .CK(clk), .Q(w_q[410]), .QN()
         );
  DFF_X2 \w_reg/q_reg_411_  ( .D(\w_reg/N414 ), .CK(clk), .Q(w_q[411]), .QN()
         );
  DFF_X2 \w_reg/q_reg_412_  ( .D(\w_reg/N415 ), .CK(clk), .Q(w_q[412]), .QN()
         );
  DFF_X2 \w_reg/q_reg_413_  ( .D(\w_reg/N416 ), .CK(clk), .Q(w_q[413]), .QN()
         );
  DFF_X2 \w_reg/q_reg_414_  ( .D(\w_reg/N417 ), .CK(clk), .Q(w_q[414]), .QN()
         );
  DFF_X2 \w_reg/q_reg_415_  ( .D(\w_reg/N418 ), .CK(clk), .Q(w_q[415]), .QN()
         );
  DFF_X2 \w_reg/q_reg_416_  ( .D(\w_reg/N419 ), .CK(clk), .Q(w_q[416]), .QN()
         );
  DFF_X2 \w_reg/q_reg_417_  ( .D(\w_reg/N420 ), .CK(clk), .Q(w_q[417]), .QN()
         );
  DFF_X2 \w_reg/q_reg_418_  ( .D(\w_reg/N421 ), .CK(clk), .Q(w_q[418]), .QN()
         );
  DFF_X2 \w_reg/q_reg_419_  ( .D(\w_reg/N422 ), .CK(clk), .Q(w_q[419]), .QN()
         );
  DFF_X2 \w_reg/q_reg_420_  ( .D(\w_reg/N423 ), .CK(clk), .Q(w_q[420]), .QN()
         );
  DFF_X2 \w_reg/q_reg_421_  ( .D(\w_reg/N424 ), .CK(clk), .Q(w_q[421]), .QN()
         );
  DFF_X2 \w_reg/q_reg_422_  ( .D(\w_reg/N425 ), .CK(clk), .Q(w_q[422]), .QN()
         );
  DFF_X2 \w_reg/q_reg_423_  ( .D(\w_reg/N426 ), .CK(clk), .Q(w_q[423]), .QN()
         );
  DFF_X2 \w_reg/q_reg_424_  ( .D(\w_reg/N427 ), .CK(clk), .Q(w_q[424]), .QN()
         );
  DFF_X2 \w_reg/q_reg_425_  ( .D(\w_reg/N428 ), .CK(clk), .Q(w_q[425]), .QN()
         );
  DFF_X2 \w_reg/q_reg_426_  ( .D(\w_reg/N429 ), .CK(clk), .Q(w_q[426]), .QN()
         );
  DFF_X2 \w_reg/q_reg_427_  ( .D(\w_reg/N430 ), .CK(clk), .Q(w_q[427]), .QN()
         );
  DFF_X2 \w_reg/q_reg_428_  ( .D(\w_reg/N431 ), .CK(clk), .Q(w_q[428]), .QN()
         );
  DFF_X2 \w_reg/q_reg_429_  ( .D(\w_reg/N432 ), .CK(clk), .Q(w_q[429]), .QN()
         );
  DFF_X2 \w_reg/q_reg_430_  ( .D(\w_reg/N433 ), .CK(clk), .Q(w_q[430]), .QN()
         );
  DFF_X2 \w_reg/q_reg_431_  ( .D(\w_reg/N434 ), .CK(clk), .Q(w_q[431]), .QN()
         );
  DFF_X2 \w_reg/q_reg_432_  ( .D(\w_reg/N435 ), .CK(clk), .Q(w_q[432]), .QN()
         );
  DFF_X2 \w_reg/q_reg_433_  ( .D(\w_reg/N436 ), .CK(clk), .Q(w_q[433]), .QN()
         );
  DFF_X2 \w_reg/q_reg_434_  ( .D(\w_reg/N437 ), .CK(clk), .Q(w_q[434]), .QN()
         );
  DFF_X2 \w_reg/q_reg_435_  ( .D(\w_reg/N438 ), .CK(clk), .Q(w_q[435]), .QN()
         );
  DFF_X2 \w_reg/q_reg_436_  ( .D(\w_reg/N439 ), .CK(clk), .Q(w_q[436]), .QN()
         );
  DFF_X2 \w_reg/q_reg_437_  ( .D(\w_reg/N440 ), .CK(clk), .Q(w_q[437]), .QN()
         );
  DFF_X2 \w_reg/q_reg_438_  ( .D(\w_reg/N441 ), .CK(clk), .Q(w_q[438]), .QN()
         );
  DFF_X2 \w_reg/q_reg_439_  ( .D(\w_reg/N442 ), .CK(clk), .Q(w_q[439]), .QN()
         );
  DFF_X2 \w_reg/q_reg_440_  ( .D(\w_reg/N443 ), .CK(clk), .Q(w_q[440]), .QN()
         );
  DFF_X2 \w_reg/q_reg_441_  ( .D(\w_reg/N444 ), .CK(clk), .Q(w_q[441]), .QN()
         );
  DFF_X2 \w_reg/q_reg_442_  ( .D(\w_reg/N445 ), .CK(clk), .Q(w_q[442]), .QN()
         );
  DFF_X2 \w_reg/q_reg_443_  ( .D(\w_reg/N446 ), .CK(clk), .Q(w_q[443]), .QN()
         );
  DFF_X2 \w_reg/q_reg_444_  ( .D(\w_reg/N447 ), .CK(clk), .Q(w_q[444]), .QN()
         );
  DFF_X2 \w_reg/q_reg_445_  ( .D(\w_reg/N448 ), .CK(clk), .Q(w_q[445]), .QN()
         );
  DFF_X2 \w_reg/q_reg_446_  ( .D(\w_reg/N449 ), .CK(clk), .Q(w_q[446]), .QN()
         );
  DFF_X2 \w_reg/q_reg_447_  ( .D(\w_reg/N450 ), .CK(clk), .Q(w_q[447]), .QN()
         );
  DFF_X2 \w_reg/q_reg_448_  ( .D(\w_reg/N451 ), .CK(clk), .Q(w_q[448]), .QN()
         );
  DFF_X2 \w_reg/q_reg_449_  ( .D(\w_reg/N452 ), .CK(clk), .Q(w_q[449]), .QN()
         );
  DFF_X2 \w_reg/q_reg_450_  ( .D(\w_reg/N453 ), .CK(clk), .Q(w_q[450]), .QN()
         );
  DFF_X2 \w_reg/q_reg_451_  ( .D(\w_reg/N454 ), .CK(clk), .Q(w_q[451]), .QN()
         );
  DFF_X2 \w_reg/q_reg_452_  ( .D(\w_reg/N455 ), .CK(clk), .Q(w_q[452]), .QN()
         );
  DFF_X2 \w_reg/q_reg_453_  ( .D(\w_reg/N456 ), .CK(clk), .Q(w_q[453]), .QN()
         );
  DFF_X2 \w_reg/q_reg_454_  ( .D(\w_reg/N457 ), .CK(clk), .Q(w_q[454]), .QN()
         );
  DFF_X2 \w_reg/q_reg_455_  ( .D(\w_reg/N458 ), .CK(clk), .Q(w_q[455]), .QN()
         );
  DFF_X2 \w_reg/q_reg_456_  ( .D(\w_reg/N459 ), .CK(clk), .Q(w_q[456]), .QN()
         );
  DFF_X2 \w_reg/q_reg_457_  ( .D(\w_reg/N460 ), .CK(clk), .Q(w_q[457]), .QN()
         );
  DFF_X2 \w_reg/q_reg_458_  ( .D(\w_reg/N461 ), .CK(clk), .Q(w_q[458]), .QN()
         );
  DFF_X2 \w_reg/q_reg_459_  ( .D(\w_reg/N462 ), .CK(clk), .Q(w_q[459]), .QN()
         );
  DFF_X2 \w_reg/q_reg_460_  ( .D(\w_reg/N463 ), .CK(clk), .Q(w_q[460]), .QN()
         );
  DFF_X2 \w_reg/q_reg_461_  ( .D(\w_reg/N464 ), .CK(clk), .Q(w_q[461]), .QN()
         );
  DFF_X2 \w_reg/q_reg_462_  ( .D(\w_reg/N465 ), .CK(clk), .Q(w_q[462]), .QN()
         );
  DFF_X2 \w_reg/q_reg_463_  ( .D(\w_reg/N466 ), .CK(clk), .Q(w_q[463]), .QN()
         );
  DFF_X2 \w_reg/q_reg_464_  ( .D(\w_reg/N467 ), .CK(clk), .Q(w_q[464]), .QN()
         );
  DFF_X2 \w_reg/q_reg_465_  ( .D(\w_reg/N468 ), .CK(clk), .Q(w_q[465]), .QN()
         );
  DFF_X2 \w_reg/q_reg_466_  ( .D(\w_reg/N469 ), .CK(clk), .Q(w_q[466]), .QN()
         );
  DFF_X2 \w_reg/q_reg_467_  ( .D(\w_reg/N470 ), .CK(clk), .Q(w_q[467]), .QN()
         );
  DFF_X2 \w_reg/q_reg_468_  ( .D(\w_reg/N471 ), .CK(clk), .Q(w_q[468]), .QN()
         );
  DFF_X2 \w_reg/q_reg_469_  ( .D(\w_reg/N472 ), .CK(clk), .Q(w_q[469]), .QN()
         );
  DFF_X2 \w_reg/q_reg_470_  ( .D(\w_reg/N473 ), .CK(clk), .Q(w_q[470]), .QN()
         );
  DFF_X2 \w_reg/q_reg_471_  ( .D(\w_reg/N474 ), .CK(clk), .Q(w_q[471]), .QN()
         );
  DFF_X2 \w_reg/q_reg_472_  ( .D(\w_reg/N475 ), .CK(clk), .Q(w_q[472]), .QN()
         );
  DFF_X2 \w_reg/q_reg_473_  ( .D(\w_reg/N476 ), .CK(clk), .Q(w_q[473]), .QN()
         );
  DFF_X2 \w_reg/q_reg_474_  ( .D(\w_reg/N477 ), .CK(clk), .Q(w_q[474]), .QN()
         );
  DFF_X2 \w_reg/q_reg_475_  ( .D(\w_reg/N478 ), .CK(clk), .Q(w_q[475]), .QN()
         );
  DFF_X2 \w_reg/q_reg_476_  ( .D(\w_reg/N479 ), .CK(clk), .Q(w_q[476]), .QN()
         );
  DFF_X2 \w_reg/q_reg_477_  ( .D(\w_reg/N480 ), .CK(clk), .Q(w_q[477]), .QN()
         );
  DFF_X2 \w_reg/q_reg_478_  ( .D(\w_reg/N481 ), .CK(clk), .Q(w_q[478]), .QN()
         );
  DFF_X2 \w_reg/q_reg_479_  ( .D(\w_reg/N482 ), .CK(clk), .Q(w_q[479]), .QN()
         );
  DFF_X2 \w_reg/q_reg_480_  ( .D(\w_reg/N483 ), .CK(clk), .Q(w[0]), .QN() );
  DFF_X2 \w_reg/q_reg_481_  ( .D(\w_reg/N484 ), .CK(clk), .Q(w[1]), .QN() );
  DFF_X2 \w_reg/q_reg_482_  ( .D(\w_reg/N485 ), .CK(clk), .Q(w[2]), .QN() );
  DFF_X2 \w_reg/q_reg_483_  ( .D(\w_reg/N486 ), .CK(clk), .Q(w[3]), .QN() );
  DFF_X2 \w_reg/q_reg_484_  ( .D(\w_reg/N487 ), .CK(clk), .Q(w[4]), .QN() );
  DFF_X2 \w_reg/q_reg_485_  ( .D(\w_reg/N488 ), .CK(clk), .Q(w[5]), .QN() );
  DFF_X2 \w_reg/q_reg_486_  ( .D(\w_reg/N489 ), .CK(clk), .Q(w[6]), .QN() );
  DFF_X2 \w_reg/q_reg_487_  ( .D(\w_reg/N490 ), .CK(clk), .Q(w[7]), .QN() );
  DFF_X2 \w_reg/q_reg_488_  ( .D(\w_reg/N491 ), .CK(clk), .Q(w[8]), .QN() );
  DFF_X2 \w_reg/q_reg_489_  ( .D(\w_reg/N492 ), .CK(clk), .Q(w[9]), .QN() );
  DFF_X2 \w_reg/q_reg_490_  ( .D(\w_reg/N493 ), .CK(clk), .Q(w[10]), .QN() );
  DFF_X2 \w_reg/q_reg_491_  ( .D(\w_reg/N494 ), .CK(clk), .Q(w[11]), .QN() );
  DFF_X2 \w_reg/q_reg_492_  ( .D(\w_reg/N495 ), .CK(clk), .Q(w[12]), .QN() );
  DFF_X2 \w_reg/q_reg_493_  ( .D(\w_reg/N496 ), .CK(clk), .Q(w[13]), .QN() );
  DFF_X2 \w_reg/q_reg_494_  ( .D(\w_reg/N497 ), .CK(clk), .Q(w[14]), .QN() );
  DFF_X2 \w_reg/q_reg_495_  ( .D(\w_reg/N498 ), .CK(clk), .Q(w[15]), .QN() );
  DFF_X2 \w_reg/q_reg_496_  ( .D(\w_reg/N499 ), .CK(clk), .Q(w[16]), .QN() );
  DFF_X2 \w_reg/q_reg_497_  ( .D(\w_reg/N500 ), .CK(clk), .Q(w[17]), .QN() );
  DFF_X2 \w_reg/q_reg_498_  ( .D(\w_reg/N501 ), .CK(clk), .Q(w[18]), .QN() );
  DFF_X2 \w_reg/q_reg_499_  ( .D(\w_reg/N502 ), .CK(clk), .Q(w[19]), .QN() );
  DFF_X2 \w_reg/q_reg_500_  ( .D(\w_reg/N503 ), .CK(clk), .Q(w[20]), .QN() );
  DFF_X2 \w_reg/q_reg_501_  ( .D(\w_reg/N504 ), .CK(clk), .Q(w[21]), .QN() );
  DFF_X2 \w_reg/q_reg_502_  ( .D(\w_reg/N505 ), .CK(clk), .Q(w[22]), .QN() );
  DFF_X2 \w_reg/q_reg_503_  ( .D(\w_reg/N506 ), .CK(clk), .Q(w[23]), .QN() );
  DFF_X2 \w_reg/q_reg_504_  ( .D(\w_reg/N507 ), .CK(clk), .Q(w[24]), .QN() );
  DFF_X2 \w_reg/q_reg_505_  ( .D(\w_reg/N508 ), .CK(clk), .Q(w[25]), .QN() );
  DFF_X2 \w_reg/q_reg_506_  ( .D(\w_reg/N509 ), .CK(clk), .Q(w[26]), .QN() );
  DFF_X2 \w_reg/q_reg_507_  ( .D(\w_reg/N510 ), .CK(clk), .Q(w[27]), .QN() );
  DFF_X2 \w_reg/q_reg_508_  ( .D(\w_reg/N511 ), .CK(clk), .Q(w[28]), .QN() );
  DFF_X2 \w_reg/q_reg_509_  ( .D(\w_reg/N512 ), .CK(clk), .Q(w[29]), .QN() );
  DFF_X2 \w_reg/q_reg_510_  ( .D(\w_reg/N513 ), .CK(clk), .Q(w[30]), .QN() );
  DFF_X2 \w_reg/q_reg_511_  ( .D(\w_reg/N514 ), .CK(clk), .Q(w[31]), .QN() );
  AND2_X2 \cv_reg/U179  ( .A1(cv_d[137]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N140 ) );
  AND2_X2 \cv_reg/U178  ( .A1(cv_d[136]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N139 ) );
  AND2_X2 \cv_reg/U177  ( .A1(cv_d[135]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N138 ) );
  AND2_X2 \cv_reg/U176  ( .A1(cv_d[134]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N137 ) );
  AND2_X2 \cv_reg/U175  ( .A1(cv_d[133]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N136 ) );
  AND2_X2 \cv_reg/U174  ( .A1(cv_d[132]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N135 ) );
  AND2_X2 \cv_reg/U173  ( .A1(cv_d[131]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N134 ) );
  AND2_X2 \cv_reg/U172  ( .A1(cv_d[130]), .A2(\cv_reg/n230 ), .ZN(
        \cv_reg/N133 ) );
  AND2_X2 \cv_reg/U171  ( .A1(cv_d[129]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N132 ) );
  AND2_X2 \cv_reg/U170  ( .A1(cv_d[128]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N131 ) );
  AND2_X2 \cv_reg/U169  ( .A1(cv_d[111]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N114 ) );
  AND2_X2 \cv_reg/U168  ( .A1(cv_d[110]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N113 ) );
  AND2_X2 \cv_reg/U167  ( .A1(cv_d[109]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N112 ) );
  AND2_X2 \cv_reg/U166  ( .A1(cv_d[108]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N111 ) );
  AND2_X2 \cv_reg/U165  ( .A1(cv_d[107]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N110 ) );
  AND2_X2 \cv_reg/U164  ( .A1(cv_d[106]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N109 ) );
  AND2_X2 \cv_reg/U163  ( .A1(cv_d[105]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N108 ) );
  AND2_X2 \cv_reg/U162  ( .A1(cv_d[104]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N107 ) );
  AND2_X2 \cv_reg/U161  ( .A1(cv_d[103]), .A2(\cv_reg/n220 ), .ZN(
        \cv_reg/N106 ) );
  AND2_X2 \cv_reg/U160  ( .A1(cv_d[102]), .A2(\cv_reg/n210 ), .ZN(
        \cv_reg/N105 ) );
  AND2_X2 \cv_reg/U159  ( .A1(cv_d[101]), .A2(\cv_reg/n210 ), .ZN(
        \cv_reg/N104 ) );
  AND2_X2 \cv_reg/U158  ( .A1(cv_d[100]), .A2(\cv_reg/n210 ), .ZN(
        \cv_reg/N103 ) );
  AND2_X2 \cv_reg/U157  ( .A1(cv_d[99]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N102 ) );
  AND2_X2 \cv_reg/U156  ( .A1(cv_d[98]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N101 ) );
  AND2_X2 \cv_reg/U155  ( .A1(cv_d[97]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N100 ) );
  AND2_X2 \cv_reg/U154  ( .A1(cv_d[96]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N99 )
         );
  AND2_X2 \cv_reg/U153  ( .A1(cv_d[79]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N82 )
         );
  AND2_X2 \cv_reg/U152  ( .A1(cv_d[78]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N81 )
         );
  AND2_X2 \cv_reg/U151  ( .A1(cv_d[77]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N80 )
         );
  AND2_X2 \cv_reg/U150  ( .A1(cv_d[76]), .A2(\cv_reg/n210 ), .ZN(\cv_reg/N79 )
         );
  AND2_X2 \cv_reg/U149  ( .A1(cv_d[75]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N78 )
         );
  AND2_X2 \cv_reg/U148  ( .A1(cv_d[74]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N77 )
         );
  AND2_X2 \cv_reg/U147  ( .A1(cv_d[73]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N76 )
         );
  AND2_X2 \cv_reg/U146  ( .A1(cv_d[72]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N75 )
         );
  AND2_X2 \cv_reg/U140  ( .A1(cv_d[71]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N74 )
         );
  AND2_X2 \cv_reg/U129  ( .A1(cv_d[70]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N73 )
         );
  AND2_X2 \cv_reg/U127  ( .A1(cv_d[69]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N72 )
         );
  AND2_X2 \cv_reg/U126  ( .A1(cv_d[68]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N71 )
         );
  AND2_X2 \cv_reg/U125  ( .A1(cv_d[67]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N70 )
         );
  AND2_X2 \cv_reg/U124  ( .A1(cv_d[66]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N69 )
         );
  AND2_X2 \cv_reg/U123  ( .A1(cv_d[65]), .A2(\cv_reg/n200 ), .ZN(\cv_reg/N68 )
         );
  AND2_X2 \cv_reg/U122  ( .A1(cv_d[64]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N67 )
         );
  AND2_X2 \cv_reg/U121  ( .A1(cv_d[47]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N50 )
         );
  AND2_X2 \cv_reg/U120  ( .A1(cv_d[46]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N49 )
         );
  AND2_X2 \cv_reg/U119  ( .A1(cv_d[45]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N48 )
         );
  AND2_X2 \cv_reg/U118  ( .A1(cv_d[44]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N47 )
         );
  AND2_X2 \cv_reg/U117  ( .A1(cv_d[43]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N46 )
         );
  AND2_X2 \cv_reg/U116  ( .A1(cv_d[42]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N45 )
         );
  AND2_X2 \cv_reg/U115  ( .A1(cv_d[41]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N44 )
         );
  AND2_X2 \cv_reg/U114  ( .A1(cv_d[40]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N43 )
         );
  AND2_X2 \cv_reg/U113  ( .A1(cv_d[39]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N42 )
         );
  AND2_X2 \cv_reg/U112  ( .A1(cv_d[38]), .A2(\cv_reg/n190 ), .ZN(\cv_reg/N41 )
         );
  AND2_X2 \cv_reg/U111  ( .A1(cv_d[37]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N40 )
         );
  AND2_X2 \cv_reg/U110  ( .A1(cv_d[36]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N39 )
         );
  AND2_X2 \cv_reg/U109  ( .A1(cv_d[35]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N38 )
         );
  AND2_X2 \cv_reg/U108  ( .A1(cv_d[34]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N37 )
         );
  AND2_X2 \cv_reg/U107  ( .A1(cv_d[33]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N36 )
         );
  AND2_X2 \cv_reg/U106  ( .A1(cv_d[32]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N35 )
         );
  AND2_X2 \cv_reg/U105  ( .A1(cv_d[15]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N18 )
         );
  AND2_X2 \cv_reg/U102  ( .A1(cv_d[14]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N17 )
         );
  AND2_X2 \cv_reg/U101  ( .A1(cv_d[13]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N16 )
         );
  AND2_X2 \cv_reg/U97  ( .A1(cv_d[12]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N15 )
         );
  AND2_X2 \cv_reg/U96  ( .A1(cv_d[11]), .A2(\cv_reg/n180 ), .ZN(\cv_reg/N14 )
         );
  AND2_X2 \cv_reg/U95  ( .A1(cv_d[10]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N13 )
         );
  AND2_X2 \cv_reg/U92  ( .A1(cv_d[9]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N12 )
         );
  AND2_X2 \cv_reg/U91  ( .A1(cv_d[8]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N11 )
         );
  AND2_X2 \cv_reg/U79  ( .A1(cv_d[7]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N10 )
         );
  AND2_X2 \cv_reg/U73  ( .A1(cv_d[6]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N9 ) );
  AND2_X2 \cv_reg/U72  ( .A1(cv_d[5]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N8 ) );
  AND2_X2 \cv_reg/U71  ( .A1(cv_d[4]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N7 ) );
  AND2_X2 \cv_reg/U70  ( .A1(cv_d[3]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N6 ) );
  AND2_X2 \cv_reg/U69  ( .A1(cv_d[2]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N5 ) );
  AND2_X2 \cv_reg/U68  ( .A1(cv_d[1]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N4 ) );
  AND2_X2 \cv_reg/U67  ( .A1(cv_d[0]), .A2(\cv_reg/n170 ), .ZN(\cv_reg/N3 ) );
  INV_X4 \cv_reg/U66  ( .A(n7117), .ZN(\cv_reg/n330 ) );
  INV_X4 \cv_reg/U65  ( .A(\cv_reg/n330 ), .ZN(\cv_reg/n320 ) );
  INV_X4 \cv_reg/U64  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n310 ) );
  INV_X4 \cv_reg/U63  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n220 ) );
  INV_X4 \cv_reg/U62  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n210 ) );
  INV_X4 \cv_reg/U61  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n200 ) );
  INV_X4 \cv_reg/U60  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n190 ) );
  INV_X4 \cv_reg/U59  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n180 ) );
  INV_X4 \cv_reg/U58  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n170 ) );
  INV_X4 \cv_reg/U57  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n280 ) );
  INV_X4 \cv_reg/U56  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n290 ) );
  INV_X4 \cv_reg/U46  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n300 ) );
  INV_X4 \cv_reg/U38  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n240 ) );
  INV_X4 \cv_reg/U37  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n230 ) );
  INV_X4 \cv_reg/U36  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n250 ) );
  INV_X4 \cv_reg/U35  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n260 ) );
  INV_X4 \cv_reg/U34  ( .A(\cv_reg/n320 ), .ZN(\cv_reg/n270 ) );
  AND2_X1 \cv_reg/U33  ( .A1(cv_d[157]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N160 ) );
  AND2_X1 \cv_reg/U32  ( .A1(cv_d[156]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N159 ) );
  AND2_X1 \cv_reg/U31  ( .A1(cv_d[152]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N155 ) );
  AND2_X1 \cv_reg/U30  ( .A1(cv_d[151]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N154 ) );
  AND2_X1 \cv_reg/U29  ( .A1(cv_d[148]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N151 ) );
  AND2_X1 \cv_reg/U28  ( .A1(cv_d[147]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N150 ) );
  AND2_X1 \cv_reg/U27  ( .A1(cv_d[146]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N149 ) );
  AND2_X1 \cv_reg/U26  ( .A1(cv_d[145]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N148 ) );
  AND2_X1 \cv_reg/U25  ( .A1(cv_d[144]), .A2(\cv_reg/n300 ), .ZN(\cv_reg/N147 ) );
  AND2_X1 \cv_reg/U24  ( .A1(cv_d[143]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N146 ) );
  AND2_X1 \cv_reg/U23  ( .A1(cv_d[142]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N145 ) );
  AND2_X1 \cv_reg/U22  ( .A1(cv_d[141]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N144 ) );
  AND2_X1 \cv_reg/U21  ( .A1(cv_d[140]), .A2(\cv_reg/n230 ), .ZN(\cv_reg/N143 ) );
  AND2_X1 \cv_reg/U13  ( .A1(cv_d[139]), .A2(\cv_reg/n230 ), .ZN(\cv_reg/N142 ) );
  AND2_X1 \cv_reg/U3  ( .A1(cv_d[138]), .A2(\cv_reg/n230 ), .ZN(\cv_reg/N141 )
         );
  AND2_X2 \cv_reg/U145  ( .A1(cv_d[112]), .A2(\cv_reg/n310 ), .ZN(
        \cv_reg/N115 ) );
  AND2_X2 \cv_reg/U144  ( .A1(cv_d[113]), .A2(\cv_reg/n310 ), .ZN(
        \cv_reg/N116 ) );
  AND2_X2 \cv_reg/U143  ( .A1(cv_d[114]), .A2(\cv_reg/n310 ), .ZN(
        \cv_reg/N117 ) );
  AND2_X2 \cv_reg/U142  ( .A1(cv_d[115]), .A2(\cv_reg/n310 ), .ZN(
        \cv_reg/N118 ) );
  AND2_X2 \cv_reg/U141  ( .A1(cv_d[116]), .A2(\cv_reg/n310 ), .ZN(
        \cv_reg/N119 ) );
  AND2_X2 \cv_reg/U139  ( .A1(cv_d[117]), .A2(\cv_reg/n310 ), .ZN(
        \cv_reg/N120 ) );
  AND2_X2 \cv_reg/U138  ( .A1(cv_d[118]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N121 ) );
  AND2_X2 \cv_reg/U137  ( .A1(cv_d[119]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N122 ) );
  AND2_X2 \cv_reg/U136  ( .A1(cv_d[120]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N123 ) );
  AND2_X2 \cv_reg/U135  ( .A1(cv_d[121]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N124 ) );
  AND2_X2 \cv_reg/U134  ( .A1(cv_d[122]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N125 ) );
  AND2_X2 \cv_reg/U133  ( .A1(cv_d[123]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N126 ) );
  AND2_X2 \cv_reg/U132  ( .A1(cv_d[124]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N127 ) );
  AND2_X2 \cv_reg/U131  ( .A1(cv_d[125]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N128 ) );
  AND2_X2 \cv_reg/U130  ( .A1(cv_d[126]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N129 ) );
  AND2_X2 \cv_reg/U128  ( .A1(cv_d[127]), .A2(\cv_reg/n300 ), .ZN(
        \cv_reg/N130 ) );
  AND2_X2 \cv_reg/U104  ( .A1(cv_d[149]), .A2(\cv_reg/n290 ), .ZN(
        \cv_reg/N152 ) );
  AND2_X2 \cv_reg/U103  ( .A1(cv_d[150]), .A2(\cv_reg/n290 ), .ZN(
        \cv_reg/N153 ) );
  AND2_X2 \cv_reg/U100  ( .A1(cv_d[153]), .A2(\cv_reg/n290 ), .ZN(
        \cv_reg/N156 ) );
  AND2_X2 \cv_reg/U99  ( .A1(cv_d[154]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N157 ) );
  AND2_X2 \cv_reg/U98  ( .A1(cv_d[155]), .A2(\cv_reg/n290 ), .ZN(\cv_reg/N158 ) );
  AND2_X2 \cv_reg/U94  ( .A1(cv_d[158]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N161 ) );
  AND2_X2 \cv_reg/U93  ( .A1(cv_d[159]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N162 ) );
  AND2_X2 \cv_reg/U90  ( .A1(cv_d[16]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N19 )
         );
  AND2_X2 \cv_reg/U89  ( .A1(cv_d[17]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N20 )
         );
  AND2_X2 \cv_reg/U88  ( .A1(cv_d[18]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N21 )
         );
  AND2_X2 \cv_reg/U87  ( .A1(cv_d[19]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N22 )
         );
  AND2_X2 \cv_reg/U86  ( .A1(cv_d[20]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N23 )
         );
  AND2_X2 \cv_reg/U85  ( .A1(cv_d[21]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N24 )
         );
  AND2_X2 \cv_reg/U84  ( .A1(cv_d[22]), .A2(\cv_reg/n280 ), .ZN(\cv_reg/N25 )
         );
  AND2_X2 \cv_reg/U83  ( .A1(cv_d[23]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N26 )
         );
  AND2_X2 \cv_reg/U82  ( .A1(cv_d[24]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N27 )
         );
  AND2_X2 \cv_reg/U81  ( .A1(cv_d[25]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N28 )
         );
  AND2_X2 \cv_reg/U80  ( .A1(cv_d[26]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N29 )
         );
  AND2_X2 \cv_reg/U78  ( .A1(cv_d[27]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N30 )
         );
  AND2_X2 \cv_reg/U77  ( .A1(cv_d[28]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N31 )
         );
  AND2_X2 \cv_reg/U76  ( .A1(cv_d[29]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N32 )
         );
  AND2_X2 \cv_reg/U75  ( .A1(cv_d[30]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N33 )
         );
  AND2_X2 \cv_reg/U74  ( .A1(cv_d[31]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N34 )
         );
  AND2_X2 \cv_reg/U55  ( .A1(cv_d[48]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N51 )
         );
  AND2_X2 \cv_reg/U54  ( .A1(cv_d[49]), .A2(\cv_reg/n270 ), .ZN(\cv_reg/N52 )
         );
  AND2_X2 \cv_reg/U53  ( .A1(cv_d[50]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N53 )
         );
  AND2_X2 \cv_reg/U52  ( .A1(cv_d[51]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N54 )
         );
  AND2_X2 \cv_reg/U51  ( .A1(cv_d[52]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N55 )
         );
  AND2_X2 \cv_reg/U50  ( .A1(cv_d[53]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N56 )
         );
  AND2_X2 \cv_reg/U49  ( .A1(cv_d[54]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N57 )
         );
  AND2_X2 \cv_reg/U48  ( .A1(cv_d[55]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N58 )
         );
  AND2_X2 \cv_reg/U47  ( .A1(cv_d[56]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N59 )
         );
  AND2_X2 \cv_reg/U45  ( .A1(cv_d[57]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N60 )
         );
  AND2_X2 \cv_reg/U44  ( .A1(cv_d[58]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N61 )
         );
  AND2_X2 \cv_reg/U43  ( .A1(cv_d[59]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N62 )
         );
  AND2_X2 \cv_reg/U42  ( .A1(cv_d[60]), .A2(\cv_reg/n260 ), .ZN(\cv_reg/N63 )
         );
  AND2_X2 \cv_reg/U41  ( .A1(cv_d[61]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N64 )
         );
  AND2_X2 \cv_reg/U40  ( .A1(cv_d[62]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N65 )
         );
  AND2_X2 \cv_reg/U39  ( .A1(cv_d[63]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N66 )
         );
  AND2_X2 \cv_reg/U20  ( .A1(cv_d[80]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N83 )
         );
  AND2_X2 \cv_reg/U19  ( .A1(cv_d[81]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N84 )
         );
  AND2_X2 \cv_reg/U18  ( .A1(cv_d[82]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N85 )
         );
  AND2_X2 \cv_reg/U17  ( .A1(cv_d[83]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N86 )
         );
  AND2_X2 \cv_reg/U16  ( .A1(cv_d[84]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N87 )
         );
  AND2_X2 \cv_reg/U15  ( .A1(cv_d[85]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N88 )
         );
  AND2_X2 \cv_reg/U14  ( .A1(cv_d[86]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N89 )
         );
  AND2_X2 \cv_reg/U12  ( .A1(cv_d[87]), .A2(\cv_reg/n250 ), .ZN(\cv_reg/N90 )
         );
  AND2_X2 \cv_reg/U11  ( .A1(cv_d[88]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N91 )
         );
  AND2_X2 \cv_reg/U10  ( .A1(cv_d[89]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N92 )
         );
  AND2_X2 \cv_reg/U9  ( .A1(cv_d[90]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N93 )
         );
  AND2_X2 \cv_reg/U8  ( .A1(cv_d[91]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N94 )
         );
  AND2_X2 \cv_reg/U7  ( .A1(cv_d[92]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N95 )
         );
  AND2_X2 \cv_reg/U6  ( .A1(cv_d[93]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N96 )
         );
  AND2_X2 \cv_reg/U5  ( .A1(cv_d[94]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N97 )
         );
  AND2_X2 \cv_reg/U4  ( .A1(cv_d[95]), .A2(\cv_reg/n240 ), .ZN(\cv_reg/N98 )
         );
  DFF_X2 \cv_reg/q_reg_0_  ( .D(\cv_reg/N3 ), .CK(clk), .Q(cv_q[0]), .QN() );
  DFF_X2 \cv_reg/q_reg_1_  ( .D(\cv_reg/N4 ), .CK(clk), .Q(cv_q[1]), .QN() );
  DFF_X2 \cv_reg/q_reg_2_  ( .D(\cv_reg/N5 ), .CK(clk), .Q(cv_q[2]), .QN() );
  DFF_X2 \cv_reg/q_reg_3_  ( .D(\cv_reg/N6 ), .CK(clk), .Q(cv_q[3]), .QN() );
  DFF_X2 \cv_reg/q_reg_4_  ( .D(\cv_reg/N7 ), .CK(clk), .Q(cv_q[4]), .QN() );
  DFF_X2 \cv_reg/q_reg_5_  ( .D(\cv_reg/N8 ), .CK(clk), .Q(cv_q[5]), .QN() );
  DFF_X2 \cv_reg/q_reg_6_  ( .D(\cv_reg/N9 ), .CK(clk), .Q(cv_q[6]), .QN() );
  DFF_X2 \cv_reg/q_reg_7_  ( .D(\cv_reg/N10 ), .CK(clk), .Q(cv_q[7]), .QN() );
  DFF_X2 \cv_reg/q_reg_8_  ( .D(\cv_reg/N11 ), .CK(clk), .Q(cv_q[8]), .QN() );
  DFF_X2 \cv_reg/q_reg_9_  ( .D(\cv_reg/N12 ), .CK(clk), .Q(cv_q[9]), .QN() );
  DFF_X2 \cv_reg/q_reg_10_  ( .D(\cv_reg/N13 ), .CK(clk), .Q(cv_q[10]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_11_  ( .D(\cv_reg/N14 ), .CK(clk), .Q(cv_q[11]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_12_  ( .D(\cv_reg/N15 ), .CK(clk), .Q(cv_q[12]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_13_  ( .D(\cv_reg/N16 ), .CK(clk), .Q(cv_q[13]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_14_  ( .D(\cv_reg/N17 ), .CK(clk), .Q(cv_q[14]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_15_  ( .D(\cv_reg/N18 ), .CK(clk), .Q(cv_q[15]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_16_  ( .D(\cv_reg/N19 ), .CK(clk), .Q(cv_q[16]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_17_  ( .D(\cv_reg/N20 ), .CK(clk), .Q(cv_q[17]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_18_  ( .D(\cv_reg/N21 ), .CK(clk), .Q(cv_q[18]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_19_  ( .D(\cv_reg/N22 ), .CK(clk), .Q(cv_q[19]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_20_  ( .D(\cv_reg/N23 ), .CK(clk), .Q(cv_q[20]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_21_  ( .D(\cv_reg/N24 ), .CK(clk), .Q(cv_q[21]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_22_  ( .D(\cv_reg/N25 ), .CK(clk), .Q(cv_q[22]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_23_  ( .D(\cv_reg/N26 ), .CK(clk), .Q(cv_q[23]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_24_  ( .D(\cv_reg/N27 ), .CK(clk), .Q(cv_q[24]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_25_  ( .D(\cv_reg/N28 ), .CK(clk), .Q(cv_q[25]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_26_  ( .D(\cv_reg/N29 ), .CK(clk), .Q(cv_q[26]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_27_  ( .D(\cv_reg/N30 ), .CK(clk), .Q(cv_q[27]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_28_  ( .D(\cv_reg/N31 ), .CK(clk), .Q(cv_q[28]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_29_  ( .D(\cv_reg/N32 ), .CK(clk), .Q(cv_q[29]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_30_  ( .D(\cv_reg/N33 ), .CK(clk), .Q(cv_q[30]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_31_  ( .D(\cv_reg/N34 ), .CK(clk), .Q(cv_q[31]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_32_  ( .D(\cv_reg/N35 ), .CK(clk), .Q(cv_q[32]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_33_  ( .D(\cv_reg/N36 ), .CK(clk), .Q(cv_q[33]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_34_  ( .D(\cv_reg/N37 ), .CK(clk), .Q(cv_q[34]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_35_  ( .D(\cv_reg/N38 ), .CK(clk), .Q(cv_q[35]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_36_  ( .D(\cv_reg/N39 ), .CK(clk), .Q(cv_q[36]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_37_  ( .D(\cv_reg/N40 ), .CK(clk), .Q(cv_q[37]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_38_  ( .D(\cv_reg/N41 ), .CK(clk), .Q(cv_q[38]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_39_  ( .D(\cv_reg/N42 ), .CK(clk), .Q(cv_q[39]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_40_  ( .D(\cv_reg/N43 ), .CK(clk), .Q(cv_q[40]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_41_  ( .D(\cv_reg/N44 ), .CK(clk), .Q(cv_q[41]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_42_  ( .D(\cv_reg/N45 ), .CK(clk), .Q(cv_q[42]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_43_  ( .D(\cv_reg/N46 ), .CK(clk), .Q(cv_q[43]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_44_  ( .D(\cv_reg/N47 ), .CK(clk), .Q(cv_q[44]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_45_  ( .D(\cv_reg/N48 ), .CK(clk), .Q(cv_q[45]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_46_  ( .D(\cv_reg/N49 ), .CK(clk), .Q(cv_q[46]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_47_  ( .D(\cv_reg/N50 ), .CK(clk), .Q(cv_q[47]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_48_  ( .D(\cv_reg/N51 ), .CK(clk), .Q(cv_q[48]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_49_  ( .D(\cv_reg/N52 ), .CK(clk), .Q(cv_q[49]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_50_  ( .D(\cv_reg/N53 ), .CK(clk), .Q(cv_q[50]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_51_  ( .D(\cv_reg/N54 ), .CK(clk), .Q(cv_q[51]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_52_  ( .D(\cv_reg/N55 ), .CK(clk), .Q(cv_q[52]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_53_  ( .D(\cv_reg/N56 ), .CK(clk), .Q(cv_q[53]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_54_  ( .D(\cv_reg/N57 ), .CK(clk), .Q(cv_q[54]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_55_  ( .D(\cv_reg/N58 ), .CK(clk), .Q(cv_q[55]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_56_  ( .D(\cv_reg/N59 ), .CK(clk), .Q(cv_q[56]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_57_  ( .D(\cv_reg/N60 ), .CK(clk), .Q(cv_q[57]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_58_  ( .D(\cv_reg/N61 ), .CK(clk), .Q(cv_q[58]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_59_  ( .D(\cv_reg/N62 ), .CK(clk), .Q(cv_q[59]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_60_  ( .D(\cv_reg/N63 ), .CK(clk), .Q(cv_q[60]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_61_  ( .D(\cv_reg/N64 ), .CK(clk), .Q(cv_q[61]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_62_  ( .D(\cv_reg/N65 ), .CK(clk), .Q(cv_q[62]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_63_  ( .D(\cv_reg/N66 ), .CK(clk), .Q(cv_q[63]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_64_  ( .D(\cv_reg/N67 ), .CK(clk), .Q(cv_q[64]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_65_  ( .D(\cv_reg/N68 ), .CK(clk), .Q(cv_q[65]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_66_  ( .D(\cv_reg/N69 ), .CK(clk), .Q(cv_q[66]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_67_  ( .D(\cv_reg/N70 ), .CK(clk), .Q(cv_q[67]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_68_  ( .D(\cv_reg/N71 ), .CK(clk), .Q(cv_q[68]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_69_  ( .D(\cv_reg/N72 ), .CK(clk), .Q(cv_q[69]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_70_  ( .D(\cv_reg/N73 ), .CK(clk), .Q(cv_q[70]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_71_  ( .D(\cv_reg/N74 ), .CK(clk), .Q(cv_q[71]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_72_  ( .D(\cv_reg/N75 ), .CK(clk), .Q(cv_q[72]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_73_  ( .D(\cv_reg/N76 ), .CK(clk), .Q(cv_q[73]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_74_  ( .D(\cv_reg/N77 ), .CK(clk), .Q(cv_q[74]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_75_  ( .D(\cv_reg/N78 ), .CK(clk), .Q(cv_q[75]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_76_  ( .D(\cv_reg/N79 ), .CK(clk), .Q(cv_q[76]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_77_  ( .D(\cv_reg/N80 ), .CK(clk), .Q(cv_q[77]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_78_  ( .D(\cv_reg/N81 ), .CK(clk), .Q(cv_q[78]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_79_  ( .D(\cv_reg/N82 ), .CK(clk), .Q(cv_q[79]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_80_  ( .D(\cv_reg/N83 ), .CK(clk), .Q(cv_q[80]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_81_  ( .D(\cv_reg/N84 ), .CK(clk), .Q(cv_q[81]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_82_  ( .D(\cv_reg/N85 ), .CK(clk), .Q(cv_q[82]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_83_  ( .D(\cv_reg/N86 ), .CK(clk), .Q(cv_q[83]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_84_  ( .D(\cv_reg/N87 ), .CK(clk), .Q(cv_q[84]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_85_  ( .D(\cv_reg/N88 ), .CK(clk), .Q(cv_q[85]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_86_  ( .D(\cv_reg/N89 ), .CK(clk), .Q(cv_q[86]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_87_  ( .D(\cv_reg/N90 ), .CK(clk), .Q(cv_q[87]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_88_  ( .D(\cv_reg/N91 ), .CK(clk), .Q(cv_q[88]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_89_  ( .D(\cv_reg/N92 ), .CK(clk), .Q(cv_q[89]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_90_  ( .D(\cv_reg/N93 ), .CK(clk), .Q(cv_q[90]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_91_  ( .D(\cv_reg/N94 ), .CK(clk), .Q(cv_q[91]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_92_  ( .D(\cv_reg/N95 ), .CK(clk), .Q(cv_q[92]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_93_  ( .D(\cv_reg/N96 ), .CK(clk), .Q(cv_q[93]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_94_  ( .D(\cv_reg/N97 ), .CK(clk), .Q(cv_q[94]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_95_  ( .D(\cv_reg/N98 ), .CK(clk), .Q(cv_q[95]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_96_  ( .D(\cv_reg/N99 ), .CK(clk), .Q(cv_q[96]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_97_  ( .D(\cv_reg/N100 ), .CK(clk), .Q(cv_q[97]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_98_  ( .D(\cv_reg/N101 ), .CK(clk), .Q(cv_q[98]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_99_  ( .D(\cv_reg/N102 ), .CK(clk), .Q(cv_q[99]), .QN()
         );
  DFF_X2 \cv_reg/q_reg_100_  ( .D(\cv_reg/N103 ), .CK(clk), .Q(cv_q[100]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_101_  ( .D(\cv_reg/N104 ), .CK(clk), .Q(cv_q[101]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_102_  ( .D(\cv_reg/N105 ), .CK(clk), .Q(cv_q[102]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_103_  ( .D(\cv_reg/N106 ), .CK(clk), .Q(cv_q[103]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_104_  ( .D(\cv_reg/N107 ), .CK(clk), .Q(cv_q[104]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_105_  ( .D(\cv_reg/N108 ), .CK(clk), .Q(cv_q[105]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_106_  ( .D(\cv_reg/N109 ), .CK(clk), .Q(cv_q[106]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_107_  ( .D(\cv_reg/N110 ), .CK(clk), .Q(cv_q[107]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_108_  ( .D(\cv_reg/N111 ), .CK(clk), .Q(cv_q[108]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_109_  ( .D(\cv_reg/N112 ), .CK(clk), .Q(cv_q[109]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_110_  ( .D(\cv_reg/N113 ), .CK(clk), .Q(cv_q[110]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_111_  ( .D(\cv_reg/N114 ), .CK(clk), .Q(cv_q[111]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_112_  ( .D(\cv_reg/N115 ), .CK(clk), .Q(cv_q[112]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_113_  ( .D(\cv_reg/N116 ), .CK(clk), .Q(cv_q[113]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_114_  ( .D(\cv_reg/N117 ), .CK(clk), .Q(cv_q[114]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_115_  ( .D(\cv_reg/N118 ), .CK(clk), .Q(cv_q[115]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_116_  ( .D(\cv_reg/N119 ), .CK(clk), .Q(cv_q[116]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_117_  ( .D(\cv_reg/N120 ), .CK(clk), .Q(cv_q[117]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_118_  ( .D(\cv_reg/N121 ), .CK(clk), .Q(cv_q[118]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_119_  ( .D(\cv_reg/N122 ), .CK(clk), .Q(cv_q[119]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_120_  ( .D(\cv_reg/N123 ), .CK(clk), .Q(cv_q[120]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_121_  ( .D(\cv_reg/N124 ), .CK(clk), .Q(cv_q[121]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_122_  ( .D(\cv_reg/N125 ), .CK(clk), .Q(cv_q[122]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_123_  ( .D(\cv_reg/N126 ), .CK(clk), .Q(cv_q[123]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_124_  ( .D(\cv_reg/N127 ), .CK(clk), .Q(cv_q[124]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_125_  ( .D(\cv_reg/N128 ), .CK(clk), .Q(cv_q[125]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_126_  ( .D(\cv_reg/N129 ), .CK(clk), .Q(cv_q[126]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_127_  ( .D(\cv_reg/N130 ), .CK(clk), .Q(cv_q[127]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_128_  ( .D(\cv_reg/N131 ), .CK(clk), .Q(cv_q[128]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_129_  ( .D(\cv_reg/N132 ), .CK(clk), .Q(cv_q[129]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_130_  ( .D(\cv_reg/N133 ), .CK(clk), .Q(cv_q[130]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_131_  ( .D(\cv_reg/N134 ), .CK(clk), .Q(cv_q[131]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_132_  ( .D(\cv_reg/N135 ), .CK(clk), .Q(cv_q[132]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_133_  ( .D(\cv_reg/N136 ), .CK(clk), .Q(cv_q[133]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_134_  ( .D(\cv_reg/N137 ), .CK(clk), .Q(cv_q[134]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_135_  ( .D(\cv_reg/N138 ), .CK(clk), .Q(cv_q[135]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_136_  ( .D(\cv_reg/N139 ), .CK(clk), .Q(cv_q[136]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_137_  ( .D(\cv_reg/N140 ), .CK(clk), .Q(cv_q[137]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_138_  ( .D(\cv_reg/N141 ), .CK(clk), .Q(cv_q[138]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_139_  ( .D(\cv_reg/N142 ), .CK(clk), .Q(cv_q[139]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_140_  ( .D(\cv_reg/N143 ), .CK(clk), .Q(cv_q[140]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_141_  ( .D(\cv_reg/N144 ), .CK(clk), .Q(cv_q[141]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_142_  ( .D(\cv_reg/N145 ), .CK(clk), .Q(cv_q[142]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_143_  ( .D(\cv_reg/N146 ), .CK(clk), .Q(cv_q[143]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_144_  ( .D(\cv_reg/N147 ), .CK(clk), .Q(cv_q[144]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_145_  ( .D(\cv_reg/N148 ), .CK(clk), .Q(cv_q[145]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_146_  ( .D(\cv_reg/N149 ), .CK(clk), .Q(cv_q[146]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_147_  ( .D(\cv_reg/N150 ), .CK(clk), .Q(cv_q[147]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_148_  ( .D(\cv_reg/N151 ), .CK(clk), .Q(cv_q[148]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_149_  ( .D(\cv_reg/N152 ), .CK(clk), .Q(cv_q[149]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_150_  ( .D(\cv_reg/N153 ), .CK(clk), .Q(cv_q[150]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_151_  ( .D(\cv_reg/N154 ), .CK(clk), .Q(cv_q[151]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_152_  ( .D(\cv_reg/N155 ), .CK(clk), .Q(cv_q[152]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_153_  ( .D(\cv_reg/N156 ), .CK(clk), .Q(cv_q[153]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_154_  ( .D(\cv_reg/N157 ), .CK(clk), .Q(cv_q[154]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_155_  ( .D(\cv_reg/N158 ), .CK(clk), .Q(cv_q[155]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_156_  ( .D(\cv_reg/N159 ), .CK(clk), .Q(cv_q[156]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_157_  ( .D(\cv_reg/N160 ), .CK(clk), .Q(cv_q[157]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_158_  ( .D(\cv_reg/N161 ), .CK(clk), .Q(cv_q[158]), 
        .QN() );
  DFF_X2 \cv_reg/q_reg_159_  ( .D(\cv_reg/N162 ), .CK(clk), .Q(cv_q[159]), 
        .QN() );
  AND2_X2 \rnd_reg/U178  ( .A1(rnd_d[159]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N162 ) );
  AND2_X2 \rnd_reg/U177  ( .A1(rnd_d[158]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N161 ) );
  AND2_X2 \rnd_reg/U176  ( .A1(rnd_d[157]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N160 ) );
  AND2_X2 \rnd_reg/U175  ( .A1(rnd_d[156]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N159 ) );
  AND2_X2 \rnd_reg/U174  ( .A1(rnd_d[154]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N157 ) );
  AND2_X2 \rnd_reg/U173  ( .A1(rnd_d[153]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N156 ) );
  AND2_X2 \rnd_reg/U172  ( .A1(rnd_d[152]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N155 ) );
  AND2_X2 \rnd_reg/U171  ( .A1(rnd_d[151]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N154 ) );
  AND2_X2 \rnd_reg/U170  ( .A1(rnd_d[149]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N152 ) );
  AND2_X2 \rnd_reg/U169  ( .A1(rnd_d[148]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N151 ) );
  AND2_X2 \rnd_reg/U168  ( .A1(rnd_d[147]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N150 ) );
  AND2_X2 \rnd_reg/U167  ( .A1(rnd_d[146]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N149 ) );
  AND2_X2 \rnd_reg/U166  ( .A1(rnd_d[145]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N148 ) );
  AND2_X2 \rnd_reg/U165  ( .A1(rnd_d[144]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N147 ) );
  AND2_X2 \rnd_reg/U164  ( .A1(rnd_d[143]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N146 ) );
  AND2_X2 \rnd_reg/U163  ( .A1(rnd_d[142]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N145 ) );
  AND2_X2 \rnd_reg/U162  ( .A1(rnd_d[141]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N144 ) );
  AND2_X2 \rnd_reg/U161  ( .A1(rnd_d[140]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N143 ) );
  AND2_X2 \rnd_reg/U160  ( .A1(rnd_d[139]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N142 ) );
  AND2_X2 \rnd_reg/U159  ( .A1(rnd_d[138]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N141 ) );
  AND2_X2 \rnd_reg/U158  ( .A1(rnd_d[137]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N140 ) );
  AND2_X2 \rnd_reg/U157  ( .A1(rnd_d[136]), .A2(\rnd_reg/n250 ), .ZN(
        \rnd_reg/N139 ) );
  AND2_X2 \rnd_reg/U156  ( .A1(rnd_d[135]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N138 ) );
  AND2_X2 \rnd_reg/U155  ( .A1(rnd_d[134]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N137 ) );
  AND2_X2 \rnd_reg/U154  ( .A1(rnd_d[133]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N136 ) );
  AND2_X2 \rnd_reg/U153  ( .A1(rnd_d[132]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N135 ) );
  AND2_X2 \rnd_reg/U152  ( .A1(rnd_d[131]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N134 ) );
  AND2_X2 \rnd_reg/U151  ( .A1(rnd_d[130]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N133 ) );
  AND2_X2 \rnd_reg/U150  ( .A1(rnd_d[129]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N132 ) );
  AND2_X2 \rnd_reg/U149  ( .A1(rnd_d[128]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N131 ) );
  AND2_X2 \rnd_reg/U148  ( .A1(rnd_d[116]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N119 ) );
  AND2_X2 \rnd_reg/U147  ( .A1(rnd_d[115]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N118 ) );
  AND2_X2 \rnd_reg/U146  ( .A1(rnd_d[114]), .A2(\rnd_reg/n240 ), .ZN(
        \rnd_reg/N117 ) );
  AND2_X2 \rnd_reg/U145  ( .A1(rnd_d[113]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N116 ) );
  AND2_X2 \rnd_reg/U144  ( .A1(rnd_d[112]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N115 ) );
  AND2_X2 \rnd_reg/U143  ( .A1(rnd_d[111]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N114 ) );
  AND2_X2 \rnd_reg/U142  ( .A1(rnd_d[110]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N113 ) );
  AND2_X2 \rnd_reg/U141  ( .A1(rnd_d[109]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N112 ) );
  AND2_X2 \rnd_reg/U140  ( .A1(rnd_d[108]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N111 ) );
  AND2_X2 \rnd_reg/U129  ( .A1(rnd_d[107]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N110 ) );
  AND2_X2 \rnd_reg/U127  ( .A1(rnd_d[106]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N109 ) );
  AND2_X2 \rnd_reg/U126  ( .A1(rnd_d[105]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N108 ) );
  AND2_X2 \rnd_reg/U125  ( .A1(rnd_d[104]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N107 ) );
  AND2_X2 \rnd_reg/U124  ( .A1(rnd_d[103]), .A2(\rnd_reg/n230 ), .ZN(
        \rnd_reg/N106 ) );
  AND2_X2 \rnd_reg/U123  ( .A1(rnd_d[102]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N105 ) );
  AND2_X2 \rnd_reg/U122  ( .A1(rnd_d[101]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N104 ) );
  AND2_X2 \rnd_reg/U121  ( .A1(rnd_d[100]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N103 ) );
  AND2_X2 \rnd_reg/U120  ( .A1(rnd_d[99]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N102 ) );
  AND2_X2 \rnd_reg/U119  ( .A1(rnd_d[98]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N101 ) );
  AND2_X2 \rnd_reg/U118  ( .A1(rnd_d[97]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N100 ) );
  AND2_X2 \rnd_reg/U117  ( .A1(rnd_d[96]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N99 ) );
  AND2_X2 \rnd_reg/U116  ( .A1(rnd_d[83]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N86 ) );
  AND2_X2 \rnd_reg/U115  ( .A1(rnd_d[82]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N85 ) );
  AND2_X2 \rnd_reg/U114  ( .A1(rnd_d[81]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N84 ) );
  AND2_X2 \rnd_reg/U113  ( .A1(rnd_d[80]), .A2(\rnd_reg/n220 ), .ZN(
        \rnd_reg/N83 ) );
  AND2_X2 \rnd_reg/U112  ( .A1(rnd_d[79]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N82 ) );
  AND2_X2 \rnd_reg/U111  ( .A1(rnd_d[78]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N81 ) );
  AND2_X2 \rnd_reg/U110  ( .A1(rnd_d[77]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N80 ) );
  AND2_X2 \rnd_reg/U109  ( .A1(rnd_d[76]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N79 ) );
  AND2_X2 \rnd_reg/U108  ( .A1(rnd_d[75]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N78 ) );
  AND2_X2 \rnd_reg/U107  ( .A1(rnd_d[74]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N77 ) );
  AND2_X2 \rnd_reg/U106  ( .A1(rnd_d[73]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N76 ) );
  AND2_X2 \rnd_reg/U105  ( .A1(rnd_d[72]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N75 ) );
  AND2_X2 \rnd_reg/U104  ( .A1(rnd_d[71]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N74 ) );
  AND2_X2 \rnd_reg/U103  ( .A1(rnd_d[70]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N73 ) );
  AND2_X2 \rnd_reg/U102  ( .A1(rnd_d[69]), .A2(\rnd_reg/n210 ), .ZN(
        \rnd_reg/N72 ) );
  AND2_X2 \rnd_reg/U101  ( .A1(rnd_d[68]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N71 ) );
  AND2_X2 \rnd_reg/U100  ( .A1(rnd_d[67]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N70 ) );
  AND2_X2 \rnd_reg/U99  ( .A1(rnd_d[66]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N69 ) );
  AND2_X2 \rnd_reg/U98  ( .A1(rnd_d[65]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N68 ) );
  AND2_X2 \rnd_reg/U97  ( .A1(rnd_d[64]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N67 ) );
  AND2_X2 \rnd_reg/U96  ( .A1(rnd_d[51]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N54 ) );
  AND2_X2 \rnd_reg/U95  ( .A1(rnd_d[50]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N53 ) );
  AND2_X2 \rnd_reg/U94  ( .A1(rnd_d[49]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N52 ) );
  AND2_X2 \rnd_reg/U93  ( .A1(rnd_d[48]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N51 ) );
  AND2_X2 \rnd_reg/U92  ( .A1(rnd_d[47]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N50 ) );
  AND2_X2 \rnd_reg/U91  ( .A1(rnd_d[46]), .A2(\rnd_reg/n200 ), .ZN(
        \rnd_reg/N49 ) );
  AND2_X2 \rnd_reg/U90  ( .A1(rnd_d[45]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N48 ) );
  AND2_X2 \rnd_reg/U89  ( .A1(rnd_d[44]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N47 ) );
  AND2_X2 \rnd_reg/U88  ( .A1(rnd_d[43]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N46 ) );
  AND2_X2 \rnd_reg/U79  ( .A1(rnd_d[42]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N45 ) );
  AND2_X2 \rnd_reg/U73  ( .A1(rnd_d[41]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N44 ) );
  AND2_X2 \rnd_reg/U72  ( .A1(rnd_d[40]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N43 ) );
  AND2_X2 \rnd_reg/U71  ( .A1(rnd_d[39]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N42 ) );
  AND2_X2 \rnd_reg/U70  ( .A1(rnd_d[38]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N41 ) );
  AND2_X2 \rnd_reg/U69  ( .A1(rnd_d[37]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N40 ) );
  AND2_X2 \rnd_reg/U68  ( .A1(rnd_d[36]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N39 ) );
  AND2_X2 \rnd_reg/U67  ( .A1(rnd_d[35]), .A2(\rnd_reg/n190 ), .ZN(
        \rnd_reg/N38 ) );
  AND2_X2 \rnd_reg/U66  ( .A1(rnd_d[34]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N37 ) );
  AND2_X2 \rnd_reg/U65  ( .A1(rnd_d[33]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N36 ) );
  AND2_X2 \rnd_reg/U64  ( .A1(rnd_d[32]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N35 ) );
  AND2_X2 \rnd_reg/U63  ( .A1(rnd_d[18]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N21 ) );
  AND2_X2 \rnd_reg/U62  ( .A1(rnd_d[17]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N20 ) );
  AND2_X2 \rnd_reg/U61  ( .A1(rnd_d[16]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N19 ) );
  AND2_X2 \rnd_reg/U60  ( .A1(rnd_d[15]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N18 ) );
  AND2_X2 \rnd_reg/U59  ( .A1(rnd_d[14]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N17 ) );
  AND2_X2 \rnd_reg/U58  ( .A1(rnd_d[13]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N16 ) );
  AND2_X2 \rnd_reg/U57  ( .A1(rnd_d[12]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N15 ) );
  AND2_X2 \rnd_reg/U56  ( .A1(rnd_d[11]), .A2(\rnd_reg/n180 ), .ZN(
        \rnd_reg/N14 ) );
  AND2_X2 \rnd_reg/U55  ( .A1(rnd_d[10]), .A2(\rnd_reg/n170 ), .ZN(
        \rnd_reg/N13 ) );
  AND2_X2 \rnd_reg/U54  ( .A1(rnd_d[9]), .A2(\rnd_reg/n170 ), .ZN(
        \rnd_reg/N12 ) );
  AND2_X2 \rnd_reg/U53  ( .A1(rnd_d[8]), .A2(\rnd_reg/n170 ), .ZN(
        \rnd_reg/N11 ) );
  AND2_X2 \rnd_reg/U52  ( .A1(rnd_d[7]), .A2(\rnd_reg/n170 ), .ZN(
        \rnd_reg/N10 ) );
  AND2_X2 \rnd_reg/U46  ( .A1(rnd_d[6]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N9 ) );
  AND2_X2 \rnd_reg/U38  ( .A1(rnd_d[5]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N8 ) );
  AND2_X2 \rnd_reg/U37  ( .A1(rnd_d[4]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N7 ) );
  AND2_X2 \rnd_reg/U36  ( .A1(rnd_d[3]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N6 ) );
  AND2_X2 \rnd_reg/U35  ( .A1(rnd_d[2]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N5 ) );
  AND2_X2 \rnd_reg/U34  ( .A1(rnd_d[1]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N4 ) );
  AND2_X2 \rnd_reg/U33  ( .A1(rnd_d[0]), .A2(\rnd_reg/n170 ), .ZN(\rnd_reg/N3 ) );
  INV_X4 \rnd_reg/U32  ( .A(\rnd_reg/n190 ), .ZN(\rnd_reg/n320 ) );
  INV_X4 \rnd_reg/U31  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n310 ) );
  INV_X4 \rnd_reg/U30  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n220 ) );
  INV_X4 \rnd_reg/U29  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n210 ) );
  INV_X4 \rnd_reg/U28  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n200 ) );
  INV_X4 \rnd_reg/U27  ( .A(n7117), .ZN(\rnd_reg/n190 ) );
  INV_X4 \rnd_reg/U26  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n180 ) );
  INV_X4 \rnd_reg/U25  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n170 ) );
  INV_X4 \rnd_reg/U24  ( .A(n7117), .ZN(\rnd_reg/n260 ) );
  INV_X4 \rnd_reg/U23  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n250 ) );
  INV_X4 \rnd_reg/U22  ( .A(n7117), .ZN(\rnd_reg/n240 ) );
  INV_X4 \rnd_reg/U21  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n300 ) );
  INV_X4 \rnd_reg/U20  ( .A(n7117), .ZN(\rnd_reg/n230 ) );
  INV_X4 \rnd_reg/U19  ( .A(n7117), .ZN(\rnd_reg/n270 ) );
  INV_X4 \rnd_reg/U18  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n280 ) );
  INV_X4 \rnd_reg/U17  ( .A(\rnd_reg/n320 ), .ZN(\rnd_reg/n290 ) );
  AND2_X4 \rnd_reg/U13  ( .A1(rnd_d[155]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N158 ) );
  AND2_X4 \rnd_reg/U3  ( .A1(rnd_d[150]), .A2(\rnd_reg/n260 ), .ZN(
        \rnd_reg/N153 ) );
  DFF_X2 \rnd_reg/q_reg_156_  ( .D(\rnd_reg/N159 ), .CK(clk), .Q(rnd_q[156]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_155_  ( .D(\rnd_reg/N158 ), .CK(clk), .Q(rnd_q[155]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_158_  ( .D(\rnd_reg/N161 ), .CK(clk), .Q(rnd_q[158]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_157_  ( .D(\rnd_reg/N160 ), .CK(clk), .Q(rnd_q[157]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_159_  ( .D(\rnd_reg/N162 ), .CK(clk), .Q(rnd_q[159]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_150_  ( .D(\rnd_reg/N153 ), .CK(clk), .Q(rnd_q[150]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_154_  ( .D(\rnd_reg/N157 ), .CK(clk), .Q(rnd_q[154]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_153_  ( .D(\rnd_reg/N156 ), .CK(clk), .Q(rnd_q[153]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_151_  ( .D(\rnd_reg/N154 ), .CK(clk), .Q(rnd_q[151]), 
        .QN() );
  AND2_X2 \rnd_reg/U139  ( .A1(rnd_d[117]), .A2(\rnd_reg/n310 ), .ZN(
        \rnd_reg/N120 ) );
  AND2_X2 \rnd_reg/U138  ( .A1(rnd_d[118]), .A2(\rnd_reg/n310 ), .ZN(
        \rnd_reg/N121 ) );
  AND2_X2 \rnd_reg/U137  ( .A1(rnd_d[119]), .A2(\rnd_reg/n310 ), .ZN(
        \rnd_reg/N122 ) );
  AND2_X2 \rnd_reg/U136  ( .A1(rnd_d[120]), .A2(\rnd_reg/n310 ), .ZN(
        \rnd_reg/N123 ) );
  AND2_X2 \rnd_reg/U135  ( .A1(rnd_d[121]), .A2(\rnd_reg/n310 ), .ZN(
        \rnd_reg/N124 ) );
  AND2_X2 \rnd_reg/U134  ( .A1(rnd_d[122]), .A2(\rnd_reg/n310 ), .ZN(
        \rnd_reg/N125 ) );
  AND2_X2 \rnd_reg/U133  ( .A1(rnd_d[123]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N126 ) );
  AND2_X2 \rnd_reg/U132  ( .A1(rnd_d[124]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N127 ) );
  AND2_X2 \rnd_reg/U131  ( .A1(rnd_d[125]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N128 ) );
  AND2_X2 \rnd_reg/U130  ( .A1(rnd_d[126]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N129 ) );
  AND2_X2 \rnd_reg/U128  ( .A1(rnd_d[127]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N130 ) );
  AND2_X2 \rnd_reg/U87  ( .A1(rnd_d[19]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N22 ) );
  AND2_X2 \rnd_reg/U86  ( .A1(rnd_d[20]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N23 ) );
  AND2_X2 \rnd_reg/U85  ( .A1(rnd_d[21]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N24 ) );
  AND2_X2 \rnd_reg/U84  ( .A1(rnd_d[22]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N25 ) );
  AND2_X2 \rnd_reg/U83  ( .A1(rnd_d[23]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N26 ) );
  AND2_X2 \rnd_reg/U82  ( .A1(rnd_d[24]), .A2(\rnd_reg/n300 ), .ZN(
        \rnd_reg/N27 ) );
  AND2_X2 \rnd_reg/U81  ( .A1(rnd_d[25]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N28 ) );
  AND2_X2 \rnd_reg/U80  ( .A1(rnd_d[26]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N29 ) );
  AND2_X2 \rnd_reg/U78  ( .A1(rnd_d[27]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N30 ) );
  AND2_X2 \rnd_reg/U77  ( .A1(rnd_d[28]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N31 ) );
  AND2_X2 \rnd_reg/U76  ( .A1(rnd_d[29]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N32 ) );
  AND2_X2 \rnd_reg/U75  ( .A1(rnd_d[30]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N33 ) );
  AND2_X2 \rnd_reg/U74  ( .A1(rnd_d[31]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N34 ) );
  AND2_X2 \rnd_reg/U51  ( .A1(rnd_d[52]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N55 ) );
  AND2_X2 \rnd_reg/U50  ( .A1(rnd_d[53]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N56 ) );
  AND2_X2 \rnd_reg/U49  ( .A1(rnd_d[54]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N57 ) );
  AND2_X2 \rnd_reg/U48  ( .A1(rnd_d[55]), .A2(\rnd_reg/n290 ), .ZN(
        \rnd_reg/N58 ) );
  AND2_X2 \rnd_reg/U47  ( .A1(rnd_d[56]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N59 ) );
  AND2_X2 \rnd_reg/U45  ( .A1(rnd_d[57]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N60 ) );
  AND2_X2 \rnd_reg/U44  ( .A1(rnd_d[58]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N61 ) );
  AND2_X2 \rnd_reg/U43  ( .A1(rnd_d[59]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N62 ) );
  AND2_X2 \rnd_reg/U42  ( .A1(rnd_d[60]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N63 ) );
  AND2_X2 \rnd_reg/U41  ( .A1(rnd_d[61]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N64 ) );
  AND2_X2 \rnd_reg/U40  ( .A1(rnd_d[62]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N65 ) );
  AND2_X2 \rnd_reg/U39  ( .A1(rnd_d[63]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N66 ) );
  AND2_X2 \rnd_reg/U16  ( .A1(rnd_d[84]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N87 ) );
  AND2_X2 \rnd_reg/U15  ( .A1(rnd_d[85]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N88 ) );
  AND2_X2 \rnd_reg/U14  ( .A1(rnd_d[86]), .A2(\rnd_reg/n280 ), .ZN(
        \rnd_reg/N89 ) );
  AND2_X2 \rnd_reg/U12  ( .A1(rnd_d[87]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N90 ) );
  AND2_X2 \rnd_reg/U11  ( .A1(rnd_d[88]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N91 ) );
  AND2_X2 \rnd_reg/U10  ( .A1(rnd_d[89]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N92 ) );
  AND2_X2 \rnd_reg/U9  ( .A1(rnd_d[90]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N93 ) );
  AND2_X2 \rnd_reg/U8  ( .A1(rnd_d[91]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N94 ) );
  AND2_X2 \rnd_reg/U7  ( .A1(rnd_d[92]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N95 ) );
  AND2_X2 \rnd_reg/U6  ( .A1(rnd_d[93]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N96 ) );
  AND2_X2 \rnd_reg/U5  ( .A1(rnd_d[94]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N97 ) );
  AND2_X2 \rnd_reg/U4  ( .A1(rnd_d[95]), .A2(\rnd_reg/n270 ), .ZN(
        \rnd_reg/N98 ) );
  DFF_X2 \rnd_reg/q_reg_0_  ( .D(\rnd_reg/N3 ), .CK(clk), .Q(rnd_q[0]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_1_  ( .D(\rnd_reg/N4 ), .CK(clk), .Q(rnd_q[1]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_2_  ( .D(\rnd_reg/N5 ), .CK(clk), .Q(rnd_q[2]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_3_  ( .D(\rnd_reg/N6 ), .CK(clk), .Q(rnd_q[3]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_4_  ( .D(\rnd_reg/N7 ), .CK(clk), .Q(rnd_q[4]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_5_  ( .D(\rnd_reg/N8 ), .CK(clk), .Q(rnd_q[5]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_6_  ( .D(\rnd_reg/N9 ), .CK(clk), .Q(rnd_q[6]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_7_  ( .D(\rnd_reg/N10 ), .CK(clk), .Q(rnd_q[7]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_8_  ( .D(\rnd_reg/N11 ), .CK(clk), .Q(rnd_q[8]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_9_  ( .D(\rnd_reg/N12 ), .CK(clk), .Q(rnd_q[9]), .QN()
         );
  DFF_X2 \rnd_reg/q_reg_10_  ( .D(\rnd_reg/N13 ), .CK(clk), .Q(rnd_q[10]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_11_  ( .D(\rnd_reg/N14 ), .CK(clk), .Q(rnd_q[11]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_12_  ( .D(\rnd_reg/N15 ), .CK(clk), .Q(rnd_q[12]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_13_  ( .D(\rnd_reg/N16 ), .CK(clk), .Q(rnd_q[13]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_14_  ( .D(\rnd_reg/N17 ), .CK(clk), .Q(rnd_q[14]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_15_  ( .D(\rnd_reg/N18 ), .CK(clk), .Q(rnd_q[15]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_16_  ( .D(\rnd_reg/N19 ), .CK(clk), .Q(rnd_q[16]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_17_  ( .D(\rnd_reg/N20 ), .CK(clk), .Q(rnd_q[17]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_18_  ( .D(\rnd_reg/N21 ), .CK(clk), .Q(rnd_q[18]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_19_  ( .D(\rnd_reg/N22 ), .CK(clk), .Q(rnd_q[19]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_20_  ( .D(\rnd_reg/N23 ), .CK(clk), .Q(rnd_q[20]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_21_  ( .D(\rnd_reg/N24 ), .CK(clk), .Q(rnd_q[21]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_22_  ( .D(\rnd_reg/N25 ), .CK(clk), .Q(rnd_q[22]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_23_  ( .D(\rnd_reg/N26 ), .CK(clk), .Q(rnd_q[23]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_24_  ( .D(\rnd_reg/N27 ), .CK(clk), .Q(rnd_q[24]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_25_  ( .D(\rnd_reg/N28 ), .CK(clk), .Q(rnd_q[25]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_26_  ( .D(\rnd_reg/N29 ), .CK(clk), .Q(rnd_q[26]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_27_  ( .D(\rnd_reg/N30 ), .CK(clk), .Q(rnd_q[27]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_28_  ( .D(\rnd_reg/N31 ), .CK(clk), .Q(rnd_q[28]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_29_  ( .D(\rnd_reg/N32 ), .CK(clk), .Q(rnd_q[29]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_30_  ( .D(\rnd_reg/N33 ), .CK(clk), .Q(rnd_q[30]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_31_  ( .D(\rnd_reg/N34 ), .CK(clk), .Q(rnd_q[31]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_32_  ( .D(\rnd_reg/N35 ), .CK(clk), .Q(rnd_q[32]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_33_  ( .D(\rnd_reg/N36 ), .CK(clk), .Q(rnd_q[33]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_34_  ( .D(\rnd_reg/N37 ), .CK(clk), .Q(rnd_q[34]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_35_  ( .D(\rnd_reg/N38 ), .CK(clk), .Q(rnd_q[35]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_36_  ( .D(\rnd_reg/N39 ), .CK(clk), .Q(rnd_q[36]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_37_  ( .D(\rnd_reg/N40 ), .CK(clk), .Q(rnd_q[37]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_38_  ( .D(\rnd_reg/N41 ), .CK(clk), .Q(rnd_q[38]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_39_  ( .D(\rnd_reg/N42 ), .CK(clk), .Q(rnd_q[39]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_40_  ( .D(\rnd_reg/N43 ), .CK(clk), .Q(rnd_q[40]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_41_  ( .D(\rnd_reg/N44 ), .CK(clk), .Q(rnd_q[41]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_42_  ( .D(\rnd_reg/N45 ), .CK(clk), .Q(rnd_q[42]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_43_  ( .D(\rnd_reg/N46 ), .CK(clk), .Q(rnd_q[43]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_44_  ( .D(\rnd_reg/N47 ), .CK(clk), .Q(rnd_q[44]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_45_  ( .D(\rnd_reg/N48 ), .CK(clk), .Q(rnd_q[45]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_46_  ( .D(\rnd_reg/N49 ), .CK(clk), .Q(rnd_q[46]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_47_  ( .D(\rnd_reg/N50 ), .CK(clk), .Q(rnd_q[47]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_48_  ( .D(\rnd_reg/N51 ), .CK(clk), .Q(rnd_q[48]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_49_  ( .D(\rnd_reg/N52 ), .CK(clk), .Q(rnd_q[49]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_50_  ( .D(\rnd_reg/N53 ), .CK(clk), .Q(rnd_q[50]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_51_  ( .D(\rnd_reg/N54 ), .CK(clk), .Q(rnd_q[51]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_52_  ( .D(\rnd_reg/N55 ), .CK(clk), .Q(rnd_q[52]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_53_  ( .D(\rnd_reg/N56 ), .CK(clk), .Q(rnd_q[53]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_54_  ( .D(\rnd_reg/N57 ), .CK(clk), .Q(rnd_q[54]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_55_  ( .D(\rnd_reg/N58 ), .CK(clk), .Q(rnd_q[55]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_56_  ( .D(\rnd_reg/N59 ), .CK(clk), .Q(rnd_q[56]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_57_  ( .D(\rnd_reg/N60 ), .CK(clk), .Q(rnd_q[57]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_58_  ( .D(\rnd_reg/N61 ), .CK(clk), .Q(rnd_q[58]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_59_  ( .D(\rnd_reg/N62 ), .CK(clk), .Q(rnd_q[59]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_60_  ( .D(\rnd_reg/N63 ), .CK(clk), .Q(rnd_q[60]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_61_  ( .D(\rnd_reg/N64 ), .CK(clk), .Q(rnd_q[61]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_62_  ( .D(\rnd_reg/N65 ), .CK(clk), .Q(rnd_q[62]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_63_  ( .D(\rnd_reg/N66 ), .CK(clk), .Q(rnd_q[63]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_64_  ( .D(\rnd_reg/N67 ), .CK(clk), .Q(rnd_q[64]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_65_  ( .D(\rnd_reg/N68 ), .CK(clk), .Q(rnd_q[65]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_66_  ( .D(\rnd_reg/N69 ), .CK(clk), .Q(rnd_q[66]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_67_  ( .D(\rnd_reg/N70 ), .CK(clk), .Q(rnd_q[67]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_68_  ( .D(\rnd_reg/N71 ), .CK(clk), .Q(rnd_q[68]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_69_  ( .D(\rnd_reg/N72 ), .CK(clk), .Q(rnd_q[69]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_70_  ( .D(\rnd_reg/N73 ), .CK(clk), .Q(rnd_q[70]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_71_  ( .D(\rnd_reg/N74 ), .CK(clk), .Q(rnd_q[71]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_72_  ( .D(\rnd_reg/N75 ), .CK(clk), .Q(rnd_q[72]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_73_  ( .D(\rnd_reg/N76 ), .CK(clk), .Q(rnd_q[73]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_74_  ( .D(\rnd_reg/N77 ), .CK(clk), .Q(rnd_q[74]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_75_  ( .D(\rnd_reg/N78 ), .CK(clk), .Q(rnd_q[75]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_76_  ( .D(\rnd_reg/N79 ), .CK(clk), .Q(rnd_q[76]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_77_  ( .D(\rnd_reg/N80 ), .CK(clk), .Q(rnd_q[77]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_78_  ( .D(\rnd_reg/N81 ), .CK(clk), .Q(rnd_q[78]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_79_  ( .D(\rnd_reg/N82 ), .CK(clk), .Q(rnd_q[79]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_80_  ( .D(\rnd_reg/N83 ), .CK(clk), .Q(rnd_q[80]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_81_  ( .D(\rnd_reg/N84 ), .CK(clk), .Q(rnd_q[81]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_82_  ( .D(\rnd_reg/N85 ), .CK(clk), .Q(rnd_q[82]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_83_  ( .D(\rnd_reg/N86 ), .CK(clk), .Q(rnd_q[83]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_84_  ( .D(\rnd_reg/N87 ), .CK(clk), .Q(rnd_q[84]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_85_  ( .D(\rnd_reg/N88 ), .CK(clk), .Q(rnd_q[85]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_86_  ( .D(\rnd_reg/N89 ), .CK(clk), .Q(rnd_q[86]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_87_  ( .D(\rnd_reg/N90 ), .CK(clk), .Q(rnd_q[87]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_88_  ( .D(\rnd_reg/N91 ), .CK(clk), .Q(rnd_q[88]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_89_  ( .D(\rnd_reg/N92 ), .CK(clk), .Q(rnd_q[89]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_90_  ( .D(\rnd_reg/N93 ), .CK(clk), .Q(rnd_q[90]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_91_  ( .D(\rnd_reg/N94 ), .CK(clk), .Q(rnd_q[91]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_92_  ( .D(\rnd_reg/N95 ), .CK(clk), .Q(rnd_q[92]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_93_  ( .D(\rnd_reg/N96 ), .CK(clk), .Q(rnd_q[93]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_94_  ( .D(\rnd_reg/N97 ), .CK(clk), .Q(rnd_q[94]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_95_  ( .D(\rnd_reg/N98 ), .CK(clk), .Q(rnd_q[95]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_96_  ( .D(\rnd_reg/N99 ), .CK(clk), .Q(rnd_q[96]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_97_  ( .D(\rnd_reg/N100 ), .CK(clk), .Q(rnd_q[97]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_98_  ( .D(\rnd_reg/N101 ), .CK(clk), .Q(rnd_q[98]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_99_  ( .D(\rnd_reg/N102 ), .CK(clk), .Q(rnd_q[99]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_100_  ( .D(\rnd_reg/N103 ), .CK(clk), .Q(rnd_q[100]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_101_  ( .D(\rnd_reg/N104 ), .CK(clk), .Q(rnd_q[101]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_102_  ( .D(\rnd_reg/N105 ), .CK(clk), .Q(rnd_q[102]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_103_  ( .D(\rnd_reg/N106 ), .CK(clk), .Q(rnd_q[103]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_104_  ( .D(\rnd_reg/N107 ), .CK(clk), .Q(rnd_q[104]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_105_  ( .D(\rnd_reg/N108 ), .CK(clk), .Q(rnd_q[105]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_106_  ( .D(\rnd_reg/N109 ), .CK(clk), .Q(rnd_q[106]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_107_  ( .D(\rnd_reg/N110 ), .CK(clk), .Q(rnd_q[107]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_108_  ( .D(\rnd_reg/N111 ), .CK(clk), .Q(rnd_q[108]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_109_  ( .D(\rnd_reg/N112 ), .CK(clk), .Q(rnd_q[109]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_110_  ( .D(\rnd_reg/N113 ), .CK(clk), .Q(rnd_q[110]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_111_  ( .D(\rnd_reg/N114 ), .CK(clk), .Q(rnd_q[111]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_112_  ( .D(\rnd_reg/N115 ), .CK(clk), .Q(rnd_q[112]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_113_  ( .D(\rnd_reg/N116 ), .CK(clk), .Q(rnd_q[113]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_114_  ( .D(\rnd_reg/N117 ), .CK(clk), .Q(rnd_q[114]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_115_  ( .D(\rnd_reg/N118 ), .CK(clk), .Q(rnd_q[115]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_116_  ( .D(\rnd_reg/N119 ), .CK(clk), .Q(rnd_q[116]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_117_  ( .D(\rnd_reg/N120 ), .CK(clk), .Q(rnd_q[117]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_118_  ( .D(\rnd_reg/N121 ), .CK(clk), .Q(rnd_q[118]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_119_  ( .D(\rnd_reg/N122 ), .CK(clk), .Q(rnd_q[119]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_120_  ( .D(\rnd_reg/N123 ), .CK(clk), .Q(rnd_q[120]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_121_  ( .D(\rnd_reg/N124 ), .CK(clk), .Q(rnd_q[121]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_122_  ( .D(\rnd_reg/N125 ), .CK(clk), .Q(rnd_q[122]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_123_  ( .D(\rnd_reg/N126 ), .CK(clk), .Q(rnd_q[123]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_124_  ( .D(\rnd_reg/N127 ), .CK(clk), .Q(rnd_q[124]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_125_  ( .D(\rnd_reg/N128 ), .CK(clk), .Q(rnd_q[125]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_126_  ( .D(\rnd_reg/N129 ), .CK(clk), .Q(rnd_q[126]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_127_  ( .D(\rnd_reg/N130 ), .CK(clk), .Q(rnd_q[127]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_128_  ( .D(\rnd_reg/N131 ), .CK(clk), .Q(rnd_q[128]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_129_  ( .D(\rnd_reg/N132 ), .CK(clk), .Q(rnd_q[129]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_130_  ( .D(\rnd_reg/N133 ), .CK(clk), .Q(rnd_q[130]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_131_  ( .D(\rnd_reg/N134 ), .CK(clk), .Q(rnd_q[131]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_132_  ( .D(\rnd_reg/N135 ), .CK(clk), .Q(rnd_q[132]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_133_  ( .D(\rnd_reg/N136 ), .CK(clk), .Q(rnd_q[133]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_134_  ( .D(\rnd_reg/N137 ), .CK(clk), .Q(rnd_q[134]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_135_  ( .D(\rnd_reg/N138 ), .CK(clk), .Q(rnd_q[135]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_136_  ( .D(\rnd_reg/N139 ), .CK(clk), .Q(rnd_q[136]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_137_  ( .D(\rnd_reg/N140 ), .CK(clk), .Q(rnd_q[137]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_138_  ( .D(\rnd_reg/N141 ), .CK(clk), .Q(rnd_q[138]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_139_  ( .D(\rnd_reg/N142 ), .CK(clk), .Q(rnd_q[139]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_140_  ( .D(\rnd_reg/N143 ), .CK(clk), .Q(rnd_q[140]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_141_  ( .D(\rnd_reg/N144 ), .CK(clk), .Q(rnd_q[141]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_142_  ( .D(\rnd_reg/N145 ), .CK(clk), .Q(rnd_q[142]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_143_  ( .D(\rnd_reg/N146 ), .CK(clk), .Q(rnd_q[143]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_144_  ( .D(\rnd_reg/N147 ), .CK(clk), .Q(rnd_q[144]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_145_  ( .D(\rnd_reg/N148 ), .CK(clk), .Q(rnd_q[145]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_146_  ( .D(\rnd_reg/N149 ), .CK(clk), .Q(rnd_q[146]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_147_  ( .D(\rnd_reg/N150 ), .CK(clk), .Q(rnd_q[147]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_148_  ( .D(\rnd_reg/N151 ), .CK(clk), .Q(rnd_q[148]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_149_  ( .D(\rnd_reg/N152 ), .CK(clk), .Q(rnd_q[149]), 
        .QN() );
  DFF_X2 \rnd_reg/q_reg_152_  ( .D(\rnd_reg/N155 ), .CK(clk), .Q(rnd_q[152]), 
        .QN() );
  AND2_X2 \cv_next_reg/U178  ( .A1(cv_next_d[159]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N162 ) );
  AND2_X2 \cv_next_reg/U177  ( .A1(cv_next_d[158]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N161 ) );
  AND2_X2 \cv_next_reg/U176  ( .A1(cv_next_d[157]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N160 ) );
  AND2_X2 \cv_next_reg/U175  ( .A1(cv_next_d[156]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N159 ) );
  AND2_X2 \cv_next_reg/U174  ( .A1(cv_next_d[155]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N158 ) );
  AND2_X2 \cv_next_reg/U173  ( .A1(cv_next_d[154]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N157 ) );
  AND2_X2 \cv_next_reg/U172  ( .A1(cv_next_d[153]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N156 ) );
  AND2_X2 \cv_next_reg/U171  ( .A1(cv_next_d[152]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N155 ) );
  AND2_X2 \cv_next_reg/U170  ( .A1(cv_next_d[151]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N154 ) );
  AND2_X2 \cv_next_reg/U169  ( .A1(cv_next_d[150]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N153 ) );
  AND2_X2 \cv_next_reg/U168  ( .A1(cv_next_d[149]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N152 ) );
  AND2_X2 \cv_next_reg/U167  ( .A1(cv_next_d[148]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N151 ) );
  AND2_X2 \cv_next_reg/U166  ( .A1(cv_next_d[147]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N150 ) );
  AND2_X2 \cv_next_reg/U165  ( .A1(cv_next_d[146]), .A2(\cv_next_reg/n230 ), 
        .ZN(\cv_next_reg/N149 ) );
  AND2_X2 \cv_next_reg/U164  ( .A1(cv_next_d[145]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N148 ) );
  AND2_X2 \cv_next_reg/U163  ( .A1(cv_next_d[144]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N147 ) );
  AND2_X2 \cv_next_reg/U145  ( .A1(cv_next_d[127]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N130 ) );
  AND2_X2 \cv_next_reg/U144  ( .A1(cv_next_d[126]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N129 ) );
  AND2_X2 \cv_next_reg/U143  ( .A1(cv_next_d[125]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N128 ) );
  AND2_X2 \cv_next_reg/U142  ( .A1(cv_next_d[124]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N127 ) );
  AND2_X2 \cv_next_reg/U141  ( .A1(cv_next_d[123]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N126 ) );
  AND2_X2 \cv_next_reg/U139  ( .A1(cv_next_d[122]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N125 ) );
  AND2_X2 \cv_next_reg/U138  ( .A1(cv_next_d[121]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N124 ) );
  AND2_X2 \cv_next_reg/U137  ( .A1(cv_next_d[120]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N123 ) );
  AND2_X2 \cv_next_reg/U136  ( .A1(cv_next_d[119]), .A2(\cv_next_reg/n220 ), 
        .ZN(\cv_next_reg/N122 ) );
  AND2_X2 \cv_next_reg/U135  ( .A1(cv_next_d[118]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N121 ) );
  AND2_X2 \cv_next_reg/U134  ( .A1(cv_next_d[117]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N120 ) );
  AND2_X2 \cv_next_reg/U133  ( .A1(cv_next_d[116]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N119 ) );
  AND2_X2 \cv_next_reg/U132  ( .A1(cv_next_d[115]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N118 ) );
  AND2_X2 \cv_next_reg/U131  ( .A1(cv_next_d[114]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N117 ) );
  AND2_X2 \cv_next_reg/U130  ( .A1(cv_next_d[113]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N116 ) );
  AND2_X2 \cv_next_reg/U128  ( .A1(cv_next_d[112]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N115 ) );
  AND2_X2 \cv_next_reg/U110  ( .A1(cv_next_d[95]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N98 ) );
  AND2_X2 \cv_next_reg/U109  ( .A1(cv_next_d[94]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N97 ) );
  AND2_X2 \cv_next_reg/U108  ( .A1(cv_next_d[93]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N96 ) );
  AND2_X2 \cv_next_reg/U106  ( .A1(cv_next_d[92]), .A2(\cv_next_reg/n210 ), 
        .ZN(\cv_next_reg/N95 ) );
  AND2_X2 \cv_next_reg/U105  ( .A1(cv_next_d[91]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N94 ) );
  AND2_X2 \cv_next_reg/U104  ( .A1(cv_next_d[90]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N93 ) );
  AND2_X2 \cv_next_reg/U103  ( .A1(cv_next_d[89]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N92 ) );
  AND2_X2 \cv_next_reg/U102  ( .A1(cv_next_d[88]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N91 ) );
  AND2_X2 \cv_next_reg/U101  ( .A1(cv_next_d[87]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N90 ) );
  AND2_X2 \cv_next_reg/U100  ( .A1(cv_next_d[86]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N89 ) );
  AND2_X2 \cv_next_reg/U99  ( .A1(cv_next_d[85]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N88 ) );
  AND2_X2 \cv_next_reg/U98  ( .A1(cv_next_d[84]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N87 ) );
  AND2_X2 \cv_next_reg/U97  ( .A1(cv_next_d[83]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N86 ) );
  AND2_X2 \cv_next_reg/U95  ( .A1(cv_next_d[82]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N85 ) );
  AND2_X2 \cv_next_reg/U94  ( .A1(cv_next_d[81]), .A2(\cv_next_reg/n200 ), 
        .ZN(\cv_next_reg/N84 ) );
  AND2_X2 \cv_next_reg/U93  ( .A1(cv_next_d[80]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N83 ) );
  AND2_X2 \cv_next_reg/U90  ( .A1(cv_next_d[63]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N66 ) );
  AND2_X2 \cv_next_reg/U89  ( .A1(cv_next_d[62]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N65 ) );
  AND2_X2 \cv_next_reg/U88  ( .A1(cv_next_d[61]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N64 ) );
  AND2_X2 \cv_next_reg/U87  ( .A1(cv_next_d[60]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N63 ) );
  AND2_X2 \cv_next_reg/U86  ( .A1(cv_next_d[59]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N62 ) );
  AND2_X2 \cv_next_reg/U85  ( .A1(cv_next_d[58]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N61 ) );
  AND2_X2 \cv_next_reg/U84  ( .A1(cv_next_d[57]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N60 ) );
  AND2_X2 \cv_next_reg/U83  ( .A1(cv_next_d[56]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N59 ) );
  AND2_X2 \cv_next_reg/U82  ( .A1(cv_next_d[55]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N58 ) );
  AND2_X2 \cv_next_reg/U81  ( .A1(cv_next_d[54]), .A2(\cv_next_reg/n190 ), 
        .ZN(\cv_next_reg/N57 ) );
  AND2_X2 \cv_next_reg/U80  ( .A1(cv_next_d[53]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N56 ) );
  AND2_X2 \cv_next_reg/U78  ( .A1(cv_next_d[52]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N55 ) );
  AND2_X2 \cv_next_reg/U77  ( .A1(cv_next_d[51]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N54 ) );
  AND2_X2 \cv_next_reg/U76  ( .A1(cv_next_d[50]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N53 ) );
  AND2_X2 \cv_next_reg/U75  ( .A1(cv_next_d[49]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N52 ) );
  AND2_X2 \cv_next_reg/U74  ( .A1(cv_next_d[48]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N51 ) );
  AND2_X2 \cv_next_reg/U55  ( .A1(cv_next_d[31]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N34 ) );
  AND2_X2 \cv_next_reg/U54  ( .A1(cv_next_d[30]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N33 ) );
  AND2_X2 \cv_next_reg/U53  ( .A1(cv_next_d[29]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N32 ) );
  AND2_X2 \cv_next_reg/U52  ( .A1(cv_next_d[28]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N31 ) );
  AND2_X2 \cv_next_reg/U51  ( .A1(cv_next_d[27]), .A2(\cv_next_reg/n180 ), 
        .ZN(\cv_next_reg/N30 ) );
  AND2_X2 \cv_next_reg/U50  ( .A1(cv_next_d[26]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N29 ) );
  AND2_X2 \cv_next_reg/U49  ( .A1(cv_next_d[25]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N28 ) );
  AND2_X2 \cv_next_reg/U48  ( .A1(cv_next_d[24]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N27 ) );
  AND2_X2 \cv_next_reg/U47  ( .A1(cv_next_d[23]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N26 ) );
  AND2_X2 \cv_next_reg/U45  ( .A1(cv_next_d[22]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N25 ) );
  AND2_X2 \cv_next_reg/U44  ( .A1(cv_next_d[21]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N24 ) );
  AND2_X2 \cv_next_reg/U43  ( .A1(cv_next_d[20]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N23 ) );
  AND2_X2 \cv_next_reg/U42  ( .A1(cv_next_d[19]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N22 ) );
  AND2_X2 \cv_next_reg/U41  ( .A1(cv_next_d[18]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N21 ) );
  AND2_X2 \cv_next_reg/U40  ( .A1(cv_next_d[17]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N20 ) );
  AND2_X2 \cv_next_reg/U39  ( .A1(cv_next_d[16]), .A2(\cv_next_reg/n170 ), 
        .ZN(\cv_next_reg/N19 ) );
  INV_X4 \cv_next_reg/U20  ( .A(\cv_next_reg/n250 ), .ZN(\cv_next_reg/n320 )
         );
  INV_X4 \cv_next_reg/U19  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n310 )
         );
  INV_X4 \cv_next_reg/U18  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n220 )
         );
  INV_X4 \cv_next_reg/U17  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n210 )
         );
  INV_X4 \cv_next_reg/U16  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n200 )
         );
  INV_X4 \cv_next_reg/U15  ( .A(n7117), .ZN(\cv_next_reg/n190 ) );
  INV_X4 \cv_next_reg/U14  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n180 )
         );
  INV_X4 \cv_next_reg/U12  ( .A(n7117), .ZN(\cv_next_reg/n170 ) );
  INV_X4 \cv_next_reg/U11  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n240 )
         );
  INV_X4 \cv_next_reg/U10  ( .A(n7117), .ZN(\cv_next_reg/n230 ) );
  INV_X4 \cv_next_reg/U9  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n280 ) );
  INV_X4 \cv_next_reg/U8  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n290 ) );
  INV_X4 \cv_next_reg/U7  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n300 ) );
  INV_X4 \cv_next_reg/U6  ( .A(n7117), .ZN(\cv_next_reg/n250 ) );
  INV_X4 \cv_next_reg/U5  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n260 ) );
  INV_X4 \cv_next_reg/U4  ( .A(\cv_next_reg/n320 ), .ZN(\cv_next_reg/n270 ) );
  AND2_X2 \cv_next_reg/U162  ( .A1(cv_next_d[7]), .A2(\cv_next_reg/n310 ), 
        .ZN(\cv_next_reg/N10 ) );
  AND2_X2 \cv_next_reg/U161  ( .A1(cv_next_d[97]), .A2(\cv_next_reg/n310 ), 
        .ZN(\cv_next_reg/N100 ) );
  AND2_X2 \cv_next_reg/U160  ( .A1(cv_next_d[98]), .A2(\cv_next_reg/n310 ), 
        .ZN(\cv_next_reg/N101 ) );
  AND2_X2 \cv_next_reg/U159  ( .A1(cv_next_d[99]), .A2(\cv_next_reg/n310 ), 
        .ZN(\cv_next_reg/N102 ) );
  AND2_X2 \cv_next_reg/U158  ( .A1(cv_next_d[100]), .A2(\cv_next_reg/n310 ), 
        .ZN(\cv_next_reg/N103 ) );
  AND2_X2 \cv_next_reg/U157  ( .A1(cv_next_d[101]), .A2(\cv_next_reg/n310 ), 
        .ZN(\cv_next_reg/N104 ) );
  AND2_X2 \cv_next_reg/U156  ( .A1(cv_next_d[102]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N105 ) );
  AND2_X2 \cv_next_reg/U155  ( .A1(cv_next_d[103]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N106 ) );
  AND2_X2 \cv_next_reg/U154  ( .A1(cv_next_d[104]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N107 ) );
  AND2_X2 \cv_next_reg/U153  ( .A1(cv_next_d[105]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N108 ) );
  AND2_X2 \cv_next_reg/U152  ( .A1(cv_next_d[106]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N109 ) );
  AND2_X2 \cv_next_reg/U151  ( .A1(cv_next_d[8]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N11 ) );
  AND2_X2 \cv_next_reg/U150  ( .A1(cv_next_d[107]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N110 ) );
  AND2_X2 \cv_next_reg/U149  ( .A1(cv_next_d[108]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N111 ) );
  AND2_X2 \cv_next_reg/U148  ( .A1(cv_next_d[109]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N112 ) );
  AND2_X2 \cv_next_reg/U147  ( .A1(cv_next_d[110]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N113 ) );
  AND2_X2 \cv_next_reg/U146  ( .A1(cv_next_d[111]), .A2(\cv_next_reg/n300 ), 
        .ZN(\cv_next_reg/N114 ) );
  AND2_X2 \cv_next_reg/U140  ( .A1(cv_next_d[9]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N12 ) );
  AND2_X2 \cv_next_reg/U129  ( .A1(cv_next_d[10]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N13 ) );
  AND2_X2 \cv_next_reg/U127  ( .A1(cv_next_d[128]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N131 ) );
  AND2_X2 \cv_next_reg/U126  ( .A1(cv_next_d[129]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N132 ) );
  AND2_X2 \cv_next_reg/U125  ( .A1(cv_next_d[130]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N133 ) );
  AND2_X2 \cv_next_reg/U124  ( .A1(cv_next_d[131]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N134 ) );
  AND2_X2 \cv_next_reg/U123  ( .A1(cv_next_d[132]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N135 ) );
  AND2_X2 \cv_next_reg/U122  ( .A1(cv_next_d[133]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N136 ) );
  AND2_X2 \cv_next_reg/U121  ( .A1(cv_next_d[134]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N137 ) );
  AND2_X2 \cv_next_reg/U120  ( .A1(cv_next_d[135]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N138 ) );
  AND2_X2 \cv_next_reg/U119  ( .A1(cv_next_d[136]), .A2(\cv_next_reg/n290 ), 
        .ZN(\cv_next_reg/N139 ) );
  AND2_X2 \cv_next_reg/U118  ( .A1(cv_next_d[11]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N14 ) );
  AND2_X2 \cv_next_reg/U117  ( .A1(cv_next_d[137]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N140 ) );
  AND2_X2 \cv_next_reg/U116  ( .A1(cv_next_d[138]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N141 ) );
  AND2_X2 \cv_next_reg/U115  ( .A1(cv_next_d[139]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N142 ) );
  AND2_X2 \cv_next_reg/U114  ( .A1(cv_next_d[140]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N143 ) );
  AND2_X2 \cv_next_reg/U113  ( .A1(cv_next_d[141]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N144 ) );
  AND2_X2 \cv_next_reg/U112  ( .A1(cv_next_d[142]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N145 ) );
  AND2_X2 \cv_next_reg/U111  ( .A1(cv_next_d[143]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N146 ) );
  AND2_X2 \cv_next_reg/U107  ( .A1(cv_next_d[12]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N15 ) );
  AND2_X2 \cv_next_reg/U96  ( .A1(cv_next_d[13]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N16 ) );
  AND2_X2 \cv_next_reg/U92  ( .A1(cv_next_d[14]), .A2(\cv_next_reg/n280 ), 
        .ZN(\cv_next_reg/N17 ) );
  AND2_X2 \cv_next_reg/U91  ( .A1(cv_next_d[15]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N18 ) );
  AND2_X2 \cv_next_reg/U79  ( .A1(cv_next_d[0]), .A2(\cv_next_reg/n270 ), .ZN(
        \cv_next_reg/N3 ) );
  AND2_X2 \cv_next_reg/U73  ( .A1(cv_next_d[32]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N35 ) );
  AND2_X2 \cv_next_reg/U72  ( .A1(cv_next_d[33]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N36 ) );
  AND2_X2 \cv_next_reg/U71  ( .A1(cv_next_d[34]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N37 ) );
  AND2_X2 \cv_next_reg/U70  ( .A1(cv_next_d[35]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N38 ) );
  AND2_X2 \cv_next_reg/U69  ( .A1(cv_next_d[36]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N39 ) );
  AND2_X2 \cv_next_reg/U68  ( .A1(cv_next_d[1]), .A2(\cv_next_reg/n270 ), .ZN(
        \cv_next_reg/N4 ) );
  AND2_X2 \cv_next_reg/U67  ( .A1(cv_next_d[37]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N40 ) );
  AND2_X2 \cv_next_reg/U66  ( .A1(cv_next_d[38]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N41 ) );
  AND2_X2 \cv_next_reg/U65  ( .A1(cv_next_d[39]), .A2(\cv_next_reg/n270 ), 
        .ZN(\cv_next_reg/N42 ) );
  AND2_X2 \cv_next_reg/U64  ( .A1(cv_next_d[40]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N43 ) );
  AND2_X2 \cv_next_reg/U63  ( .A1(cv_next_d[41]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N44 ) );
  AND2_X2 \cv_next_reg/U62  ( .A1(cv_next_d[42]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N45 ) );
  AND2_X2 \cv_next_reg/U61  ( .A1(cv_next_d[43]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N46 ) );
  AND2_X2 \cv_next_reg/U60  ( .A1(cv_next_d[44]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N47 ) );
  AND2_X2 \cv_next_reg/U59  ( .A1(cv_next_d[45]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N48 ) );
  AND2_X2 \cv_next_reg/U58  ( .A1(cv_next_d[46]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N49 ) );
  AND2_X2 \cv_next_reg/U57  ( .A1(cv_next_d[2]), .A2(\cv_next_reg/n260 ), .ZN(
        \cv_next_reg/N5 ) );
  AND2_X2 \cv_next_reg/U56  ( .A1(cv_next_d[47]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N50 ) );
  AND2_X2 \cv_next_reg/U46  ( .A1(cv_next_d[3]), .A2(\cv_next_reg/n260 ), .ZN(
        \cv_next_reg/N6 ) );
  AND2_X2 \cv_next_reg/U38  ( .A1(cv_next_d[64]), .A2(\cv_next_reg/n260 ), 
        .ZN(\cv_next_reg/N67 ) );
  AND2_X2 \cv_next_reg/U37  ( .A1(cv_next_d[65]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N68 ) );
  AND2_X2 \cv_next_reg/U36  ( .A1(cv_next_d[66]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N69 ) );
  AND2_X2 \cv_next_reg/U35  ( .A1(cv_next_d[4]), .A2(\cv_next_reg/n250 ), .ZN(
        \cv_next_reg/N7 ) );
  AND2_X2 \cv_next_reg/U34  ( .A1(cv_next_d[67]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N70 ) );
  AND2_X2 \cv_next_reg/U33  ( .A1(cv_next_d[68]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N71 ) );
  AND2_X2 \cv_next_reg/U32  ( .A1(cv_next_d[69]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N72 ) );
  AND2_X2 \cv_next_reg/U31  ( .A1(cv_next_d[70]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N73 ) );
  AND2_X2 \cv_next_reg/U30  ( .A1(cv_next_d[71]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N74 ) );
  AND2_X2 \cv_next_reg/U29  ( .A1(cv_next_d[72]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N75 ) );
  AND2_X2 \cv_next_reg/U28  ( .A1(cv_next_d[73]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N76 ) );
  AND2_X2 \cv_next_reg/U27  ( .A1(cv_next_d[74]), .A2(\cv_next_reg/n250 ), 
        .ZN(\cv_next_reg/N77 ) );
  AND2_X2 \cv_next_reg/U26  ( .A1(cv_next_d[75]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N78 ) );
  AND2_X2 \cv_next_reg/U25  ( .A1(cv_next_d[76]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N79 ) );
  AND2_X2 \cv_next_reg/U24  ( .A1(cv_next_d[5]), .A2(\cv_next_reg/n240 ), .ZN(
        \cv_next_reg/N8 ) );
  AND2_X2 \cv_next_reg/U23  ( .A1(cv_next_d[77]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N80 ) );
  AND2_X2 \cv_next_reg/U22  ( .A1(cv_next_d[78]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N81 ) );
  AND2_X2 \cv_next_reg/U21  ( .A1(cv_next_d[79]), .A2(\cv_next_reg/n240 ), 
        .ZN(\cv_next_reg/N82 ) );
  AND2_X2 \cv_next_reg/U13  ( .A1(cv_next_d[6]), .A2(\cv_next_reg/n240 ), .ZN(
        \cv_next_reg/N9 ) );
  AND2_X2 \cv_next_reg/U3  ( .A1(cv_next_d[96]), .A2(\cv_next_reg/n240 ), .ZN(
        \cv_next_reg/N99 ) );
  DFF_X2 \cv_next_reg/q_reg_0_  ( .D(\cv_next_reg/N3 ), .CK(clk), .Q(
        cv_next[0]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_1_  ( .D(\cv_next_reg/N4 ), .CK(clk), .Q(
        cv_next[1]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_2_  ( .D(\cv_next_reg/N5 ), .CK(clk), .Q(
        cv_next[2]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_3_  ( .D(\cv_next_reg/N6 ), .CK(clk), .Q(
        cv_next[3]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_4_  ( .D(\cv_next_reg/N7 ), .CK(clk), .Q(
        cv_next[4]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_5_  ( .D(\cv_next_reg/N8 ), .CK(clk), .Q(
        cv_next[5]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_6_  ( .D(\cv_next_reg/N9 ), .CK(clk), .Q(
        cv_next[6]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_7_  ( .D(\cv_next_reg/N10 ), .CK(clk), .Q(
        cv_next[7]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_8_  ( .D(\cv_next_reg/N11 ), .CK(clk), .Q(
        cv_next[8]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_9_  ( .D(\cv_next_reg/N12 ), .CK(clk), .Q(
        cv_next[9]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_10_  ( .D(\cv_next_reg/N13 ), .CK(clk), .Q(
        cv_next[10]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_11_  ( .D(\cv_next_reg/N14 ), .CK(clk), .Q(
        cv_next[11]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_12_  ( .D(\cv_next_reg/N15 ), .CK(clk), .Q(
        cv_next[12]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_13_  ( .D(\cv_next_reg/N16 ), .CK(clk), .Q(
        cv_next[13]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_14_  ( .D(\cv_next_reg/N17 ), .CK(clk), .Q(
        cv_next[14]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_15_  ( .D(\cv_next_reg/N18 ), .CK(clk), .Q(
        cv_next[15]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_16_  ( .D(\cv_next_reg/N19 ), .CK(clk), .Q(
        cv_next[16]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_17_  ( .D(\cv_next_reg/N20 ), .CK(clk), .Q(
        cv_next[17]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_18_  ( .D(\cv_next_reg/N21 ), .CK(clk), .Q(
        cv_next[18]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_19_  ( .D(\cv_next_reg/N22 ), .CK(clk), .Q(
        cv_next[19]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_20_  ( .D(\cv_next_reg/N23 ), .CK(clk), .Q(
        cv_next[20]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_21_  ( .D(\cv_next_reg/N24 ), .CK(clk), .Q(
        cv_next[21]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_22_  ( .D(\cv_next_reg/N25 ), .CK(clk), .Q(
        cv_next[22]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_23_  ( .D(\cv_next_reg/N26 ), .CK(clk), .Q(
        cv_next[23]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_24_  ( .D(\cv_next_reg/N27 ), .CK(clk), .Q(
        cv_next[24]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_25_  ( .D(\cv_next_reg/N28 ), .CK(clk), .Q(
        cv_next[25]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_26_  ( .D(\cv_next_reg/N29 ), .CK(clk), .Q(
        cv_next[26]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_27_  ( .D(\cv_next_reg/N30 ), .CK(clk), .Q(
        cv_next[27]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_28_  ( .D(\cv_next_reg/N31 ), .CK(clk), .Q(
        cv_next[28]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_29_  ( .D(\cv_next_reg/N32 ), .CK(clk), .Q(
        cv_next[29]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_30_  ( .D(\cv_next_reg/N33 ), .CK(clk), .Q(
        cv_next[30]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_31_  ( .D(\cv_next_reg/N34 ), .CK(clk), .Q(
        cv_next[31]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_32_  ( .D(\cv_next_reg/N35 ), .CK(clk), .Q(
        cv_next[32]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_33_  ( .D(\cv_next_reg/N36 ), .CK(clk), .Q(
        cv_next[33]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_34_  ( .D(\cv_next_reg/N37 ), .CK(clk), .Q(
        cv_next[34]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_35_  ( .D(\cv_next_reg/N38 ), .CK(clk), .Q(
        cv_next[35]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_36_  ( .D(\cv_next_reg/N39 ), .CK(clk), .Q(
        cv_next[36]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_37_  ( .D(\cv_next_reg/N40 ), .CK(clk), .Q(
        cv_next[37]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_38_  ( .D(\cv_next_reg/N41 ), .CK(clk), .Q(
        cv_next[38]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_39_  ( .D(\cv_next_reg/N42 ), .CK(clk), .Q(
        cv_next[39]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_40_  ( .D(\cv_next_reg/N43 ), .CK(clk), .Q(
        cv_next[40]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_41_  ( .D(\cv_next_reg/N44 ), .CK(clk), .Q(
        cv_next[41]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_42_  ( .D(\cv_next_reg/N45 ), .CK(clk), .Q(
        cv_next[42]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_43_  ( .D(\cv_next_reg/N46 ), .CK(clk), .Q(
        cv_next[43]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_44_  ( .D(\cv_next_reg/N47 ), .CK(clk), .Q(
        cv_next[44]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_45_  ( .D(\cv_next_reg/N48 ), .CK(clk), .Q(
        cv_next[45]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_46_  ( .D(\cv_next_reg/N49 ), .CK(clk), .Q(
        cv_next[46]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_47_  ( .D(\cv_next_reg/N50 ), .CK(clk), .Q(
        cv_next[47]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_48_  ( .D(\cv_next_reg/N51 ), .CK(clk), .Q(
        cv_next[48]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_49_  ( .D(\cv_next_reg/N52 ), .CK(clk), .Q(
        cv_next[49]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_50_  ( .D(\cv_next_reg/N53 ), .CK(clk), .Q(
        cv_next[50]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_51_  ( .D(\cv_next_reg/N54 ), .CK(clk), .Q(
        cv_next[51]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_52_  ( .D(\cv_next_reg/N55 ), .CK(clk), .Q(
        cv_next[52]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_53_  ( .D(\cv_next_reg/N56 ), .CK(clk), .Q(
        cv_next[53]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_54_  ( .D(\cv_next_reg/N57 ), .CK(clk), .Q(
        cv_next[54]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_55_  ( .D(\cv_next_reg/N58 ), .CK(clk), .Q(
        cv_next[55]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_56_  ( .D(\cv_next_reg/N59 ), .CK(clk), .Q(
        cv_next[56]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_57_  ( .D(\cv_next_reg/N60 ), .CK(clk), .Q(
        cv_next[57]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_58_  ( .D(\cv_next_reg/N61 ), .CK(clk), .Q(
        cv_next[58]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_59_  ( .D(\cv_next_reg/N62 ), .CK(clk), .Q(
        cv_next[59]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_60_  ( .D(\cv_next_reg/N63 ), .CK(clk), .Q(
        cv_next[60]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_61_  ( .D(\cv_next_reg/N64 ), .CK(clk), .Q(
        cv_next[61]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_62_  ( .D(\cv_next_reg/N65 ), .CK(clk), .Q(
        cv_next[62]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_63_  ( .D(\cv_next_reg/N66 ), .CK(clk), .Q(
        cv_next[63]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_64_  ( .D(\cv_next_reg/N67 ), .CK(clk), .Q(
        cv_next[64]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_65_  ( .D(\cv_next_reg/N68 ), .CK(clk), .Q(
        cv_next[65]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_66_  ( .D(\cv_next_reg/N69 ), .CK(clk), .Q(
        cv_next[66]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_67_  ( .D(\cv_next_reg/N70 ), .CK(clk), .Q(
        cv_next[67]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_68_  ( .D(\cv_next_reg/N71 ), .CK(clk), .Q(
        cv_next[68]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_69_  ( .D(\cv_next_reg/N72 ), .CK(clk), .Q(
        cv_next[69]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_70_  ( .D(\cv_next_reg/N73 ), .CK(clk), .Q(
        cv_next[70]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_71_  ( .D(\cv_next_reg/N74 ), .CK(clk), .Q(
        cv_next[71]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_72_  ( .D(\cv_next_reg/N75 ), .CK(clk), .Q(
        cv_next[72]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_73_  ( .D(\cv_next_reg/N76 ), .CK(clk), .Q(
        cv_next[73]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_74_  ( .D(\cv_next_reg/N77 ), .CK(clk), .Q(
        cv_next[74]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_75_  ( .D(\cv_next_reg/N78 ), .CK(clk), .Q(
        cv_next[75]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_76_  ( .D(\cv_next_reg/N79 ), .CK(clk), .Q(
        cv_next[76]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_77_  ( .D(\cv_next_reg/N80 ), .CK(clk), .Q(
        cv_next[77]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_78_  ( .D(\cv_next_reg/N81 ), .CK(clk), .Q(
        cv_next[78]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_79_  ( .D(\cv_next_reg/N82 ), .CK(clk), .Q(
        cv_next[79]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_80_  ( .D(\cv_next_reg/N83 ), .CK(clk), .Q(
        cv_next[80]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_81_  ( .D(\cv_next_reg/N84 ), .CK(clk), .Q(
        cv_next[81]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_82_  ( .D(\cv_next_reg/N85 ), .CK(clk), .Q(
        cv_next[82]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_83_  ( .D(\cv_next_reg/N86 ), .CK(clk), .Q(
        cv_next[83]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_84_  ( .D(\cv_next_reg/N87 ), .CK(clk), .Q(
        cv_next[84]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_85_  ( .D(\cv_next_reg/N88 ), .CK(clk), .Q(
        cv_next[85]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_86_  ( .D(\cv_next_reg/N89 ), .CK(clk), .Q(
        cv_next[86]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_87_  ( .D(\cv_next_reg/N90 ), .CK(clk), .Q(
        cv_next[87]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_88_  ( .D(\cv_next_reg/N91 ), .CK(clk), .Q(
        cv_next[88]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_89_  ( .D(\cv_next_reg/N92 ), .CK(clk), .Q(
        cv_next[89]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_90_  ( .D(\cv_next_reg/N93 ), .CK(clk), .Q(
        cv_next[90]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_91_  ( .D(\cv_next_reg/N94 ), .CK(clk), .Q(
        cv_next[91]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_92_  ( .D(\cv_next_reg/N95 ), .CK(clk), .Q(
        cv_next[92]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_93_  ( .D(\cv_next_reg/N96 ), .CK(clk), .Q(
        cv_next[93]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_94_  ( .D(\cv_next_reg/N97 ), .CK(clk), .Q(
        cv_next[94]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_95_  ( .D(\cv_next_reg/N98 ), .CK(clk), .Q(
        cv_next[95]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_96_  ( .D(\cv_next_reg/N99 ), .CK(clk), .Q(
        cv_next[96]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_97_  ( .D(\cv_next_reg/N100 ), .CK(clk), .Q(
        cv_next[97]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_98_  ( .D(\cv_next_reg/N101 ), .CK(clk), .Q(
        cv_next[98]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_99_  ( .D(\cv_next_reg/N102 ), .CK(clk), .Q(
        cv_next[99]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_100_  ( .D(\cv_next_reg/N103 ), .CK(clk), .Q(
        cv_next[100]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_101_  ( .D(\cv_next_reg/N104 ), .CK(clk), .Q(
        cv_next[101]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_102_  ( .D(\cv_next_reg/N105 ), .CK(clk), .Q(
        cv_next[102]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_103_  ( .D(\cv_next_reg/N106 ), .CK(clk), .Q(
        cv_next[103]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_104_  ( .D(\cv_next_reg/N107 ), .CK(clk), .Q(
        cv_next[104]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_105_  ( .D(\cv_next_reg/N108 ), .CK(clk), .Q(
        cv_next[105]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_106_  ( .D(\cv_next_reg/N109 ), .CK(clk), .Q(
        cv_next[106]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_107_  ( .D(\cv_next_reg/N110 ), .CK(clk), .Q(
        cv_next[107]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_108_  ( .D(\cv_next_reg/N111 ), .CK(clk), .Q(
        cv_next[108]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_109_  ( .D(\cv_next_reg/N112 ), .CK(clk), .Q(
        cv_next[109]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_110_  ( .D(\cv_next_reg/N113 ), .CK(clk), .Q(
        cv_next[110]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_111_  ( .D(\cv_next_reg/N114 ), .CK(clk), .Q(
        cv_next[111]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_112_  ( .D(\cv_next_reg/N115 ), .CK(clk), .Q(
        cv_next[112]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_113_  ( .D(\cv_next_reg/N116 ), .CK(clk), .Q(
        cv_next[113]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_114_  ( .D(\cv_next_reg/N117 ), .CK(clk), .Q(
        cv_next[114]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_115_  ( .D(\cv_next_reg/N118 ), .CK(clk), .Q(
        cv_next[115]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_116_  ( .D(\cv_next_reg/N119 ), .CK(clk), .Q(
        cv_next[116]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_117_  ( .D(\cv_next_reg/N120 ), .CK(clk), .Q(
        cv_next[117]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_118_  ( .D(\cv_next_reg/N121 ), .CK(clk), .Q(
        cv_next[118]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_119_  ( .D(\cv_next_reg/N122 ), .CK(clk), .Q(
        cv_next[119]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_120_  ( .D(\cv_next_reg/N123 ), .CK(clk), .Q(
        cv_next[120]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_121_  ( .D(\cv_next_reg/N124 ), .CK(clk), .Q(
        cv_next[121]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_122_  ( .D(\cv_next_reg/N125 ), .CK(clk), .Q(
        cv_next[122]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_123_  ( .D(\cv_next_reg/N126 ), .CK(clk), .Q(
        cv_next[123]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_124_  ( .D(\cv_next_reg/N127 ), .CK(clk), .Q(
        cv_next[124]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_125_  ( .D(\cv_next_reg/N128 ), .CK(clk), .Q(
        cv_next[125]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_126_  ( .D(\cv_next_reg/N129 ), .CK(clk), .Q(
        cv_next[126]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_127_  ( .D(\cv_next_reg/N130 ), .CK(clk), .Q(
        cv_next[127]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_128_  ( .D(\cv_next_reg/N131 ), .CK(clk), .Q(
        cv_next[128]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_129_  ( .D(\cv_next_reg/N132 ), .CK(clk), .Q(
        cv_next[129]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_130_  ( .D(\cv_next_reg/N133 ), .CK(clk), .Q(
        cv_next[130]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_131_  ( .D(\cv_next_reg/N134 ), .CK(clk), .Q(
        cv_next[131]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_132_  ( .D(\cv_next_reg/N135 ), .CK(clk), .Q(
        cv_next[132]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_133_  ( .D(\cv_next_reg/N136 ), .CK(clk), .Q(
        cv_next[133]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_134_  ( .D(\cv_next_reg/N137 ), .CK(clk), .Q(
        cv_next[134]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_135_  ( .D(\cv_next_reg/N138 ), .CK(clk), .Q(
        cv_next[135]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_136_  ( .D(\cv_next_reg/N139 ), .CK(clk), .Q(
        cv_next[136]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_137_  ( .D(\cv_next_reg/N140 ), .CK(clk), .Q(
        cv_next[137]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_138_  ( .D(\cv_next_reg/N141 ), .CK(clk), .Q(
        cv_next[138]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_139_  ( .D(\cv_next_reg/N142 ), .CK(clk), .Q(
        cv_next[139]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_140_  ( .D(\cv_next_reg/N143 ), .CK(clk), .Q(
        cv_next[140]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_141_  ( .D(\cv_next_reg/N144 ), .CK(clk), .Q(
        cv_next[141]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_142_  ( .D(\cv_next_reg/N145 ), .CK(clk), .Q(
        cv_next[142]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_143_  ( .D(\cv_next_reg/N146 ), .CK(clk), .Q(
        cv_next[143]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_144_  ( .D(\cv_next_reg/N147 ), .CK(clk), .Q(
        cv_next[144]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_145_  ( .D(\cv_next_reg/N148 ), .CK(clk), .Q(
        cv_next[145]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_146_  ( .D(\cv_next_reg/N149 ), .CK(clk), .Q(
        cv_next[146]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_147_  ( .D(\cv_next_reg/N150 ), .CK(clk), .Q(
        cv_next[147]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_148_  ( .D(\cv_next_reg/N151 ), .CK(clk), .Q(
        cv_next[148]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_149_  ( .D(\cv_next_reg/N152 ), .CK(clk), .Q(
        cv_next[149]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_150_  ( .D(\cv_next_reg/N153 ), .CK(clk), .Q(
        cv_next[150]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_151_  ( .D(\cv_next_reg/N154 ), .CK(clk), .Q(
        cv_next[151]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_152_  ( .D(\cv_next_reg/N155 ), .CK(clk), .Q(
        cv_next[152]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_153_  ( .D(\cv_next_reg/N156 ), .CK(clk), .Q(
        cv_next[153]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_154_  ( .D(\cv_next_reg/N157 ), .CK(clk), .Q(
        cv_next[154]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_155_  ( .D(\cv_next_reg/N158 ), .CK(clk), .Q(
        cv_next[155]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_156_  ( .D(\cv_next_reg/N159 ), .CK(clk), .Q(
        cv_next[156]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_157_  ( .D(\cv_next_reg/N160 ), .CK(clk), .Q(
        cv_next[157]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_158_  ( .D(\cv_next_reg/N161 ), .CK(clk), .Q(
        cv_next[158]), .QN() );
  DFF_X2 \cv_next_reg/q_reg_159_  ( .D(\cv_next_reg/N162 ), .CK(clk), .Q(
        cv_next[159]), .QN() );
  NAND2_X2 \add_98_2/U411  ( .A1(rnd_q[96]), .A2(cv_q[96]), .ZN(
        \add_98_2/n222 ) );
  INV_X4 \add_98_2/U410  ( .A(\add_98_2/n343 ), .ZN(\add_98_2/n379 ) );
  NAND2_X2 \add_98_2/U409  ( .A1(rnd_q[106]), .A2(cv_q[106]), .ZN(
        \add_98_2/n342 ) );
  NAND2_X2 \add_98_2/U408  ( .A1(\add_98_2/n379 ), .A2(\add_98_2/n342 ), .ZN(
        \add_98_2/n359 ) );
  NAND2_X2 \add_98_2/U407  ( .A1(rnd_q[104]), .A2(cv_q[104]), .ZN(
        \add_98_2/n52 ) );
  NAND2_X2 \add_98_2/U406  ( .A1(rnd_q[97]), .A2(cv_q[97]), .ZN(
        \add_98_2/n375 ) );
  NAND2_X2 \add_98_2/U405  ( .A1(\add_98_2/n375 ), .A2(\add_98_2/n222 ), .ZN(
        \add_98_2/n374 ) );
  NAND2_X2 \add_98_2/U404  ( .A1(\add_98_2/n1 ), .A2(\add_98_2/n374 ), .ZN(
        \add_98_2/n370 ) );
  NAND2_X2 \add_98_2/U403  ( .A1(cv_q[98]), .A2(rnd_q[98]), .ZN(
        \add_98_2/n373 ) );
  INV_X4 \add_98_2/U402  ( .A(\add_98_2/n219 ), .ZN(\add_98_2/n371 ) );
  NAND2_X2 \add_98_2/U401  ( .A1(rnd_q[99]), .A2(cv_q[99]), .ZN(
        \add_98_2/n217 ) );
  INV_X4 \add_98_2/U400  ( .A(\add_98_2/n29 ), .ZN(\add_98_2/n369 ) );
  NAND2_X2 \add_98_2/U399  ( .A1(rnd_q[103]), .A2(cv_q[103]), .ZN(
        \add_98_2/n56 ) );
  NAND2_X2 \add_98_2/U398  ( .A1(rnd_q[102]), .A2(cv_q[102]), .ZN(
        \add_98_2/n368 ) );
  NAND2_X2 \add_98_2/U397  ( .A1(rnd_q[100]), .A2(cv_q[100]), .ZN(
        \add_98_2/n66 ) );
  NAND2_X2 \add_98_2/U396  ( .A1(rnd_q[101]), .A2(cv_q[101]), .ZN(
        \add_98_2/n63 ) );
  NAND2_X2 \add_98_2/U395  ( .A1(\add_98_2/n66 ), .A2(\add_98_2/n63 ), .ZN(
        \add_98_2/n367 ) );
  NAND2_X2 \add_98_2/U394  ( .A1(\add_98_2/n366 ), .A2(\add_98_2/n367 ), .ZN(
        \add_98_2/n365 ) );
  NAND2_X2 \add_98_2/U393  ( .A1(\add_98_2/n35 ), .A2(\add_98_2/n365 ), .ZN(
        \add_98_2/n364 ) );
  NAND2_X2 \add_98_2/U392  ( .A1(\add_98_2/n9 ), .A2(\add_98_2/n363 ), .ZN(
        \add_98_2/n362 ) );
  XNOR2_X2 \add_98_2/U391  ( .A(\add_98_2/n359 ), .B(\add_98_2/n358 ), .ZN(N71) );
  NAND2_X2 \add_98_2/U390  ( .A1(\add_98_2/n358 ), .A2(\add_98_2/n379 ), .ZN(
        \add_98_2/n357 ) );
  NAND2_X2 \add_98_2/U389  ( .A1(\add_98_2/n357 ), .A2(\add_98_2/n342 ), .ZN(
        \add_98_2/n355 ) );
  NAND2_X2 \add_98_2/U388  ( .A1(rnd_q[107]), .A2(cv_q[107]), .ZN(
        \add_98_2/n341 ) );
  NAND2_X2 \add_98_2/U387  ( .A1(\add_98_2/n341 ), .A2(\add_98_2/n308 ), .ZN(
        \add_98_2/n356 ) );
  XNOR2_X2 \add_98_2/U386  ( .A(\add_98_2/n355 ), .B(\add_98_2/n356 ), .ZN(N72) );
  INV_X4 \add_98_2/U385  ( .A(\add_98_2/n43 ), .ZN(\add_98_2/n350 ) );
  INV_X4 \add_98_2/U384  ( .A(\add_98_2/n46 ), .ZN(\add_98_2/n351 ) );
  INV_X4 \add_98_2/U383  ( .A(\add_98_2/n308 ), .ZN(\add_98_2/n353 ) );
  NAND2_X2 \add_98_2/U382  ( .A1(\add_98_2/n345 ), .A2(\add_98_2/n346 ), .ZN(
        \add_98_2/n337 ) );
  NAND2_X2 \add_98_2/U381  ( .A1(cv_q[105]), .A2(rnd_q[105]), .ZN(
        \add_98_2/n344 ) );
  INV_X4 \add_98_2/U380  ( .A(\add_98_2/n342 ), .ZN(\add_98_2/n339 ) );
  INV_X4 \add_98_2/U379  ( .A(\add_98_2/n341 ), .ZN(\add_98_2/n340 ) );
  NAND2_X2 \add_98_2/U378  ( .A1(\add_98_2/n309 ), .A2(\add_98_2/n308 ), .ZN(
        \add_98_2/n332 ) );
  INV_X4 \add_98_2/U377  ( .A(\add_98_2/n332 ), .ZN(\add_98_2/n321 ) );
  NAND2_X2 \add_98_2/U376  ( .A1(rnd_q[108]), .A2(cv_q[108]), .ZN(
        \add_98_2/n322 ) );
  INV_X4 \add_98_2/U375  ( .A(\add_98_2/n322 ), .ZN(\add_98_2/n335 ) );
  XNOR2_X2 \add_98_2/U374  ( .A(\add_98_2/n333 ), .B(\add_98_2/n334 ), .ZN(N73) );
  NAND2_X2 \add_98_2/U373  ( .A1(\add_98_2/n328 ), .A2(\add_98_2/n4 ), .ZN(
        \add_98_2/n331 ) );
  NAND2_X2 \add_98_2/U372  ( .A1(\add_98_2/n331 ), .A2(\add_98_2/n322 ), .ZN(
        \add_98_2/n329 ) );
  NAND2_X2 \add_98_2/U371  ( .A1(rnd_q[109]), .A2(cv_q[109]), .ZN(
        \add_98_2/n323 ) );
  NAND2_X2 \add_98_2/U370  ( .A1(\add_98_2/n323 ), .A2(\add_98_2/n6 ), .ZN(
        \add_98_2/n330 ) );
  XNOR2_X2 \add_98_2/U369  ( .A(\add_98_2/n329 ), .B(\add_98_2/n330 ), .ZN(N74) );
  NAND2_X2 \add_98_2/U368  ( .A1(rnd_q[110]), .A2(cv_q[110]), .ZN(
        \add_98_2/n324 ) );
  NAND2_X2 \add_98_2/U367  ( .A1(\add_98_2/n11 ), .A2(\add_98_2/n324 ), .ZN(
        \add_98_2/n326 ) );
  XNOR2_X2 \add_98_2/U366  ( .A(\add_98_2/n325 ), .B(\add_98_2/n326 ), .ZN(N75) );
  INV_X4 \add_98_2/U365  ( .A(\add_98_2/n300 ), .ZN(\add_98_2/n311 ) );
  INV_X4 \add_98_2/U364  ( .A(\add_98_2/n324 ), .ZN(\add_98_2/n306 ) );
  NAND2_X2 \add_98_2/U363  ( .A1(\add_98_2/n322 ), .A2(\add_98_2/n323 ), .ZN(
        \add_98_2/n319 ) );
  XNOR2_X2 \add_98_2/U362  ( .A(\add_98_2/n313 ), .B(\add_98_2/n314 ), .ZN(N76) );
  NAND2_X2 \add_98_2/U361  ( .A1(rnd_q[112]), .A2(cv_q[112]), .ZN(
        \add_98_2/n280 ) );
  NAND2_X2 \add_98_2/U360  ( .A1(\add_98_2/n280 ), .A2(\add_98_2/n282 ), .ZN(
        \add_98_2/n283 ) );
  INV_X4 \add_98_2/U359  ( .A(\add_98_2/n133 ), .ZN(\add_98_2/n211 ) );
  NAND2_X2 \add_98_2/U358  ( .A1(cv_q[109]), .A2(rnd_q[109]), .ZN(
        \add_98_2/n307 ) );
  NAND2_X2 \add_98_2/U357  ( .A1(rnd_q[108]), .A2(cv_q[108]), .ZN(
        \add_98_2/n302 ) );
  NAND2_X2 \add_98_2/U356  ( .A1(\add_98_2/n299 ), .A2(\add_98_2/n300 ), .ZN(
        \add_98_2/n132 ) );
  INV_X4 \add_98_2/U355  ( .A(\add_98_2/n132 ), .ZN(\add_98_2/n210 ) );
  INV_X4 \add_98_2/U354  ( .A(\add_98_2/n222 ), .ZN(\add_98_2/n298 ) );
  NAND2_X2 \add_98_2/U353  ( .A1(rnd_q[97]), .A2(cv_q[97]), .ZN(
        \add_98_2/n138 ) );
  INV_X4 \add_98_2/U352  ( .A(\add_98_2/n138 ), .ZN(\add_98_2/n260 ) );
  INV_X4 \add_98_2/U351  ( .A(\add_98_2/n217 ), .ZN(\add_98_2/n77 ) );
  NAND2_X2 \add_98_2/U350  ( .A1(\add_98_2/n296 ), .A2(\add_98_2/n297 ), .ZN(
        \add_98_2/n293 ) );
  NAND2_X2 \add_98_2/U349  ( .A1(rnd_q[101]), .A2(cv_q[101]), .ZN(
        \add_98_2/n289 ) );
  NAND2_X2 \add_98_2/U348  ( .A1(\add_98_2/n66 ), .A2(\add_98_2/n289 ), .ZN(
        \add_98_2/n288 ) );
  NAND2_X2 \add_98_2/U347  ( .A1(\add_98_2/n227 ), .A2(\add_98_2/n288 ), .ZN(
        \add_98_2/n287 ) );
  NAND2_X2 \add_98_2/U346  ( .A1(\add_98_2/n35 ), .A2(\add_98_2/n287 ), .ZN(
        \add_98_2/n285 ) );
  NAND3_X2 \add_98_2/U345  ( .A1(\add_98_2/n285 ), .A2(\add_98_2/n3 ), .A3(
        \add_98_2/n286 ), .ZN(\add_98_2/n258 ) );
  INV_X4 \add_98_2/U344  ( .A(\add_98_2/n258 ), .ZN(\add_98_2/n135 ) );
  XNOR2_X2 \add_98_2/U343  ( .A(\add_98_2/n283 ), .B(\add_98_2/n88 ), .ZN(N77)
         );
  INV_X4 \add_98_2/U342  ( .A(\add_98_2/n274 ), .ZN(\add_98_2/n282 ) );
  NAND2_X2 \add_98_2/U341  ( .A1(\add_98_2/n88 ), .A2(\add_98_2/n282 ), .ZN(
        \add_98_2/n281 ) );
  NAND2_X2 \add_98_2/U340  ( .A1(\add_98_2/n280 ), .A2(\add_98_2/n281 ), .ZN(
        \add_98_2/n278 ) );
  NAND2_X2 \add_98_2/U339  ( .A1(rnd_q[113]), .A2(cv_q[113]), .ZN(
        \add_98_2/n275 ) );
  NAND2_X2 \add_98_2/U338  ( .A1(\add_98_2/n40 ), .A2(\add_98_2/n275 ), .ZN(
        \add_98_2/n279 ) );
  XNOR2_X2 \add_98_2/U337  ( .A(\add_98_2/n278 ), .B(\add_98_2/n279 ), .ZN(N78) );
  NAND2_X2 \add_98_2/U336  ( .A1(\add_98_2/n33 ), .A2(\add_98_2/n275 ), .ZN(
        \add_98_2/n265 ) );
  INV_X4 \add_98_2/U335  ( .A(\add_98_2/n265 ), .ZN(\add_98_2/n271 ) );
  NAND2_X2 \add_98_2/U334  ( .A1(\add_98_2/n268 ), .A2(\add_98_2/n88 ), .ZN(
        \add_98_2/n272 ) );
  NAND2_X2 \add_98_2/U333  ( .A1(\add_98_2/n271 ), .A2(\add_98_2/n272 ), .ZN(
        \add_98_2/n269 ) );
  NAND2_X2 \add_98_2/U332  ( .A1(rnd_q[114]), .A2(cv_q[114]), .ZN(
        \add_98_2/n264 ) );
  NAND2_X2 \add_98_2/U331  ( .A1(\add_98_2/n264 ), .A2(\add_98_2/n266 ), .ZN(
        \add_98_2/n270 ) );
  XNOR2_X2 \add_98_2/U330  ( .A(\add_98_2/n269 ), .B(\add_98_2/n270 ), .ZN(N79) );
  INV_X4 \add_98_2/U329  ( .A(\add_98_2/n88 ), .ZN(\add_98_2/n267 ) );
  NAND2_X2 \add_98_2/U328  ( .A1(\add_98_2/n268 ), .A2(\add_98_2/n266 ), .ZN(
        \add_98_2/n256 ) );
  NAND2_X2 \add_98_2/U327  ( .A1(\add_98_2/n265 ), .A2(\add_98_2/n266 ), .ZN(
        \add_98_2/n263 ) );
  NAND2_X2 \add_98_2/U326  ( .A1(\add_98_2/n263 ), .A2(\add_98_2/n264 ), .ZN(
        \add_98_2/n197 ) );
  NAND2_X2 \add_98_2/U325  ( .A1(rnd_q[115]), .A2(cv_q[115]), .ZN(
        \add_98_2/n127 ) );
  XNOR2_X2 \add_98_2/U324  ( .A(\add_98_2/n261 ), .B(\add_98_2/n23 ), .ZN(N80)
         );
  XNOR2_X2 \add_98_2/U323  ( .A(\add_98_2/n222 ), .B(\add_98_2/n259 ), .ZN(N62) );
  INV_X4 \add_98_2/U322  ( .A(\add_98_2/n256 ), .ZN(\add_98_2/n255 ) );
  NAND2_X2 \add_98_2/U321  ( .A1(\add_98_2/n255 ), .A2(\add_98_2/n196 ), .ZN(
        \add_98_2/n129 ) );
  NAND2_X2 \add_98_2/U320  ( .A1(\add_98_2/n197 ), .A2(\add_98_2/n196 ), .ZN(
        \add_98_2/n126 ) );
  NAND2_X2 \add_98_2/U319  ( .A1(\add_98_2/n126 ), .A2(\add_98_2/n127 ), .ZN(
        \add_98_2/n253 ) );
  XNOR2_X2 \add_98_2/U318  ( .A(\add_98_2/n235 ), .B(\add_98_2/n251 ), .ZN(N81) );
  NAND2_X2 \add_98_2/U317  ( .A1(rnd_q[117]), .A2(cv_q[117]), .ZN(
        \add_98_2/n202 ) );
  INV_X4 \add_98_2/U316  ( .A(\add_98_2/n202 ), .ZN(\add_98_2/n248 ) );
  XNOR2_X2 \add_98_2/U315  ( .A(\add_98_2/n246 ), .B(\add_98_2/n247 ), .ZN(N82) );
  INV_X4 \add_98_2/U314  ( .A(\add_98_2/n236 ), .ZN(\add_98_2/n243 ) );
  INV_X4 \add_98_2/U313  ( .A(\add_98_2/n242 ), .ZN(\add_98_2/n241 ) );
  NAND2_X2 \add_98_2/U312  ( .A1(\add_98_2/n203 ), .A2(\add_98_2/n202 ), .ZN(
        \add_98_2/n240 ) );
  NAND2_X2 \add_98_2/U311  ( .A1(rnd_q[118]), .A2(cv_q[118]), .ZN(
        \add_98_2/n204 ) );
  XNOR2_X2 \add_98_2/U310  ( .A(\add_98_2/n238 ), .B(\add_98_2/n26 ), .ZN(N83)
         );
  NAND2_X2 \add_98_2/U309  ( .A1(\add_98_2/n203 ), .A2(\add_98_2/n202 ), .ZN(
        \add_98_2/n237 ) );
  NAND2_X2 \add_98_2/U308  ( .A1(\add_98_2/n237 ), .A2(\add_98_2/n199 ), .ZN(
        \add_98_2/n234 ) );
  NAND2_X2 \add_98_2/U307  ( .A1(\add_98_2/n236 ), .A2(\add_98_2/n199 ), .ZN(
        \add_98_2/n231 ) );
  NAND2_X2 \add_98_2/U306  ( .A1(rnd_q[119]), .A2(cv_q[119]), .ZN(
        \add_98_2/n152 ) );
  NAND2_X2 \add_98_2/U305  ( .A1(\add_98_2/n200 ), .A2(\add_98_2/n152 ), .ZN(
        \add_98_2/n233 ) );
  XNOR2_X2 \add_98_2/U304  ( .A(\add_98_2/n232 ), .B(\add_98_2/n233 ), .ZN(N84) );
  INV_X4 \add_98_2/U303  ( .A(\add_98_2/n231 ), .ZN(\add_98_2/n230 ) );
  NAND2_X2 \add_98_2/U302  ( .A1(\add_98_2/n230 ), .A2(\add_98_2/n200 ), .ZN(
        \add_98_2/n147 ) );
  NAND2_X2 \add_98_2/U301  ( .A1(rnd_q[101]), .A2(cv_q[101]), .ZN(
        \add_98_2/n229 ) );
  NAND2_X2 \add_98_2/U300  ( .A1(\add_98_2/n66 ), .A2(\add_98_2/n229 ), .ZN(
        \add_98_2/n228 ) );
  NAND2_X2 \add_98_2/U299  ( .A1(\add_98_2/n227 ), .A2(\add_98_2/n228 ), .ZN(
        \add_98_2/n226 ) );
  NAND2_X2 \add_98_2/U298  ( .A1(\add_98_2/n35 ), .A2(\add_98_2/n226 ), .ZN(
        \add_98_2/n223 ) );
  INV_X4 \add_98_2/U297  ( .A(\add_98_2/n215 ), .ZN(\add_98_2/n224 ) );
  INV_X4 \add_98_2/U296  ( .A(\add_98_2/n216 ), .ZN(\add_98_2/n225 ) );
  NAND4_X2 \add_98_2/U295  ( .A1(\add_98_2/n223 ), .A2(\add_98_2/n3 ), .A3(
        \add_98_2/n224 ), .A4(\add_98_2/n225 ), .ZN(\add_98_2/n207 ) );
  NAND2_X2 \add_98_2/U294  ( .A1(rnd_q[97]), .A2(cv_q[97]), .ZN(
        \add_98_2/n221 ) );
  NAND2_X2 \add_98_2/U293  ( .A1(\add_98_2/n221 ), .A2(\add_98_2/n222 ), .ZN(
        \add_98_2/n220 ) );
  NAND2_X2 \add_98_2/U292  ( .A1(\add_98_2/n1 ), .A2(\add_98_2/n220 ), .ZN(
        \add_98_2/n218 ) );
  INV_X4 \add_98_2/U291  ( .A(\add_98_2/n49 ), .ZN(\add_98_2/n214 ) );
  NAND2_X2 \add_98_2/U290  ( .A1(\add_98_2/n205 ), .A2(\add_98_2/n206 ), .ZN(
        \add_98_2/n189 ) );
  INV_X4 \add_98_2/U289  ( .A(\add_98_2/n146 ), .ZN(\add_98_2/n198 ) );
  NAND2_X2 \add_98_2/U288  ( .A1(\add_98_2/n198 ), .A2(\add_98_2/n152 ), .ZN(
        \add_98_2/n191 ) );
  INV_X4 \add_98_2/U287  ( .A(\add_98_2/n197 ), .ZN(\add_98_2/n194 ) );
  INV_X4 \add_98_2/U286  ( .A(\add_98_2/n196 ), .ZN(\add_98_2/n195 ) );
  NAND2_X2 \add_98_2/U285  ( .A1(\add_98_2/n189 ), .A2(\add_98_2/n190 ), .ZN(
        \add_98_2/n163 ) );
  NAND2_X2 \add_98_2/U284  ( .A1(rnd_q[120]), .A2(cv_q[120]), .ZN(
        \add_98_2/n187 ) );
  NAND2_X2 \add_98_2/U283  ( .A1(\add_98_2/n187 ), .A2(\add_98_2/n172 ), .ZN(
        \add_98_2/n188 ) );
  XNOR2_X2 \add_98_2/U282  ( .A(\add_98_2/n163 ), .B(\add_98_2/n188 ), .ZN(N85) );
  INV_X4 \add_98_2/U281  ( .A(\add_98_2/n181 ), .ZN(\add_98_2/n172 ) );
  NAND2_X2 \add_98_2/U280  ( .A1(\add_98_2/n172 ), .A2(\add_98_2/n163 ), .ZN(
        \add_98_2/n186 ) );
  NAND2_X2 \add_98_2/U279  ( .A1(\add_98_2/n186 ), .A2(\add_98_2/n187 ), .ZN(
        \add_98_2/n182 ) );
  NAND2_X2 \add_98_2/U278  ( .A1(rnd_q[121]), .A2(cv_q[121]), .ZN(
        \add_98_2/n161 ) );
  INV_X4 \add_98_2/U277  ( .A(rnd_q[121]), .ZN(\add_98_2/n184 ) );
  INV_X4 \add_98_2/U276  ( .A(cv_q[121]), .ZN(\add_98_2/n185 ) );
  NAND2_X2 \add_98_2/U275  ( .A1(\add_98_2/n184 ), .A2(\add_98_2/n185 ), .ZN(
        \add_98_2/n171 ) );
  NAND2_X2 \add_98_2/U274  ( .A1(\add_98_2/n161 ), .A2(\add_98_2/n171 ), .ZN(
        \add_98_2/n183 ) );
  XNOR2_X2 \add_98_2/U273  ( .A(\add_98_2/n182 ), .B(\add_98_2/n183 ), .ZN(N86) );
  INV_X4 \add_98_2/U272  ( .A(\add_98_2/n163 ), .ZN(\add_98_2/n180 ) );
  INV_X4 \add_98_2/U271  ( .A(\add_98_2/n171 ), .ZN(\add_98_2/n178 ) );
  NAND2_X2 \add_98_2/U270  ( .A1(cv_q[120]), .A2(rnd_q[120]), .ZN(
        \add_98_2/n179 ) );
  NAND2_X2 \add_98_2/U269  ( .A1(\add_98_2/n10 ), .A2(\add_98_2/n161 ), .ZN(
        \add_98_2/n177 ) );
  INV_X4 \add_98_2/U268  ( .A(rnd_q[122]), .ZN(\add_98_2/n174 ) );
  INV_X4 \add_98_2/U267  ( .A(cv_q[122]), .ZN(\add_98_2/n175 ) );
  NAND2_X2 \add_98_2/U266  ( .A1(\add_98_2/n174 ), .A2(\add_98_2/n175 ), .ZN(
        \add_98_2/n159 ) );
  NAND2_X2 \add_98_2/U265  ( .A1(rnd_q[122]), .A2(cv_q[122]), .ZN(
        \add_98_2/n162 ) );
  XNOR2_X2 \add_98_2/U264  ( .A(\add_98_2/n173 ), .B(\add_98_2/n24 ), .ZN(N87)
         );
  NAND2_X2 \add_98_2/U263  ( .A1(\add_98_2/n30 ), .A2(\add_98_2/n163 ), .ZN(
        \add_98_2/n168 ) );
  NAND2_X2 \add_98_2/U262  ( .A1(\add_98_2/n170 ), .A2(\add_98_2/n159 ), .ZN(
        \add_98_2/n169 ) );
  NAND2_X2 \add_98_2/U261  ( .A1(\add_98_2/n168 ), .A2(\add_98_2/n169 ), .ZN(
        \add_98_2/n164 ) );
  INV_X4 \add_98_2/U260  ( .A(rnd_q[123]), .ZN(\add_98_2/n166 ) );
  INV_X4 \add_98_2/U259  ( .A(cv_q[123]), .ZN(\add_98_2/n167 ) );
  NAND2_X2 \add_98_2/U258  ( .A1(\add_98_2/n166 ), .A2(\add_98_2/n167 ), .ZN(
        \add_98_2/n150 ) );
  NAND2_X2 \add_98_2/U257  ( .A1(rnd_q[123]), .A2(cv_q[123]), .ZN(
        \add_98_2/n158 ) );
  NAND2_X2 \add_98_2/U256  ( .A1(\add_98_2/n150 ), .A2(\add_98_2/n158 ), .ZN(
        \add_98_2/n165 ) );
  XNOR2_X2 \add_98_2/U255  ( .A(\add_98_2/n164 ), .B(\add_98_2/n165 ), .ZN(N88) );
  NAND2_X2 \add_98_2/U254  ( .A1(\add_98_2/n157 ), .A2(\add_98_2/n158 ), .ZN(
        \add_98_2/n153 ) );
  INV_X4 \add_98_2/U253  ( .A(rnd_q[124]), .ZN(\add_98_2/n155 ) );
  INV_X4 \add_98_2/U252  ( .A(cv_q[124]), .ZN(\add_98_2/n156 ) );
  NAND2_X2 \add_98_2/U251  ( .A1(\add_98_2/n155 ), .A2(\add_98_2/n156 ), .ZN(
        \add_98_2/n151 ) );
  NAND2_X2 \add_98_2/U250  ( .A1(rnd_q[124]), .A2(cv_q[124]), .ZN(
        \add_98_2/n101 ) );
  XNOR2_X2 \add_98_2/U249  ( .A(\add_98_2/n154 ), .B(\add_98_2/n25 ), .ZN(N89)
         );
  INV_X4 \add_98_2/U248  ( .A(\add_98_2/n152 ), .ZN(\add_98_2/n149 ) );
  INV_X4 \add_98_2/U247  ( .A(\add_98_2/n122 ), .ZN(\add_98_2/n104 ) );
  INV_X4 \add_98_2/U246  ( .A(\add_98_2/n101 ), .ZN(\add_98_2/n148 ) );
  INV_X4 \add_98_2/U245  ( .A(\add_98_2/n147 ), .ZN(\add_98_2/n103 ) );
  INV_X4 \add_98_2/U244  ( .A(\add_98_2/n129 ), .ZN(\add_98_2/n87 ) );
  NAND2_X2 \add_98_2/U243  ( .A1(\add_98_2/n126 ), .A2(\add_98_2/n127 ), .ZN(
        \add_98_2/n102 ) );
  NAND2_X2 \add_98_2/U242  ( .A1(\add_98_2/n102 ), .A2(\add_98_2/n14 ), .ZN(
        \add_98_2/n145 ) );
  NAND2_X2 \add_98_2/U241  ( .A1(\add_98_2/n146 ), .A2(\add_98_2/n104 ), .ZN(
        \add_98_2/n93 ) );
  NAND4_X2 \add_98_2/U240  ( .A1(\add_98_2/n143 ), .A2(\add_98_2/n144 ), .A3(
        \add_98_2/n145 ), .A4(\add_98_2/n93 ), .ZN(\add_98_2/n139 ) );
  NAND2_X2 \add_98_2/U239  ( .A1(rnd_q[125]), .A2(cv_q[125]), .ZN(
        \add_98_2/n91 ) );
  INV_X4 \add_98_2/U238  ( .A(rnd_q[125]), .ZN(\add_98_2/n141 ) );
  INV_X4 \add_98_2/U237  ( .A(cv_q[125]), .ZN(\add_98_2/n142 ) );
  NAND2_X2 \add_98_2/U236  ( .A1(\add_98_2/n141 ), .A2(\add_98_2/n142 ), .ZN(
        \add_98_2/n117 ) );
  NAND2_X2 \add_98_2/U235  ( .A1(\add_98_2/n91 ), .A2(\add_98_2/n117 ), .ZN(
        \add_98_2/n140 ) );
  XNOR2_X2 \add_98_2/U234  ( .A(\add_98_2/n139 ), .B(\add_98_2/n140 ), .ZN(N90) );
  XNOR2_X2 \add_98_2/U233  ( .A(\add_98_2/n80 ), .B(\add_98_2/n136 ), .ZN(N63)
         );
  INV_X4 \add_98_2/U232  ( .A(\add_98_2/n134 ), .ZN(\add_98_2/n130 ) );
  NAND2_X2 \add_98_2/U231  ( .A1(\add_98_2/n132 ), .A2(\add_98_2/n133 ), .ZN(
        \add_98_2/n131 ) );
  NAND2_X2 \add_98_2/U230  ( .A1(\add_98_2/n126 ), .A2(\add_98_2/n127 ), .ZN(
        \add_98_2/n125 ) );
  NAND2_X2 \add_98_2/U229  ( .A1(\add_98_2/n103 ), .A2(\add_98_2/n117 ), .ZN(
        \add_98_2/n123 ) );
  NAND2_X2 \add_98_2/U228  ( .A1(\add_98_2/n12 ), .A2(\add_98_2/n117 ), .ZN(
        \add_98_2/n113 ) );
  INV_X4 \add_98_2/U227  ( .A(\add_98_2/n93 ), .ZN(\add_98_2/n120 ) );
  NAND2_X2 \add_98_2/U226  ( .A1(\add_98_2/n120 ), .A2(\add_98_2/n117 ), .ZN(
        \add_98_2/n114 ) );
  INV_X4 \add_98_2/U225  ( .A(\add_98_2/n91 ), .ZN(\add_98_2/n118 ) );
  INV_X4 \add_98_2/U224  ( .A(\add_98_2/n117 ), .ZN(\add_98_2/n105 ) );
  NAND2_X2 \add_98_2/U223  ( .A1(\add_98_2/n19 ), .A2(\add_98_2/n117 ), .ZN(
        \add_98_2/n116 ) );
  NAND4_X2 \add_98_2/U222  ( .A1(\add_98_2/n113 ), .A2(\add_98_2/n114 ), .A3(
        \add_98_2/n115 ), .A4(\add_98_2/n116 ), .ZN(\add_98_2/n112 ) );
  INV_X4 \add_98_2/U221  ( .A(rnd_q[126]), .ZN(\add_98_2/n109 ) );
  INV_X4 \add_98_2/U220  ( .A(cv_q[126]), .ZN(\add_98_2/n110 ) );
  NAND2_X2 \add_98_2/U219  ( .A1(rnd_q[126]), .A2(cv_q[126]), .ZN(
        \add_98_2/n100 ) );
  INV_X4 \add_98_2/U218  ( .A(\add_98_2/n100 ), .ZN(\add_98_2/n108 ) );
  XNOR2_X2 \add_98_2/U217  ( .A(\add_98_2/n106 ), .B(\add_98_2/n107 ), .ZN(N91) );
  NAND2_X2 \add_98_2/U216  ( .A1(\add_98_2/n13 ), .A2(\add_98_2/n102 ), .ZN(
        \add_98_2/n83 ) );
  NAND2_X2 \add_98_2/U215  ( .A1(\add_98_2/n94 ), .A2(\add_98_2/n148 ), .ZN(
        \add_98_2/n99 ) );
  NAND2_X2 \add_98_2/U214  ( .A1(\add_98_2/n99 ), .A2(\add_98_2/n100 ), .ZN(
        \add_98_2/n95 ) );
  NAND2_X2 \add_98_2/U213  ( .A1(\add_98_2/n12 ), .A2(\add_98_2/n94 ), .ZN(
        \add_98_2/n97 ) );
  NAND2_X2 \add_98_2/U212  ( .A1(\add_98_2/n19 ), .A2(\add_98_2/n94 ), .ZN(
        \add_98_2/n98 ) );
  NAND2_X2 \add_98_2/U211  ( .A1(\add_98_2/n97 ), .A2(\add_98_2/n98 ), .ZN(
        \add_98_2/n96 ) );
  INV_X4 \add_98_2/U210  ( .A(\add_98_2/n94 ), .ZN(\add_98_2/n92 ) );
  NAND4_X2 \add_98_2/U209  ( .A1(\add_98_2/n83 ), .A2(\add_98_2/n84 ), .A3(
        \add_98_2/n85 ), .A4(\add_98_2/n86 ), .ZN(\add_98_2/n81 ) );
  XNOR2_X2 \add_98_2/U208  ( .A(rnd_q[127]), .B(cv_q[127]), .ZN(\add_98_2/n82 ) );
  XNOR2_X2 \add_98_2/U207  ( .A(\add_98_2/n81 ), .B(\add_98_2/n82 ), .ZN(N92)
         );
  XNOR2_X2 \add_98_2/U206  ( .A(\add_98_2/n74 ), .B(\add_98_2/n75 ), .ZN(N64)
         );
  INV_X4 \add_98_2/U205  ( .A(\add_98_2/n66 ), .ZN(\add_98_2/n72 ) );
  XNOR2_X2 \add_98_2/U204  ( .A(\add_98_2/n29 ), .B(\add_98_2/n73 ), .ZN(N65)
         );
  INV_X4 \add_98_2/U203  ( .A(\add_98_2/n63 ), .ZN(\add_98_2/n70 ) );
  XNOR2_X2 \add_98_2/U202  ( .A(\add_98_2/n68 ), .B(\add_98_2/n69 ), .ZN(N66)
         );
  NAND2_X2 \add_98_2/U201  ( .A1(rnd_q[102]), .A2(cv_q[102]), .ZN(
        \add_98_2/n58 ) );
  NAND2_X2 \add_98_2/U200  ( .A1(\add_98_2/n58 ), .A2(\add_98_2/n7 ), .ZN(
        \add_98_2/n61 ) );
  NAND2_X2 \add_98_2/U199  ( .A1(\add_98_2/n29 ), .A2(\add_98_2/n66 ), .ZN(
        \add_98_2/n65 ) );
  NAND2_X2 \add_98_2/U198  ( .A1(\add_98_2/n64 ), .A2(\add_98_2/n65 ), .ZN(
        \add_98_2/n62 ) );
  NAND2_X2 \add_98_2/U197  ( .A1(\add_98_2/n62 ), .A2(\add_98_2/n63 ), .ZN(
        \add_98_2/n59 ) );
  XNOR2_X2 \add_98_2/U196  ( .A(\add_98_2/n61 ), .B(\add_98_2/n59 ), .ZN(N67)
         );
  NAND2_X2 \add_98_2/U195  ( .A1(\add_98_2/n59 ), .A2(\add_98_2/n7 ), .ZN(
        \add_98_2/n57 ) );
  NAND2_X2 \add_98_2/U194  ( .A1(\add_98_2/n57 ), .A2(\add_98_2/n58 ), .ZN(
        \add_98_2/n54 ) );
  NAND2_X2 \add_98_2/U193  ( .A1(\add_98_2/n56 ), .A2(\add_98_2/n3 ), .ZN(
        \add_98_2/n55 ) );
  XNOR2_X2 \add_98_2/U192  ( .A(\add_98_2/n54 ), .B(\add_98_2/n55 ), .ZN(N68)
         );
  INV_X4 \add_98_2/U191  ( .A(\add_98_2/n52 ), .ZN(\add_98_2/n45 ) );
  XNOR2_X2 \add_98_2/U190  ( .A(\add_98_2/n50 ), .B(\add_98_2/n51 ), .ZN(N69)
         );
  XNOR2_X2 \add_98_2/U189  ( .A(\add_98_2/n41 ), .B(\add_98_2/n42 ), .ZN(N70)
         );
  NAND2_X2 \add_98_2/U188  ( .A1(\add_98_2/n258 ), .A2(\add_98_2/n134 ), .ZN(
        \add_98_2/n257 ) );
  NOR2_X2 \add_98_2/U187  ( .A1(\add_98_2/n20 ), .A2(\add_98_2/n108 ), .ZN(
        \add_98_2/n107 ) );
  NOR2_X2 \add_98_2/U186  ( .A1(\add_98_2/n242 ), .A2(\add_98_2/n248 ), .ZN(
        \add_98_2/n247 ) );
  NOR2_X2 \add_98_2/U185  ( .A1(\add_98_2/n38 ), .A2(\add_98_2/n43 ), .ZN(
        \add_98_2/n42 ) );
  NOR2_X2 \add_98_2/U184  ( .A1(\add_98_2/n70 ), .A2(\add_98_2/n67 ), .ZN(
        \add_98_2/n69 ) );
  NOR2_X2 \add_98_2/U183  ( .A1(\add_98_2/n36 ), .A2(\add_98_2/n72 ), .ZN(
        \add_98_2/n73 ) );
  NOR2_X2 \add_98_2/U182  ( .A1(\add_98_2/n39 ), .A2(\add_98_2/n79 ), .ZN(
        \add_98_2/n136 ) );
  NOR2_X2 \add_98_2/U181  ( .A1(\add_98_2/n260 ), .A2(\add_98_2/n137 ), .ZN(
        \add_98_2/n259 ) );
  AND2_X2 \add_98_2/U180  ( .A1(cv_q[104]), .A2(rnd_q[104]), .ZN(
        \add_98_2/n345 ) );
  NOR2_X1 \add_98_2/U179  ( .A1(cv_q[105]), .A2(rnd_q[105]), .ZN(
        \add_98_2/n347 ) );
  NOR2_X1 \add_98_2/U178  ( .A1(cv_q[106]), .A2(rnd_q[106]), .ZN(
        \add_98_2/n348 ) );
  NOR2_X2 \add_98_2/U177  ( .A1(\add_98_2/n347 ), .A2(\add_98_2/n348 ), .ZN(
        \add_98_2/n346 ) );
  NOR2_X2 \add_98_2/U176  ( .A1(\add_98_2/n311 ), .A2(\add_98_2/n34 ), .ZN(
        \add_98_2/n313 ) );
  NOR2_X2 \add_98_2/U175  ( .A1(\add_98_2/n335 ), .A2(\add_98_2/n312 ), .ZN(
        \add_98_2/n334 ) );
  NOR2_X2 \add_98_2/U174  ( .A1(\add_98_2/n76 ), .A2(\add_98_2/n77 ), .ZN(
        \add_98_2/n75 ) );
  AND2_X2 \add_98_2/U173  ( .A1(rnd_q[98]), .A2(cv_q[98]), .ZN(\add_98_2/n39 )
         );
  AND2_X2 \add_98_2/U172  ( .A1(rnd_q[105]), .A2(cv_q[105]), .ZN(
        \add_98_2/n38 ) );
  AND2_X2 \add_98_2/U171  ( .A1(rnd_q[116]), .A2(cv_q[116]), .ZN(
        \add_98_2/n37 ) );
  NOR2_X1 \add_98_2/U170  ( .A1(cv_q[113]), .A2(rnd_q[113]), .ZN(
        \add_98_2/n273 ) );
  NOR2_X2 \add_98_2/U169  ( .A1(\add_98_2/n273 ), .A2(\add_98_2/n274 ), .ZN(
        \add_98_2/n268 ) );
  NOR2_X1 \add_98_2/U168  ( .A1(cv_q[101]), .A2(rnd_q[101]), .ZN(
        \add_98_2/n290 ) );
  NOR2_X1 \add_98_2/U167  ( .A1(cv_q[102]), .A2(rnd_q[102]), .ZN(
        \add_98_2/n291 ) );
  NOR2_X2 \add_98_2/U166  ( .A1(\add_98_2/n290 ), .A2(\add_98_2/n291 ), .ZN(
        \add_98_2/n227 ) );
  AND2_X2 \add_98_2/U165  ( .A1(\add_98_2/n56 ), .A2(\add_98_2/n368 ), .ZN(
        \add_98_2/n35 ) );
  AND2_X2 \add_98_2/U164  ( .A1(rnd_q[111]), .A2(cv_q[111]), .ZN(
        \add_98_2/n34 ) );
  NOR2_X1 \add_98_2/U163  ( .A1(cv_q[113]), .A2(rnd_q[113]), .ZN(
        \add_98_2/n276 ) );
  NOR2_X2 \add_98_2/U162  ( .A1(\add_98_2/n46 ), .A2(\add_98_2/n45 ), .ZN(
        \add_98_2/n51 ) );
  NOR2_X2 \add_98_2/U161  ( .A1(\add_98_2/n37 ), .A2(\add_98_2/n250 ), .ZN(
        \add_98_2/n251 ) );
  NOR2_X1 \add_98_2/U160  ( .A1(cv_q[116]), .A2(rnd_q[116]), .ZN(
        \add_98_2/n245 ) );
  NOR2_X1 \add_98_2/U159  ( .A1(cv_q[117]), .A2(rnd_q[117]), .ZN(
        \add_98_2/n244 ) );
  NOR2_X2 \add_98_2/U158  ( .A1(\add_98_2/n244 ), .A2(\add_98_2/n245 ), .ZN(
        \add_98_2/n236 ) );
  NOR2_X1 \add_98_2/U157  ( .A1(cv_q[101]), .A2(rnd_q[101]), .ZN(
        \add_98_2/n377 ) );
  NOR2_X1 \add_98_2/U156  ( .A1(cv_q[117]), .A2(rnd_q[117]), .ZN(
        \add_98_2/n242 ) );
  OR2_X2 \add_98_2/U155  ( .A1(\add_98_2/n276 ), .A2(\add_98_2/n277 ), .ZN(
        \add_98_2/n33 ) );
  NOR2_X1 \add_98_2/U154  ( .A1(cv_q[99]), .A2(rnd_q[99]), .ZN(\add_98_2/n76 )
         );
  NOR2_X1 \add_98_2/U153  ( .A1(cv_q[98]), .A2(rnd_q[98]), .ZN(\add_98_2/n79 )
         );
  NOR2_X1 \add_98_2/U152  ( .A1(cv_q[97]), .A2(rnd_q[97]), .ZN(\add_98_2/n137 ) );
  NAND3_X1 \add_98_2/U151  ( .A1(cv_q[116]), .A2(rnd_q[116]), .A3(
        \add_98_2/n241 ), .ZN(\add_98_2/n203 ) );
  NOR2_X1 \add_98_2/U150  ( .A1(cv_q[116]), .A2(rnd_q[116]), .ZN(
        \add_98_2/n250 ) );
  OR2_X2 \add_98_2/U149  ( .A1(rnd_q[119]), .A2(cv_q[119]), .ZN(
        \add_98_2/n200 ) );
  NOR2_X1 \add_98_2/U148  ( .A1(cv_q[112]), .A2(rnd_q[112]), .ZN(
        \add_98_2/n274 ) );
  NOR2_X1 \add_98_2/U147  ( .A1(cv_q[102]), .A2(rnd_q[102]), .ZN(
        \add_98_2/n60 ) );
  NOR2_X2 \add_98_2/U146  ( .A1(cv_q[120]), .A2(rnd_q[120]), .ZN(
        \add_98_2/n181 ) );
  NOR2_X1 \add_98_2/U145  ( .A1(cv_q[101]), .A2(rnd_q[101]), .ZN(
        \add_98_2/n67 ) );
  NOR2_X2 \add_98_2/U144  ( .A1(\add_98_2/n76 ), .A2(\add_98_2/n373 ), .ZN(
        \add_98_2/n219 ) );
  NOR2_X2 \add_98_2/U143  ( .A1(\add_98_2/n303 ), .A2(\add_98_2/n307 ), .ZN(
        \add_98_2/n305 ) );
  NOR3_X2 \add_98_2/U142  ( .A1(\add_98_2/n302 ), .A2(\add_98_2/n303 ), .A3(
        \add_98_2/n304 ), .ZN(\add_98_2/n301 ) );
  NOR2_X2 \add_98_2/U141  ( .A1(\add_98_2/n298 ), .A2(\add_98_2/n219 ), .ZN(
        \add_98_2/n296 ) );
  NAND3_X2 \add_98_2/U140  ( .A1(\add_98_2/n214 ), .A2(\add_98_2/n363 ), .A3(
        \add_98_2/n369 ), .ZN(\add_98_2/n361 ) );
  NOR2_X2 \add_98_2/U139  ( .A1(\add_98_2/n38 ), .A2(\add_98_2/n378 ), .ZN(
        \add_98_2/n360 ) );
  NAND3_X2 \add_98_2/U138  ( .A1(\add_98_2/n360 ), .A2(\add_98_2/n361 ), .A3(
        \add_98_2/n362 ), .ZN(\add_98_2/n358 ) );
  NAND3_X2 \add_98_2/U137  ( .A1(\add_98_2/n328 ), .A2(\add_98_2/n6 ), .A3(
        \add_98_2/n4 ), .ZN(\add_98_2/n327 ) );
  NAND3_X2 \add_98_2/U136  ( .A1(\add_98_2/n22 ), .A2(\add_98_2/n323 ), .A3(
        \add_98_2/n327 ), .ZN(\add_98_2/n325 ) );
  NOR2_X2 \add_98_2/U135  ( .A1(\add_98_2/n79 ), .A2(\add_98_2/n80 ), .ZN(
        \add_98_2/n78 ) );
  NOR2_X2 \add_98_2/U134  ( .A1(\add_98_2/n78 ), .A2(\add_98_2/n39 ), .ZN(
        \add_98_2/n74 ) );
  NOR2_X2 \add_98_2/U133  ( .A1(\add_98_2/n18 ), .A2(\add_98_2/n153 ), .ZN(
        \add_98_2/n154 ) );
  NOR2_X2 \add_98_2/U132  ( .A1(\add_98_2/n29 ), .A2(\add_98_2/n49 ), .ZN(
        \add_98_2/n48 ) );
  NOR2_X2 \add_98_2/U131  ( .A1(\add_98_2/n48 ), .A2(\add_98_2/n9 ), .ZN(
        \add_98_2/n47 ) );
  NOR2_X2 \add_98_2/U130  ( .A1(\add_98_2/n46 ), .A2(\add_98_2/n47 ), .ZN(
        \add_98_2/n44 ) );
  NOR2_X2 \add_98_2/U129  ( .A1(\add_98_2/n44 ), .A2(\add_98_2/n45 ), .ZN(
        \add_98_2/n41 ) );
  NOR2_X2 \add_98_2/U128  ( .A1(\add_98_2/n29 ), .A2(\add_98_2/n36 ), .ZN(
        \add_98_2/n71 ) );
  NOR2_X2 \add_98_2/U127  ( .A1(\add_98_2/n71 ), .A2(\add_98_2/n72 ), .ZN(
        \add_98_2/n68 ) );
  NOR2_X2 \add_98_2/U126  ( .A1(\add_98_2/n60 ), .A2(\add_98_2/n67 ), .ZN(
        \add_98_2/n366 ) );
  NOR2_X2 \add_98_2/U125  ( .A1(\add_98_2/n235 ), .A2(\add_98_2/n243 ), .ZN(
        \add_98_2/n239 ) );
  NOR2_X2 \add_98_2/U124  ( .A1(\add_98_2/n239 ), .A2(\add_98_2/n240 ), .ZN(
        \add_98_2/n238 ) );
  NOR2_X2 \add_98_2/U123  ( .A1(\add_98_2/n36 ), .A2(\add_98_2/n67 ), .ZN(
        \add_98_2/n64 ) );
  NOR2_X2 \add_98_2/U122  ( .A1(\add_98_2/n20 ), .A2(\add_98_2/n91 ), .ZN(
        \add_98_2/n90 ) );
  NAND3_X2 \add_98_2/U121  ( .A1(\add_98_2/n202 ), .A2(\add_98_2/n203 ), .A3(
        \add_98_2/n204 ), .ZN(\add_98_2/n201 ) );
  AND2_X4 \add_98_2/U120  ( .A1(\add_98_2/n199 ), .A2(\add_98_2/n200 ), .ZN(
        \add_98_2/n32 ) );
  AND2_X2 \add_98_2/U119  ( .A1(\add_98_2/n201 ), .A2(\add_98_2/n32 ), .ZN(
        \add_98_2/n146 ) );
  OR2_X4 \add_98_2/U118  ( .A1(\add_98_2/n137 ), .A2(\add_98_2/n222 ), .ZN(
        \add_98_2/n31 ) );
  AND2_X2 \add_98_2/U117  ( .A1(\add_98_2/n138 ), .A2(\add_98_2/n31 ), .ZN(
        \add_98_2/n80 ) );
  NOR2_X2 \add_98_2/U116  ( .A1(\add_98_2/n105 ), .A2(\add_98_2/n101 ), .ZN(
        \add_98_2/n119 ) );
  NOR2_X2 \add_98_2/U115  ( .A1(\add_98_2/n250 ), .A2(\add_98_2/n235 ), .ZN(
        \add_98_2/n249 ) );
  NOR2_X2 \add_98_2/U114  ( .A1(\add_98_2/n249 ), .A2(\add_98_2/n37 ), .ZN(
        \add_98_2/n246 ) );
  NOR3_X2 \add_98_2/U113  ( .A1(\add_98_2/n135 ), .A2(\add_98_2/n130 ), .A3(
        \add_98_2/n131 ), .ZN(\add_98_2/n128 ) );
  NOR2_X2 \add_98_2/U112  ( .A1(\add_98_2/n128 ), .A2(\add_98_2/n129 ), .ZN(
        \add_98_2/n124 ) );
  NOR2_X2 \add_98_2/U111  ( .A1(\add_98_2/n124 ), .A2(\add_98_2/n125 ), .ZN(
        \add_98_2/n121 ) );
  NOR2_X2 \add_98_2/U110  ( .A1(\add_98_2/n312 ), .A2(\add_98_2/n15 ), .ZN(
        \add_98_2/n318 ) );
  NOR2_X2 \add_98_2/U109  ( .A1(\add_98_2/n43 ), .A2(\add_98_2/n52 ), .ZN(
        \add_98_2/n378 ) );
  NOR2_X2 \add_98_2/U108  ( .A1(\add_98_2/n147 ), .A2(\add_98_2/n127 ), .ZN(
        \add_98_2/n193 ) );
  AND3_X2 \add_98_2/U107  ( .A1(\add_98_2/n171 ), .A2(\add_98_2/n159 ), .A3(
        \add_98_2/n172 ), .ZN(\add_98_2/n30 ) );
  NAND3_X2 \add_98_2/U106  ( .A1(\add_98_2/n150 ), .A2(\add_98_2/n151 ), .A3(
        \add_98_2/n30 ), .ZN(\add_98_2/n122 ) );
  NOR3_X2 \add_98_2/U105  ( .A1(\add_98_2/n194 ), .A2(\add_98_2/n147 ), .A3(
        \add_98_2/n195 ), .ZN(\add_98_2/n192 ) );
  NOR2_X2 \add_98_2/U104  ( .A1(\add_98_2/n312 ), .A2(\add_98_2/n15 ), .ZN(
        \add_98_2/n328 ) );
  NOR2_X2 \add_98_2/U103  ( .A1(\add_98_2/n46 ), .A2(\add_98_2/n43 ), .ZN(
        \add_98_2/n363 ) );
  NAND3_X2 \add_98_2/U102  ( .A1(\add_98_2/n217 ), .A2(\add_98_2/n218 ), .A3(
        \add_98_2/n371 ), .ZN(\add_98_2/n212 ) );
  NAND3_X2 \add_98_2/U101  ( .A1(\add_98_2/n161 ), .A2(\add_98_2/n10 ), .A3(
        \add_98_2/n162 ), .ZN(\add_98_2/n160 ) );
  NAND3_X2 \add_98_2/U100  ( .A1(\add_98_2/n159 ), .A2(\add_98_2/n150 ), .A3(
        \add_98_2/n160 ), .ZN(\add_98_2/n157 ) );
  NOR2_X2 \add_98_2/U99  ( .A1(\add_98_2/n36 ), .A2(\add_98_2/n377 ), .ZN(
        \add_98_2/n376 ) );
  NAND3_X2 \add_98_2/U98  ( .A1(\add_98_2/n3 ), .A2(\add_98_2/n7 ), .A3(
        \add_98_2/n376 ), .ZN(\add_98_2/n49 ) );
  NOR2_X2 \add_98_2/U97  ( .A1(\add_98_2/n20 ), .A2(\add_98_2/n105 ), .ZN(
        \add_98_2/n94 ) );
  AND3_X2 \add_98_2/U96  ( .A1(\add_98_2/n371 ), .A2(\add_98_2/n217 ), .A3(
        \add_98_2/n370 ), .ZN(\add_98_2/n29 ) );
  OR3_X4 \add_98_2/U95  ( .A1(\add_98_2/n305 ), .A2(\add_98_2/n306 ), .A3(
        \add_98_2/n34 ), .ZN(\add_98_2/n28 ) );
  OR2_X2 \add_98_2/U94  ( .A1(\add_98_2/n28 ), .A2(\add_98_2/n301 ), .ZN(
        \add_98_2/n299 ) );
  NOR2_X2 \add_98_2/U93  ( .A1(\add_98_2/n210 ), .A2(\add_98_2/n211 ), .ZN(
        \add_98_2/n209 ) );
  NAND3_X2 \add_98_2/U92  ( .A1(\add_98_2/n212 ), .A2(\add_98_2/n213 ), .A3(
        \add_98_2/n214 ), .ZN(\add_98_2/n208 ) );
  NAND3_X2 \add_98_2/U91  ( .A1(\add_98_2/n208 ), .A2(\add_98_2/n209 ), .A3(
        \add_98_2/n207 ), .ZN(\add_98_2/n206 ) );
  NAND3_X2 \add_98_2/U90  ( .A1(\add_98_2/n234 ), .A2(\add_98_2/n204 ), .A3(
        \add_98_2/n17 ), .ZN(\add_98_2/n232 ) );
  NOR3_X2 \add_98_2/U89  ( .A1(\add_98_2/n180 ), .A2(\add_98_2/n178 ), .A3(
        \add_98_2/n181 ), .ZN(\add_98_2/n176 ) );
  NOR2_X2 \add_98_2/U88  ( .A1(\add_98_2/n176 ), .A2(\add_98_2/n177 ), .ZN(
        \add_98_2/n173 ) );
  NOR2_X2 \add_98_2/U87  ( .A1(\add_98_2/n339 ), .A2(\add_98_2/n340 ), .ZN(
        \add_98_2/n338 ) );
  NAND3_X2 \add_98_2/U86  ( .A1(\add_98_2/n337 ), .A2(\add_98_2/n16 ), .A3(
        \add_98_2/n338 ), .ZN(\add_98_2/n309 ) );
  NAND3_X2 \add_98_2/U85  ( .A1(\add_98_2/n224 ), .A2(\add_98_2/n308 ), .A3(
        \add_98_2/n309 ), .ZN(\add_98_2/n133 ) );
  NAND3_X2 \add_98_2/U84  ( .A1(\add_98_2/n162 ), .A2(\add_98_2/n10 ), .A3(
        \add_98_2/n161 ), .ZN(\add_98_2/n170 ) );
  NOR2_X2 \add_98_2/U83  ( .A1(\add_98_2/n311 ), .A2(\add_98_2/n312 ), .ZN(
        \add_98_2/n310 ) );
  NAND3_X2 \add_98_2/U82  ( .A1(\add_98_2/n6 ), .A2(\add_98_2/n11 ), .A3(
        \add_98_2/n310 ), .ZN(\add_98_2/n215 ) );
  NOR3_X2 \add_98_2/U81  ( .A1(\add_98_2/n257 ), .A2(\add_98_2/n211 ), .A3(
        \add_98_2/n210 ), .ZN(\add_98_2/n254 ) );
  NOR2_X2 \add_98_2/U80  ( .A1(\add_98_2/n254 ), .A2(\add_98_2/n129 ), .ZN(
        \add_98_2/n252 ) );
  NOR2_X2 \add_98_2/U79  ( .A1(\add_98_2/n252 ), .A2(\add_98_2/n253 ), .ZN(
        \add_98_2/n235 ) );
  NOR3_X2 \add_98_2/U78  ( .A1(\add_98_2/n219 ), .A2(\add_98_2/n77 ), .A3(
        \add_98_2/n1 ), .ZN(\add_98_2/n295 ) );
  NOR2_X2 \add_98_2/U77  ( .A1(\add_98_2/n343 ), .A2(\add_98_2/n353 ), .ZN(
        \add_98_2/n352 ) );
  NAND3_X2 \add_98_2/U76  ( .A1(\add_98_2/n350 ), .A2(\add_98_2/n351 ), .A3(
        \add_98_2/n352 ), .ZN(\add_98_2/n216 ) );
  NOR2_X2 \add_98_2/U75  ( .A1(\add_98_2/n215 ), .A2(\add_98_2/n216 ), .ZN(
        \add_98_2/n286 ) );
  NOR3_X2 \add_98_2/U74  ( .A1(\add_98_2/n191 ), .A2(\add_98_2/n192 ), .A3(
        \add_98_2/n193 ), .ZN(\add_98_2/n190 ) );
  NOR2_X2 \add_98_2/U73  ( .A1(\add_98_2/n267 ), .A2(\add_98_2/n256 ), .ZN(
        \add_98_2/n262 ) );
  NOR2_X2 \add_98_2/U72  ( .A1(\add_98_2/n262 ), .A2(\add_98_2/n197 ), .ZN(
        \add_98_2/n261 ) );
  NOR2_X2 \add_98_2/U71  ( .A1(\add_98_2/n118 ), .A2(\add_98_2/n119 ), .ZN(
        \add_98_2/n115 ) );
  NOR3_X2 \add_98_2/U70  ( .A1(\add_98_2/n121 ), .A2(\add_98_2/n122 ), .A3(
        \add_98_2/n123 ), .ZN(\add_98_2/n111 ) );
  NOR2_X2 \add_98_2/U69  ( .A1(\add_98_2/n111 ), .A2(\add_98_2/n112 ), .ZN(
        \add_98_2/n106 ) );
  NOR2_X2 \add_98_2/U68  ( .A1(\add_98_2/n29 ), .A2(\add_98_2/n49 ), .ZN(
        \add_98_2/n53 ) );
  NOR2_X2 \add_98_2/U67  ( .A1(\add_98_2/n53 ), .A2(\add_98_2/n9 ), .ZN(
        \add_98_2/n50 ) );
  NOR2_X2 \add_98_2/U66  ( .A1(\add_98_2/n129 ), .A2(\add_98_2/n147 ), .ZN(
        \add_98_2/n205 ) );
  NOR2_X2 \add_98_2/U65  ( .A1(\add_98_2/n92 ), .A2(\add_98_2/n93 ), .ZN(
        \add_98_2/n89 ) );
  NOR2_X2 \add_98_2/U64  ( .A1(\add_98_2/n29 ), .A2(\add_98_2/n49 ), .ZN(
        \add_98_2/n354 ) );
  NOR2_X2 \add_98_2/U63  ( .A1(\add_98_2/n354 ), .A2(\add_98_2/n9 ), .ZN(
        \add_98_2/n349 ) );
  NOR2_X2 \add_98_2/U62  ( .A1(\add_98_2/n349 ), .A2(\add_98_2/n216 ), .ZN(
        \add_98_2/n336 ) );
  NOR2_X2 \add_98_2/U61  ( .A1(\add_98_2/n336 ), .A2(\add_98_2/n321 ), .ZN(
        \add_98_2/n333 ) );
  NOR2_X2 \add_98_2/U60  ( .A1(\add_98_2/n215 ), .A2(\add_98_2/n216 ), .ZN(
        \add_98_2/n213 ) );
  NOR2_X2 \add_98_2/U59  ( .A1(\add_98_2/n318 ), .A2(\add_98_2/n319 ), .ZN(
        \add_98_2/n317 ) );
  NOR3_X2 \add_98_2/U58  ( .A1(\add_98_2/n316 ), .A2(\add_98_2/n317 ), .A3(
        \add_98_2/n21 ), .ZN(\add_98_2/n315 ) );
  NOR2_X2 \add_98_2/U57  ( .A1(\add_98_2/n306 ), .A2(\add_98_2/n315 ), .ZN(
        \add_98_2/n314 ) );
  NOR2_X2 \add_98_2/U56  ( .A1(\add_98_2/n29 ), .A2(\add_98_2/n49 ), .ZN(
        \add_98_2/n320 ) );
  NAND3_X2 \add_98_2/U55  ( .A1(\add_98_2/n88 ), .A2(\add_98_2/n14 ), .A3(
        \add_98_2/n87 ), .ZN(\add_98_2/n144 ) );
  NOR3_X2 \add_98_2/U54  ( .A1(\add_98_2/n19 ), .A2(\add_98_2/n12 ), .A3(
        \add_98_2/n148 ), .ZN(\add_98_2/n143 ) );
  NOR2_X2 \add_98_2/U53  ( .A1(\add_98_2/n95 ), .A2(\add_98_2/n96 ), .ZN(
        \add_98_2/n84 ) );
  NOR2_X2 \add_98_2/U52  ( .A1(\add_98_2/n89 ), .A2(\add_98_2/n90 ), .ZN(
        \add_98_2/n85 ) );
  NOR4_X2 \add_98_2/U51  ( .A1(\add_98_2/n320 ), .A2(\add_98_2/n321 ), .A3(
        \add_98_2/n9 ), .A4(\add_98_2/n319 ), .ZN(\add_98_2/n316 ) );
  NOR2_X2 \add_98_2/U50  ( .A1(\add_98_2/n260 ), .A2(\add_98_2/n77 ), .ZN(
        \add_98_2/n297 ) );
  NOR2_X2 \add_98_2/U49  ( .A1(\add_98_2/n49 ), .A2(\add_98_2/n295 ), .ZN(
        \add_98_2/n294 ) );
  NOR2_X2 \add_98_2/U48  ( .A1(\add_98_2/n215 ), .A2(\add_98_2/n216 ), .ZN(
        \add_98_2/n292 ) );
  NAND3_X2 \add_98_2/U47  ( .A1(\add_98_2/n292 ), .A2(\add_98_2/n293 ), .A3(
        \add_98_2/n294 ), .ZN(\add_98_2/n134 ) );
  NAND3_X2 \add_98_2/U46  ( .A1(\add_98_2/n87 ), .A2(\add_98_2/n88 ), .A3(
        \add_98_2/n13 ), .ZN(\add_98_2/n86 ) );
  NOR2_X2 \add_98_2/U45  ( .A1(\add_98_2/n211 ), .A2(\add_98_2/n210 ), .ZN(
        \add_98_2/n284 ) );
  NAND3_X2 \add_98_2/U44  ( .A1(\add_98_2/n284 ), .A2(\add_98_2/n134 ), .A3(
        \add_98_2/n258 ), .ZN(\add_98_2/n88 ) );
  OR2_X4 \add_98_2/U43  ( .A1(rnd_q[96]), .A2(cv_q[96]), .ZN(\add_98_2/n372 )
         );
  OR2_X1 \add_98_2/U42  ( .A1(cv_q[113]), .A2(rnd_q[113]), .ZN(\add_98_2/n40 )
         );
  OR2_X4 \add_98_2/U41  ( .A1(rnd_q[114]), .A2(cv_q[114]), .ZN(\add_98_2/n266 ) );
  NAND2_X1 \add_98_2/U40  ( .A1(cv_q[112]), .A2(rnd_q[112]), .ZN(
        \add_98_2/n277 ) );
  OR2_X4 \add_98_2/U39  ( .A1(rnd_q[118]), .A2(cv_q[118]), .ZN(\add_98_2/n199 ) );
  OR2_X4 \add_98_2/U38  ( .A1(rnd_q[115]), .A2(cv_q[115]), .ZN(\add_98_2/n196 ) );
  OR2_X4 \add_98_2/U37  ( .A1(rnd_q[111]), .A2(cv_q[111]), .ZN(\add_98_2/n300 ) );
  OR2_X4 \add_98_2/U36  ( .A1(rnd_q[107]), .A2(cv_q[107]), .ZN(\add_98_2/n308 ) );
  NOR2_X1 \add_98_2/U35  ( .A1(cv_q[108]), .A2(rnd_q[108]), .ZN(
        \add_98_2/n312 ) );
  NOR2_X1 \add_98_2/U34  ( .A1(rnd_q[100]), .A2(cv_q[100]), .ZN(\add_98_2/n36 ) );
  NOR2_X1 \add_98_2/U33  ( .A1(cv_q[105]), .A2(rnd_q[105]), .ZN(\add_98_2/n43 ) );
  NOR2_X1 \add_98_2/U32  ( .A1(cv_q[104]), .A2(rnd_q[104]), .ZN(\add_98_2/n46 ) );
  NOR2_X1 \add_98_2/U31  ( .A1(cv_q[110]), .A2(rnd_q[110]), .ZN(
        \add_98_2/n303 ) );
  NOR2_X1 \add_98_2/U30  ( .A1(cv_q[106]), .A2(rnd_q[106]), .ZN(
        \add_98_2/n343 ) );
  NOR2_X1 \add_98_2/U29  ( .A1(cv_q[109]), .A2(rnd_q[109]), .ZN(
        \add_98_2/n304 ) );
  AND2_X4 \add_98_2/U28  ( .A1(\add_98_2/n372 ), .A2(\add_98_2/n222 ), .ZN(N61) );
  AND2_X4 \add_98_2/U27  ( .A1(\add_98_2/n199 ), .A2(\add_98_2/n204 ), .ZN(
        \add_98_2/n26 ) );
  AND2_X4 \add_98_2/U26  ( .A1(\add_98_2/n151 ), .A2(\add_98_2/n101 ), .ZN(
        \add_98_2/n25 ) );
  AND2_X4 \add_98_2/U25  ( .A1(\add_98_2/n159 ), .A2(\add_98_2/n162 ), .ZN(
        \add_98_2/n24 ) );
  AND2_X4 \add_98_2/U24  ( .A1(\add_98_2/n127 ), .A2(\add_98_2/n196 ), .ZN(
        \add_98_2/n23 ) );
  OR2_X4 \add_98_2/U23  ( .A1(\add_98_2/n304 ), .A2(\add_98_2/n322 ), .ZN(
        \add_98_2/n22 ) );
  OR2_X4 \add_98_2/U22  ( .A1(\add_98_2/n303 ), .A2(\add_98_2/n304 ), .ZN(
        \add_98_2/n21 ) );
  AND2_X4 \add_98_2/U21  ( .A1(\add_98_2/n109 ), .A2(\add_98_2/n110 ), .ZN(
        \add_98_2/n20 ) );
  AND2_X4 \add_98_2/U20  ( .A1(\add_98_2/n153 ), .A2(\add_98_2/n151 ), .ZN(
        \add_98_2/n19 ) );
  AND3_X4 \add_98_2/U19  ( .A1(\add_98_2/n30 ), .A2(\add_98_2/n150 ), .A3(
        \add_98_2/n163 ), .ZN(\add_98_2/n18 ) );
  OR2_X4 \add_98_2/U18  ( .A1(\add_98_2/n235 ), .A2(\add_98_2/n231 ), .ZN(
        \add_98_2/n17 ) );
  OR2_X4 \add_98_2/U17  ( .A1(\add_98_2/n343 ), .A2(\add_98_2/n344 ), .ZN(
        \add_98_2/n16 ) );
  AND2_X4 \add_98_2/U16  ( .A1(\add_98_2/n216 ), .A2(\add_98_2/n332 ), .ZN(
        \add_98_2/n15 ) );
  AND2_X4 \add_98_2/U15  ( .A1(\add_98_2/n103 ), .A2(\add_98_2/n104 ), .ZN(
        \add_98_2/n14 ) );
  AND3_X4 \add_98_2/U14  ( .A1(\add_98_2/n103 ), .A2(\add_98_2/n94 ), .A3(
        \add_98_2/n104 ), .ZN(\add_98_2/n13 ) );
  AND2_X4 \add_98_2/U13  ( .A1(\add_98_2/n149 ), .A2(\add_98_2/n104 ), .ZN(
        \add_98_2/n12 ) );
  OR2_X4 \add_98_2/U12  ( .A1(cv_q[110]), .A2(rnd_q[110]), .ZN(\add_98_2/n11 )
         );
  OR2_X4 \add_98_2/U11  ( .A1(\add_98_2/n178 ), .A2(\add_98_2/n179 ), .ZN(
        \add_98_2/n10 ) );
  AND2_X4 \add_98_2/U10  ( .A1(\add_98_2/n364 ), .A2(\add_98_2/n3 ), .ZN(
        \add_98_2/n9 ) );
  OR2_X4 \add_98_2/U9  ( .A1(cv_q[99]), .A2(rnd_q[99]), .ZN(\add_98_2/n8 ) );
  OR2_X4 \add_98_2/U8  ( .A1(cv_q[102]), .A2(rnd_q[102]), .ZN(\add_98_2/n7 )
         );
  OR2_X4 \add_98_2/U7  ( .A1(cv_q[109]), .A2(rnd_q[109]), .ZN(\add_98_2/n6 )
         );
  OR2_X4 \add_98_2/U6  ( .A1(cv_q[98]), .A2(rnd_q[98]), .ZN(\add_98_2/n5 ) );
  OR3_X4 \add_98_2/U5  ( .A1(\add_98_2/n320 ), .A2(\add_98_2/n9 ), .A3(
        \add_98_2/n321 ), .ZN(\add_98_2/n4 ) );
  OR2_X4 \add_98_2/U4  ( .A1(cv_q[103]), .A2(rnd_q[103]), .ZN(\add_98_2/n3 )
         );
  OR2_X4 \add_98_2/U3  ( .A1(cv_q[97]), .A2(rnd_q[97]), .ZN(\add_98_2/n2 ) );
  AND3_X4 \add_98_2/U2  ( .A1(\add_98_2/n5 ), .A2(\add_98_2/n8 ), .A3(
        \add_98_2/n2 ), .ZN(\add_98_2/n1 ) );
  NAND2_X2 \add_98_3/U413  ( .A1(rnd_q[64]), .A2(cv_q[64]), .ZN(
        \add_98_3/n222 ) );
  INV_X4 \add_98_3/U412  ( .A(\add_98_3/n345 ), .ZN(\add_98_3/n381 ) );
  NAND2_X2 \add_98_3/U411  ( .A1(rnd_q[74]), .A2(cv_q[74]), .ZN(
        \add_98_3/n344 ) );
  NAND2_X2 \add_98_3/U410  ( .A1(\add_98_3/n381 ), .A2(\add_98_3/n344 ), .ZN(
        \add_98_3/n361 ) );
  NAND2_X2 \add_98_3/U409  ( .A1(rnd_q[72]), .A2(cv_q[72]), .ZN(\add_98_3/n52 ) );
  NAND2_X2 \add_98_3/U408  ( .A1(rnd_q[65]), .A2(cv_q[65]), .ZN(
        \add_98_3/n377 ) );
  NAND2_X2 \add_98_3/U407  ( .A1(\add_98_3/n377 ), .A2(\add_98_3/n222 ), .ZN(
        \add_98_3/n376 ) );
  NAND2_X2 \add_98_3/U406  ( .A1(\add_98_3/n1 ), .A2(\add_98_3/n376 ), .ZN(
        \add_98_3/n372 ) );
  NAND2_X2 \add_98_3/U405  ( .A1(cv_q[66]), .A2(rnd_q[66]), .ZN(
        \add_98_3/n375 ) );
  INV_X4 \add_98_3/U404  ( .A(\add_98_3/n219 ), .ZN(\add_98_3/n373 ) );
  NAND2_X2 \add_98_3/U403  ( .A1(rnd_q[67]), .A2(cv_q[67]), .ZN(
        \add_98_3/n217 ) );
  INV_X4 \add_98_3/U402  ( .A(\add_98_3/n29 ), .ZN(\add_98_3/n371 ) );
  NAND2_X2 \add_98_3/U401  ( .A1(rnd_q[71]), .A2(cv_q[71]), .ZN(\add_98_3/n56 ) );
  NAND2_X2 \add_98_3/U400  ( .A1(rnd_q[70]), .A2(cv_q[70]), .ZN(
        \add_98_3/n370 ) );
  NAND2_X2 \add_98_3/U399  ( .A1(rnd_q[68]), .A2(cv_q[68]), .ZN(\add_98_3/n66 ) );
  NAND2_X2 \add_98_3/U398  ( .A1(rnd_q[69]), .A2(cv_q[69]), .ZN(\add_98_3/n63 ) );
  NAND2_X2 \add_98_3/U397  ( .A1(\add_98_3/n66 ), .A2(\add_98_3/n63 ), .ZN(
        \add_98_3/n369 ) );
  NAND2_X2 \add_98_3/U396  ( .A1(\add_98_3/n368 ), .A2(\add_98_3/n369 ), .ZN(
        \add_98_3/n367 ) );
  NAND2_X2 \add_98_3/U395  ( .A1(\add_98_3/n40 ), .A2(\add_98_3/n367 ), .ZN(
        \add_98_3/n366 ) );
  NAND2_X2 \add_98_3/U394  ( .A1(\add_98_3/n9 ), .A2(\add_98_3/n365 ), .ZN(
        \add_98_3/n364 ) );
  XNOR2_X2 \add_98_3/U393  ( .A(\add_98_3/n361 ), .B(\add_98_3/n360 ), .ZN(
        N103) );
  NAND2_X2 \add_98_3/U392  ( .A1(\add_98_3/n360 ), .A2(\add_98_3/n381 ), .ZN(
        \add_98_3/n359 ) );
  NAND2_X2 \add_98_3/U391  ( .A1(\add_98_3/n359 ), .A2(\add_98_3/n344 ), .ZN(
        \add_98_3/n357 ) );
  NAND2_X2 \add_98_3/U390  ( .A1(rnd_q[75]), .A2(cv_q[75]), .ZN(
        \add_98_3/n343 ) );
  NAND2_X2 \add_98_3/U389  ( .A1(\add_98_3/n343 ), .A2(\add_98_3/n310 ), .ZN(
        \add_98_3/n358 ) );
  XNOR2_X2 \add_98_3/U388  ( .A(\add_98_3/n357 ), .B(\add_98_3/n358 ), .ZN(
        N104) );
  INV_X4 \add_98_3/U387  ( .A(\add_98_3/n43 ), .ZN(\add_98_3/n352 ) );
  INV_X4 \add_98_3/U386  ( .A(\add_98_3/n46 ), .ZN(\add_98_3/n353 ) );
  INV_X4 \add_98_3/U385  ( .A(\add_98_3/n310 ), .ZN(\add_98_3/n355 ) );
  NAND2_X2 \add_98_3/U384  ( .A1(\add_98_3/n347 ), .A2(\add_98_3/n348 ), .ZN(
        \add_98_3/n339 ) );
  NAND2_X2 \add_98_3/U383  ( .A1(cv_q[73]), .A2(rnd_q[73]), .ZN(
        \add_98_3/n346 ) );
  INV_X4 \add_98_3/U382  ( .A(\add_98_3/n344 ), .ZN(\add_98_3/n341 ) );
  INV_X4 \add_98_3/U381  ( .A(\add_98_3/n343 ), .ZN(\add_98_3/n342 ) );
  NAND2_X2 \add_98_3/U380  ( .A1(\add_98_3/n311 ), .A2(\add_98_3/n310 ), .ZN(
        \add_98_3/n334 ) );
  INV_X4 \add_98_3/U379  ( .A(\add_98_3/n334 ), .ZN(\add_98_3/n323 ) );
  NAND2_X2 \add_98_3/U378  ( .A1(rnd_q[76]), .A2(cv_q[76]), .ZN(
        \add_98_3/n324 ) );
  INV_X4 \add_98_3/U377  ( .A(\add_98_3/n324 ), .ZN(\add_98_3/n337 ) );
  XNOR2_X2 \add_98_3/U376  ( .A(\add_98_3/n335 ), .B(\add_98_3/n336 ), .ZN(
        N105) );
  NAND2_X2 \add_98_3/U375  ( .A1(\add_98_3/n330 ), .A2(\add_98_3/n5 ), .ZN(
        \add_98_3/n333 ) );
  NAND2_X2 \add_98_3/U374  ( .A1(\add_98_3/n333 ), .A2(\add_98_3/n324 ), .ZN(
        \add_98_3/n331 ) );
  NAND2_X2 \add_98_3/U373  ( .A1(rnd_q[77]), .A2(cv_q[77]), .ZN(
        \add_98_3/n325 ) );
  NAND2_X2 \add_98_3/U372  ( .A1(\add_98_3/n325 ), .A2(\add_98_3/n6 ), .ZN(
        \add_98_3/n332 ) );
  XNOR2_X2 \add_98_3/U371  ( .A(\add_98_3/n331 ), .B(\add_98_3/n332 ), .ZN(
        N106) );
  NAND2_X2 \add_98_3/U370  ( .A1(rnd_q[78]), .A2(cv_q[78]), .ZN(
        \add_98_3/n326 ) );
  NAND2_X2 \add_98_3/U369  ( .A1(\add_98_3/n11 ), .A2(\add_98_3/n326 ), .ZN(
        \add_98_3/n328 ) );
  XNOR2_X2 \add_98_3/U368  ( .A(\add_98_3/n327 ), .B(\add_98_3/n328 ), .ZN(
        N107) );
  INV_X4 \add_98_3/U367  ( .A(\add_98_3/n302 ), .ZN(\add_98_3/n313 ) );
  INV_X4 \add_98_3/U366  ( .A(\add_98_3/n326 ), .ZN(\add_98_3/n308 ) );
  NAND2_X2 \add_98_3/U365  ( .A1(\add_98_3/n324 ), .A2(\add_98_3/n325 ), .ZN(
        \add_98_3/n321 ) );
  XNOR2_X2 \add_98_3/U364  ( .A(\add_98_3/n315 ), .B(\add_98_3/n316 ), .ZN(
        N108) );
  NAND2_X2 \add_98_3/U363  ( .A1(rnd_q[80]), .A2(cv_q[80]), .ZN(
        \add_98_3/n282 ) );
  NAND2_X2 \add_98_3/U362  ( .A1(\add_98_3/n282 ), .A2(\add_98_3/n284 ), .ZN(
        \add_98_3/n285 ) );
  INV_X4 \add_98_3/U361  ( .A(\add_98_3/n133 ), .ZN(\add_98_3/n211 ) );
  NAND2_X2 \add_98_3/U360  ( .A1(cv_q[77]), .A2(rnd_q[77]), .ZN(
        \add_98_3/n309 ) );
  NAND2_X2 \add_98_3/U359  ( .A1(rnd_q[76]), .A2(cv_q[76]), .ZN(
        \add_98_3/n304 ) );
  NAND2_X2 \add_98_3/U358  ( .A1(\add_98_3/n301 ), .A2(\add_98_3/n302 ), .ZN(
        \add_98_3/n132 ) );
  INV_X4 \add_98_3/U357  ( .A(\add_98_3/n132 ), .ZN(\add_98_3/n210 ) );
  INV_X4 \add_98_3/U356  ( .A(\add_98_3/n222 ), .ZN(\add_98_3/n300 ) );
  NAND2_X2 \add_98_3/U355  ( .A1(rnd_q[65]), .A2(cv_q[65]), .ZN(
        \add_98_3/n138 ) );
  INV_X4 \add_98_3/U354  ( .A(\add_98_3/n138 ), .ZN(\add_98_3/n262 ) );
  INV_X4 \add_98_3/U353  ( .A(\add_98_3/n217 ), .ZN(\add_98_3/n77 ) );
  NAND2_X2 \add_98_3/U352  ( .A1(\add_98_3/n298 ), .A2(\add_98_3/n299 ), .ZN(
        \add_98_3/n295 ) );
  NAND2_X2 \add_98_3/U351  ( .A1(rnd_q[69]), .A2(cv_q[69]), .ZN(
        \add_98_3/n291 ) );
  NAND2_X2 \add_98_3/U350  ( .A1(\add_98_3/n66 ), .A2(\add_98_3/n291 ), .ZN(
        \add_98_3/n290 ) );
  NAND2_X2 \add_98_3/U349  ( .A1(\add_98_3/n227 ), .A2(\add_98_3/n290 ), .ZN(
        \add_98_3/n289 ) );
  NAND2_X2 \add_98_3/U348  ( .A1(\add_98_3/n40 ), .A2(\add_98_3/n289 ), .ZN(
        \add_98_3/n287 ) );
  NAND3_X2 \add_98_3/U347  ( .A1(\add_98_3/n287 ), .A2(\add_98_3/n3 ), .A3(
        \add_98_3/n288 ), .ZN(\add_98_3/n260 ) );
  INV_X4 \add_98_3/U346  ( .A(\add_98_3/n260 ), .ZN(\add_98_3/n135 ) );
  XNOR2_X2 \add_98_3/U345  ( .A(\add_98_3/n285 ), .B(\add_98_3/n88 ), .ZN(N109) );
  INV_X4 \add_98_3/U344  ( .A(\add_98_3/n276 ), .ZN(\add_98_3/n284 ) );
  NAND2_X2 \add_98_3/U343  ( .A1(\add_98_3/n88 ), .A2(\add_98_3/n284 ), .ZN(
        \add_98_3/n283 ) );
  NAND2_X2 \add_98_3/U342  ( .A1(\add_98_3/n282 ), .A2(\add_98_3/n283 ), .ZN(
        \add_98_3/n280 ) );
  NAND2_X2 \add_98_3/U341  ( .A1(rnd_q[81]), .A2(cv_q[81]), .ZN(
        \add_98_3/n277 ) );
  NAND2_X2 \add_98_3/U340  ( .A1(\add_98_3/n33 ), .A2(\add_98_3/n277 ), .ZN(
        \add_98_3/n281 ) );
  XNOR2_X2 \add_98_3/U339  ( .A(\add_98_3/n280 ), .B(\add_98_3/n281 ), .ZN(
        N110) );
  NAND2_X2 \add_98_3/U338  ( .A1(\add_98_3/n39 ), .A2(\add_98_3/n277 ), .ZN(
        \add_98_3/n267 ) );
  INV_X4 \add_98_3/U337  ( .A(\add_98_3/n267 ), .ZN(\add_98_3/n273 ) );
  NAND2_X2 \add_98_3/U336  ( .A1(\add_98_3/n270 ), .A2(\add_98_3/n88 ), .ZN(
        \add_98_3/n274 ) );
  NAND2_X2 \add_98_3/U335  ( .A1(\add_98_3/n273 ), .A2(\add_98_3/n274 ), .ZN(
        \add_98_3/n271 ) );
  NAND2_X2 \add_98_3/U334  ( .A1(rnd_q[82]), .A2(cv_q[82]), .ZN(
        \add_98_3/n266 ) );
  NAND2_X2 \add_98_3/U333  ( .A1(\add_98_3/n266 ), .A2(\add_98_3/n268 ), .ZN(
        \add_98_3/n272 ) );
  XNOR2_X2 \add_98_3/U332  ( .A(\add_98_3/n271 ), .B(\add_98_3/n272 ), .ZN(
        N111) );
  INV_X4 \add_98_3/U331  ( .A(\add_98_3/n88 ), .ZN(\add_98_3/n269 ) );
  NAND2_X2 \add_98_3/U330  ( .A1(\add_98_3/n270 ), .A2(\add_98_3/n268 ), .ZN(
        \add_98_3/n258 ) );
  NAND2_X2 \add_98_3/U329  ( .A1(\add_98_3/n267 ), .A2(\add_98_3/n268 ), .ZN(
        \add_98_3/n265 ) );
  NAND2_X2 \add_98_3/U328  ( .A1(\add_98_3/n265 ), .A2(\add_98_3/n266 ), .ZN(
        \add_98_3/n197 ) );
  NAND2_X2 \add_98_3/U327  ( .A1(rnd_q[83]), .A2(cv_q[83]), .ZN(
        \add_98_3/n127 ) );
  XNOR2_X2 \add_98_3/U326  ( .A(\add_98_3/n263 ), .B(\add_98_3/n23 ), .ZN(N112) );
  XNOR2_X2 \add_98_3/U325  ( .A(\add_98_3/n222 ), .B(\add_98_3/n261 ), .ZN(N94) );
  INV_X4 \add_98_3/U324  ( .A(\add_98_3/n258 ), .ZN(\add_98_3/n257 ) );
  NAND2_X2 \add_98_3/U323  ( .A1(\add_98_3/n257 ), .A2(\add_98_3/n196 ), .ZN(
        \add_98_3/n129 ) );
  NAND2_X2 \add_98_3/U322  ( .A1(\add_98_3/n197 ), .A2(\add_98_3/n196 ), .ZN(
        \add_98_3/n126 ) );
  NAND2_X2 \add_98_3/U321  ( .A1(\add_98_3/n126 ), .A2(\add_98_3/n127 ), .ZN(
        \add_98_3/n255 ) );
  XNOR2_X2 \add_98_3/U320  ( .A(\add_98_3/n237 ), .B(\add_98_3/n253 ), .ZN(
        N113) );
  NAND2_X2 \add_98_3/U319  ( .A1(rnd_q[85]), .A2(cv_q[85]), .ZN(
        \add_98_3/n202 ) );
  INV_X4 \add_98_3/U318  ( .A(\add_98_3/n202 ), .ZN(\add_98_3/n250 ) );
  XNOR2_X2 \add_98_3/U317  ( .A(\add_98_3/n248 ), .B(\add_98_3/n249 ), .ZN(
        N114) );
  INV_X4 \add_98_3/U316  ( .A(\add_98_3/n238 ), .ZN(\add_98_3/n245 ) );
  INV_X4 \add_98_3/U315  ( .A(\add_98_3/n244 ), .ZN(\add_98_3/n243 ) );
  NAND2_X2 \add_98_3/U314  ( .A1(\add_98_3/n203 ), .A2(\add_98_3/n202 ), .ZN(
        \add_98_3/n242 ) );
  NAND2_X2 \add_98_3/U313  ( .A1(rnd_q[86]), .A2(cv_q[86]), .ZN(
        \add_98_3/n204 ) );
  XNOR2_X2 \add_98_3/U312  ( .A(\add_98_3/n240 ), .B(\add_98_3/n26 ), .ZN(N115) );
  NAND2_X2 \add_98_3/U311  ( .A1(\add_98_3/n203 ), .A2(\add_98_3/n202 ), .ZN(
        \add_98_3/n239 ) );
  NAND2_X2 \add_98_3/U310  ( .A1(\add_98_3/n239 ), .A2(\add_98_3/n199 ), .ZN(
        \add_98_3/n236 ) );
  NAND2_X2 \add_98_3/U309  ( .A1(\add_98_3/n238 ), .A2(\add_98_3/n199 ), .ZN(
        \add_98_3/n231 ) );
  INV_X4 \add_98_3/U308  ( .A(rnd_q[87]), .ZN(\add_98_3/n234 ) );
  INV_X4 \add_98_3/U307  ( .A(cv_q[87]), .ZN(\add_98_3/n235 ) );
  NAND2_X2 \add_98_3/U306  ( .A1(\add_98_3/n234 ), .A2(\add_98_3/n235 ), .ZN(
        \add_98_3/n200 ) );
  NAND2_X2 \add_98_3/U305  ( .A1(rnd_q[87]), .A2(cv_q[87]), .ZN(
        \add_98_3/n152 ) );
  NAND2_X2 \add_98_3/U304  ( .A1(\add_98_3/n200 ), .A2(\add_98_3/n152 ), .ZN(
        \add_98_3/n233 ) );
  XNOR2_X2 \add_98_3/U303  ( .A(\add_98_3/n232 ), .B(\add_98_3/n233 ), .ZN(
        N116) );
  INV_X4 \add_98_3/U302  ( .A(\add_98_3/n231 ), .ZN(\add_98_3/n230 ) );
  NAND2_X2 \add_98_3/U301  ( .A1(\add_98_3/n230 ), .A2(\add_98_3/n200 ), .ZN(
        \add_98_3/n147 ) );
  NAND2_X2 \add_98_3/U300  ( .A1(rnd_q[69]), .A2(cv_q[69]), .ZN(
        \add_98_3/n229 ) );
  NAND2_X2 \add_98_3/U299  ( .A1(\add_98_3/n66 ), .A2(\add_98_3/n229 ), .ZN(
        \add_98_3/n228 ) );
  NAND2_X2 \add_98_3/U298  ( .A1(\add_98_3/n227 ), .A2(\add_98_3/n228 ), .ZN(
        \add_98_3/n226 ) );
  NAND2_X2 \add_98_3/U297  ( .A1(\add_98_3/n40 ), .A2(\add_98_3/n226 ), .ZN(
        \add_98_3/n223 ) );
  INV_X4 \add_98_3/U296  ( .A(\add_98_3/n215 ), .ZN(\add_98_3/n224 ) );
  INV_X4 \add_98_3/U295  ( .A(\add_98_3/n216 ), .ZN(\add_98_3/n225 ) );
  NAND4_X2 \add_98_3/U294  ( .A1(\add_98_3/n223 ), .A2(\add_98_3/n3 ), .A3(
        \add_98_3/n224 ), .A4(\add_98_3/n225 ), .ZN(\add_98_3/n207 ) );
  NAND2_X2 \add_98_3/U293  ( .A1(rnd_q[65]), .A2(cv_q[65]), .ZN(
        \add_98_3/n221 ) );
  NAND2_X2 \add_98_3/U292  ( .A1(\add_98_3/n221 ), .A2(\add_98_3/n222 ), .ZN(
        \add_98_3/n220 ) );
  NAND2_X2 \add_98_3/U291  ( .A1(\add_98_3/n1 ), .A2(\add_98_3/n220 ), .ZN(
        \add_98_3/n218 ) );
  INV_X4 \add_98_3/U290  ( .A(\add_98_3/n49 ), .ZN(\add_98_3/n214 ) );
  NAND2_X2 \add_98_3/U289  ( .A1(\add_98_3/n205 ), .A2(\add_98_3/n206 ), .ZN(
        \add_98_3/n189 ) );
  INV_X4 \add_98_3/U288  ( .A(\add_98_3/n146 ), .ZN(\add_98_3/n198 ) );
  NAND2_X2 \add_98_3/U287  ( .A1(\add_98_3/n198 ), .A2(\add_98_3/n152 ), .ZN(
        \add_98_3/n191 ) );
  INV_X4 \add_98_3/U286  ( .A(\add_98_3/n197 ), .ZN(\add_98_3/n194 ) );
  INV_X4 \add_98_3/U285  ( .A(\add_98_3/n196 ), .ZN(\add_98_3/n195 ) );
  NAND2_X2 \add_98_3/U284  ( .A1(\add_98_3/n189 ), .A2(\add_98_3/n190 ), .ZN(
        \add_98_3/n163 ) );
  NAND2_X2 \add_98_3/U283  ( .A1(rnd_q[88]), .A2(cv_q[88]), .ZN(
        \add_98_3/n187 ) );
  NAND2_X2 \add_98_3/U282  ( .A1(\add_98_3/n187 ), .A2(\add_98_3/n172 ), .ZN(
        \add_98_3/n188 ) );
  XNOR2_X2 \add_98_3/U281  ( .A(\add_98_3/n163 ), .B(\add_98_3/n188 ), .ZN(
        N117) );
  INV_X4 \add_98_3/U280  ( .A(\add_98_3/n181 ), .ZN(\add_98_3/n172 ) );
  NAND2_X2 \add_98_3/U279  ( .A1(\add_98_3/n172 ), .A2(\add_98_3/n163 ), .ZN(
        \add_98_3/n186 ) );
  NAND2_X2 \add_98_3/U278  ( .A1(\add_98_3/n186 ), .A2(\add_98_3/n187 ), .ZN(
        \add_98_3/n182 ) );
  NAND2_X2 \add_98_3/U277  ( .A1(rnd_q[89]), .A2(cv_q[89]), .ZN(
        \add_98_3/n161 ) );
  INV_X4 \add_98_3/U276  ( .A(rnd_q[89]), .ZN(\add_98_3/n184 ) );
  INV_X4 \add_98_3/U275  ( .A(cv_q[89]), .ZN(\add_98_3/n185 ) );
  NAND2_X2 \add_98_3/U274  ( .A1(\add_98_3/n184 ), .A2(\add_98_3/n185 ), .ZN(
        \add_98_3/n171 ) );
  NAND2_X2 \add_98_3/U273  ( .A1(\add_98_3/n161 ), .A2(\add_98_3/n171 ), .ZN(
        \add_98_3/n183 ) );
  XNOR2_X2 \add_98_3/U272  ( .A(\add_98_3/n182 ), .B(\add_98_3/n183 ), .ZN(
        N118) );
  INV_X4 \add_98_3/U271  ( .A(\add_98_3/n163 ), .ZN(\add_98_3/n180 ) );
  INV_X4 \add_98_3/U270  ( .A(\add_98_3/n171 ), .ZN(\add_98_3/n178 ) );
  NAND2_X2 \add_98_3/U269  ( .A1(cv_q[88]), .A2(rnd_q[88]), .ZN(
        \add_98_3/n179 ) );
  NAND2_X2 \add_98_3/U268  ( .A1(\add_98_3/n10 ), .A2(\add_98_3/n161 ), .ZN(
        \add_98_3/n177 ) );
  INV_X4 \add_98_3/U267  ( .A(rnd_q[90]), .ZN(\add_98_3/n174 ) );
  INV_X4 \add_98_3/U266  ( .A(cv_q[90]), .ZN(\add_98_3/n175 ) );
  NAND2_X2 \add_98_3/U265  ( .A1(\add_98_3/n174 ), .A2(\add_98_3/n175 ), .ZN(
        \add_98_3/n159 ) );
  NAND2_X2 \add_98_3/U264  ( .A1(rnd_q[90]), .A2(cv_q[90]), .ZN(
        \add_98_3/n162 ) );
  XNOR2_X2 \add_98_3/U263  ( .A(\add_98_3/n173 ), .B(\add_98_3/n24 ), .ZN(N119) );
  NAND2_X2 \add_98_3/U262  ( .A1(\add_98_3/n30 ), .A2(\add_98_3/n163 ), .ZN(
        \add_98_3/n168 ) );
  NAND2_X2 \add_98_3/U261  ( .A1(\add_98_3/n170 ), .A2(\add_98_3/n159 ), .ZN(
        \add_98_3/n169 ) );
  NAND2_X2 \add_98_3/U260  ( .A1(\add_98_3/n168 ), .A2(\add_98_3/n169 ), .ZN(
        \add_98_3/n164 ) );
  INV_X4 \add_98_3/U259  ( .A(rnd_q[91]), .ZN(\add_98_3/n166 ) );
  INV_X4 \add_98_3/U258  ( .A(cv_q[91]), .ZN(\add_98_3/n167 ) );
  NAND2_X2 \add_98_3/U257  ( .A1(\add_98_3/n166 ), .A2(\add_98_3/n167 ), .ZN(
        \add_98_3/n150 ) );
  NAND2_X2 \add_98_3/U256  ( .A1(rnd_q[91]), .A2(cv_q[91]), .ZN(
        \add_98_3/n158 ) );
  NAND2_X2 \add_98_3/U255  ( .A1(\add_98_3/n150 ), .A2(\add_98_3/n158 ), .ZN(
        \add_98_3/n165 ) );
  XNOR2_X2 \add_98_3/U254  ( .A(\add_98_3/n164 ), .B(\add_98_3/n165 ), .ZN(
        N120) );
  NAND2_X2 \add_98_3/U253  ( .A1(\add_98_3/n157 ), .A2(\add_98_3/n158 ), .ZN(
        \add_98_3/n153 ) );
  INV_X4 \add_98_3/U252  ( .A(rnd_q[92]), .ZN(\add_98_3/n155 ) );
  INV_X4 \add_98_3/U251  ( .A(cv_q[92]), .ZN(\add_98_3/n156 ) );
  NAND2_X2 \add_98_3/U250  ( .A1(\add_98_3/n155 ), .A2(\add_98_3/n156 ), .ZN(
        \add_98_3/n151 ) );
  NAND2_X2 \add_98_3/U249  ( .A1(rnd_q[92]), .A2(cv_q[92]), .ZN(
        \add_98_3/n101 ) );
  XNOR2_X2 \add_98_3/U248  ( .A(\add_98_3/n154 ), .B(\add_98_3/n25 ), .ZN(N121) );
  INV_X4 \add_98_3/U247  ( .A(\add_98_3/n152 ), .ZN(\add_98_3/n149 ) );
  INV_X4 \add_98_3/U246  ( .A(\add_98_3/n122 ), .ZN(\add_98_3/n104 ) );
  INV_X4 \add_98_3/U245  ( .A(\add_98_3/n101 ), .ZN(\add_98_3/n148 ) );
  INV_X4 \add_98_3/U244  ( .A(\add_98_3/n147 ), .ZN(\add_98_3/n103 ) );
  INV_X4 \add_98_3/U243  ( .A(\add_98_3/n129 ), .ZN(\add_98_3/n87 ) );
  NAND2_X2 \add_98_3/U242  ( .A1(\add_98_3/n126 ), .A2(\add_98_3/n127 ), .ZN(
        \add_98_3/n102 ) );
  NAND2_X2 \add_98_3/U241  ( .A1(\add_98_3/n102 ), .A2(\add_98_3/n14 ), .ZN(
        \add_98_3/n145 ) );
  NAND2_X2 \add_98_3/U240  ( .A1(\add_98_3/n146 ), .A2(\add_98_3/n104 ), .ZN(
        \add_98_3/n93 ) );
  NAND4_X2 \add_98_3/U239  ( .A1(\add_98_3/n143 ), .A2(\add_98_3/n144 ), .A3(
        \add_98_3/n145 ), .A4(\add_98_3/n93 ), .ZN(\add_98_3/n139 ) );
  NAND2_X2 \add_98_3/U238  ( .A1(rnd_q[93]), .A2(cv_q[93]), .ZN(\add_98_3/n91 ) );
  INV_X4 \add_98_3/U237  ( .A(rnd_q[93]), .ZN(\add_98_3/n141 ) );
  INV_X4 \add_98_3/U236  ( .A(cv_q[93]), .ZN(\add_98_3/n142 ) );
  NAND2_X2 \add_98_3/U235  ( .A1(\add_98_3/n141 ), .A2(\add_98_3/n142 ), .ZN(
        \add_98_3/n117 ) );
  NAND2_X2 \add_98_3/U234  ( .A1(\add_98_3/n91 ), .A2(\add_98_3/n117 ), .ZN(
        \add_98_3/n140 ) );
  XNOR2_X2 \add_98_3/U233  ( .A(\add_98_3/n139 ), .B(\add_98_3/n140 ), .ZN(
        N122) );
  XNOR2_X2 \add_98_3/U232  ( .A(\add_98_3/n80 ), .B(\add_98_3/n136 ), .ZN(N95)
         );
  INV_X4 \add_98_3/U231  ( .A(\add_98_3/n134 ), .ZN(\add_98_3/n130 ) );
  NAND2_X2 \add_98_3/U230  ( .A1(\add_98_3/n132 ), .A2(\add_98_3/n133 ), .ZN(
        \add_98_3/n131 ) );
  NAND2_X2 \add_98_3/U229  ( .A1(\add_98_3/n126 ), .A2(\add_98_3/n127 ), .ZN(
        \add_98_3/n125 ) );
  NAND2_X2 \add_98_3/U228  ( .A1(\add_98_3/n103 ), .A2(\add_98_3/n117 ), .ZN(
        \add_98_3/n123 ) );
  NAND2_X2 \add_98_3/U227  ( .A1(\add_98_3/n12 ), .A2(\add_98_3/n117 ), .ZN(
        \add_98_3/n113 ) );
  INV_X4 \add_98_3/U226  ( .A(\add_98_3/n93 ), .ZN(\add_98_3/n120 ) );
  NAND2_X2 \add_98_3/U225  ( .A1(\add_98_3/n120 ), .A2(\add_98_3/n117 ), .ZN(
        \add_98_3/n114 ) );
  INV_X4 \add_98_3/U224  ( .A(\add_98_3/n91 ), .ZN(\add_98_3/n118 ) );
  INV_X4 \add_98_3/U223  ( .A(\add_98_3/n117 ), .ZN(\add_98_3/n105 ) );
  NAND2_X2 \add_98_3/U222  ( .A1(\add_98_3/n19 ), .A2(\add_98_3/n117 ), .ZN(
        \add_98_3/n116 ) );
  NAND4_X2 \add_98_3/U221  ( .A1(\add_98_3/n113 ), .A2(\add_98_3/n114 ), .A3(
        \add_98_3/n115 ), .A4(\add_98_3/n116 ), .ZN(\add_98_3/n112 ) );
  INV_X4 \add_98_3/U220  ( .A(rnd_q[94]), .ZN(\add_98_3/n109 ) );
  INV_X4 \add_98_3/U219  ( .A(cv_q[94]), .ZN(\add_98_3/n110 ) );
  NAND2_X2 \add_98_3/U218  ( .A1(rnd_q[94]), .A2(cv_q[94]), .ZN(
        \add_98_3/n100 ) );
  INV_X4 \add_98_3/U217  ( .A(\add_98_3/n100 ), .ZN(\add_98_3/n108 ) );
  XNOR2_X2 \add_98_3/U216  ( .A(\add_98_3/n106 ), .B(\add_98_3/n107 ), .ZN(
        N123) );
  NAND2_X2 \add_98_3/U215  ( .A1(\add_98_3/n13 ), .A2(\add_98_3/n102 ), .ZN(
        \add_98_3/n83 ) );
  NAND2_X2 \add_98_3/U214  ( .A1(\add_98_3/n94 ), .A2(\add_98_3/n148 ), .ZN(
        \add_98_3/n99 ) );
  NAND2_X2 \add_98_3/U213  ( .A1(\add_98_3/n99 ), .A2(\add_98_3/n100 ), .ZN(
        \add_98_3/n95 ) );
  NAND2_X2 \add_98_3/U212  ( .A1(\add_98_3/n12 ), .A2(\add_98_3/n94 ), .ZN(
        \add_98_3/n97 ) );
  NAND2_X2 \add_98_3/U211  ( .A1(\add_98_3/n19 ), .A2(\add_98_3/n94 ), .ZN(
        \add_98_3/n98 ) );
  NAND2_X2 \add_98_3/U210  ( .A1(\add_98_3/n97 ), .A2(\add_98_3/n98 ), .ZN(
        \add_98_3/n96 ) );
  INV_X4 \add_98_3/U209  ( .A(\add_98_3/n94 ), .ZN(\add_98_3/n92 ) );
  NAND4_X2 \add_98_3/U208  ( .A1(\add_98_3/n83 ), .A2(\add_98_3/n84 ), .A3(
        \add_98_3/n85 ), .A4(\add_98_3/n86 ), .ZN(\add_98_3/n81 ) );
  XNOR2_X2 \add_98_3/U207  ( .A(rnd_q[95]), .B(cv_q[95]), .ZN(\add_98_3/n82 )
         );
  XNOR2_X2 \add_98_3/U206  ( .A(\add_98_3/n81 ), .B(\add_98_3/n82 ), .ZN(N124)
         );
  XNOR2_X2 \add_98_3/U205  ( .A(\add_98_3/n74 ), .B(\add_98_3/n75 ), .ZN(N96)
         );
  INV_X4 \add_98_3/U204  ( .A(\add_98_3/n66 ), .ZN(\add_98_3/n72 ) );
  XNOR2_X2 \add_98_3/U203  ( .A(\add_98_3/n29 ), .B(\add_98_3/n73 ), .ZN(N97)
         );
  INV_X4 \add_98_3/U202  ( .A(\add_98_3/n63 ), .ZN(\add_98_3/n70 ) );
  XNOR2_X2 \add_98_3/U201  ( .A(\add_98_3/n68 ), .B(\add_98_3/n69 ), .ZN(N98)
         );
  NAND2_X2 \add_98_3/U200  ( .A1(rnd_q[70]), .A2(cv_q[70]), .ZN(\add_98_3/n58 ) );
  NAND2_X2 \add_98_3/U199  ( .A1(\add_98_3/n58 ), .A2(\add_98_3/n7 ), .ZN(
        \add_98_3/n61 ) );
  NAND2_X2 \add_98_3/U198  ( .A1(\add_98_3/n29 ), .A2(\add_98_3/n66 ), .ZN(
        \add_98_3/n65 ) );
  NAND2_X2 \add_98_3/U197  ( .A1(\add_98_3/n64 ), .A2(\add_98_3/n65 ), .ZN(
        \add_98_3/n62 ) );
  NAND2_X2 \add_98_3/U196  ( .A1(\add_98_3/n62 ), .A2(\add_98_3/n63 ), .ZN(
        \add_98_3/n59 ) );
  XNOR2_X2 \add_98_3/U195  ( .A(\add_98_3/n61 ), .B(\add_98_3/n59 ), .ZN(N99)
         );
  NAND2_X2 \add_98_3/U194  ( .A1(\add_98_3/n59 ), .A2(\add_98_3/n7 ), .ZN(
        \add_98_3/n57 ) );
  NAND2_X2 \add_98_3/U193  ( .A1(\add_98_3/n57 ), .A2(\add_98_3/n58 ), .ZN(
        \add_98_3/n54 ) );
  NAND2_X2 \add_98_3/U192  ( .A1(\add_98_3/n56 ), .A2(\add_98_3/n3 ), .ZN(
        \add_98_3/n55 ) );
  XNOR2_X2 \add_98_3/U191  ( .A(\add_98_3/n54 ), .B(\add_98_3/n55 ), .ZN(N100)
         );
  INV_X4 \add_98_3/U190  ( .A(\add_98_3/n52 ), .ZN(\add_98_3/n45 ) );
  XNOR2_X2 \add_98_3/U189  ( .A(\add_98_3/n50 ), .B(\add_98_3/n51 ), .ZN(N101)
         );
  XNOR2_X2 \add_98_3/U188  ( .A(\add_98_3/n41 ), .B(\add_98_3/n42 ), .ZN(N102)
         );
  NAND2_X2 \add_98_3/U187  ( .A1(\add_98_3/n260 ), .A2(\add_98_3/n134 ), .ZN(
        \add_98_3/n259 ) );
  NOR2_X2 \add_98_3/U186  ( .A1(\add_98_3/n313 ), .A2(\add_98_3/n38 ), .ZN(
        \add_98_3/n315 ) );
  NOR2_X2 \add_98_3/U185  ( .A1(\add_98_3/n70 ), .A2(\add_98_3/n67 ), .ZN(
        \add_98_3/n69 ) );
  NOR2_X2 \add_98_3/U184  ( .A1(\add_98_3/n34 ), .A2(\add_98_3/n72 ), .ZN(
        \add_98_3/n73 ) );
  NOR2_X2 \add_98_3/U183  ( .A1(\add_98_3/n36 ), .A2(\add_98_3/n79 ), .ZN(
        \add_98_3/n136 ) );
  AND2_X2 \add_98_3/U182  ( .A1(cv_q[72]), .A2(rnd_q[72]), .ZN(\add_98_3/n347 ) );
  AND2_X2 \add_98_3/U181  ( .A1(\add_98_3/n56 ), .A2(\add_98_3/n370 ), .ZN(
        \add_98_3/n40 ) );
  NOR2_X2 \add_98_3/U180  ( .A1(\add_98_3/n20 ), .A2(\add_98_3/n108 ), .ZN(
        \add_98_3/n107 ) );
  NOR2_X2 \add_98_3/U179  ( .A1(\add_98_3/n244 ), .A2(\add_98_3/n250 ), .ZN(
        \add_98_3/n249 ) );
  NOR2_X2 \add_98_3/U178  ( .A1(\add_98_3/n46 ), .A2(\add_98_3/n45 ), .ZN(
        \add_98_3/n51 ) );
  NOR2_X2 \add_98_3/U177  ( .A1(\add_98_3/n76 ), .A2(\add_98_3/n77 ), .ZN(
        \add_98_3/n75 ) );
  NOR2_X2 \add_98_3/U176  ( .A1(\add_98_3/n262 ), .A2(\add_98_3/n137 ), .ZN(
        \add_98_3/n261 ) );
  OR2_X2 \add_98_3/U175  ( .A1(\add_98_3/n278 ), .A2(\add_98_3/n279 ), .ZN(
        \add_98_3/n39 ) );
  AND2_X2 \add_98_3/U174  ( .A1(rnd_q[79]), .A2(cv_q[79]), .ZN(\add_98_3/n38 )
         );
  AND2_X2 \add_98_3/U173  ( .A1(rnd_q[73]), .A2(cv_q[73]), .ZN(\add_98_3/n37 )
         );
  AND2_X2 \add_98_3/U172  ( .A1(rnd_q[66]), .A2(cv_q[66]), .ZN(\add_98_3/n36 )
         );
  AND2_X2 \add_98_3/U171  ( .A1(rnd_q[84]), .A2(cv_q[84]), .ZN(\add_98_3/n35 )
         );
  NOR2_X2 \add_98_3/U170  ( .A1(\add_98_3/n275 ), .A2(\add_98_3/n276 ), .ZN(
        \add_98_3/n270 ) );
  NOR2_X1 \add_98_3/U169  ( .A1(cv_q[73]), .A2(rnd_q[73]), .ZN(\add_98_3/n349 ) );
  NOR2_X1 \add_98_3/U168  ( .A1(cv_q[74]), .A2(rnd_q[74]), .ZN(\add_98_3/n350 ) );
  NOR2_X2 \add_98_3/U167  ( .A1(\add_98_3/n349 ), .A2(\add_98_3/n350 ), .ZN(
        \add_98_3/n348 ) );
  NOR2_X2 \add_98_3/U166  ( .A1(\add_98_3/n246 ), .A2(\add_98_3/n247 ), .ZN(
        \add_98_3/n238 ) );
  NOR2_X2 \add_98_3/U165  ( .A1(\add_98_3/n35 ), .A2(\add_98_3/n252 ), .ZN(
        \add_98_3/n253 ) );
  NOR2_X2 \add_98_3/U164  ( .A1(\add_98_3/n337 ), .A2(\add_98_3/n314 ), .ZN(
        \add_98_3/n336 ) );
  NOR2_X2 \add_98_3/U163  ( .A1(\add_98_3/n37 ), .A2(\add_98_3/n43 ), .ZN(
        \add_98_3/n42 ) );
  NOR2_X1 \add_98_3/U162  ( .A1(cv_q[69]), .A2(rnd_q[69]), .ZN(\add_98_3/n292 ) );
  NOR2_X1 \add_98_3/U161  ( .A1(cv_q[70]), .A2(rnd_q[70]), .ZN(\add_98_3/n293 ) );
  NOR2_X2 \add_98_3/U160  ( .A1(\add_98_3/n292 ), .A2(\add_98_3/n293 ), .ZN(
        \add_98_3/n227 ) );
  NOR2_X1 \add_98_3/U159  ( .A1(cv_q[69]), .A2(rnd_q[69]), .ZN(\add_98_3/n379 ) );
  NOR2_X1 \add_98_3/U158  ( .A1(cv_q[67]), .A2(rnd_q[67]), .ZN(\add_98_3/n76 )
         );
  NOR2_X1 \add_98_3/U157  ( .A1(cv_q[66]), .A2(rnd_q[66]), .ZN(\add_98_3/n79 )
         );
  NOR2_X2 \add_98_3/U156  ( .A1(cv_q[88]), .A2(rnd_q[88]), .ZN(\add_98_3/n181 ) );
  NOR2_X1 \add_98_3/U155  ( .A1(cv_q[70]), .A2(rnd_q[70]), .ZN(\add_98_3/n60 )
         );
  NOR2_X1 \add_98_3/U154  ( .A1(cv_q[69]), .A2(rnd_q[69]), .ZN(\add_98_3/n67 )
         );
  NOR2_X2 \add_98_3/U153  ( .A1(\add_98_3/n76 ), .A2(\add_98_3/n375 ), .ZN(
        \add_98_3/n219 ) );
  NOR2_X2 \add_98_3/U152  ( .A1(\add_98_3/n305 ), .A2(\add_98_3/n309 ), .ZN(
        \add_98_3/n307 ) );
  NOR3_X2 \add_98_3/U151  ( .A1(\add_98_3/n304 ), .A2(\add_98_3/n305 ), .A3(
        \add_98_3/n306 ), .ZN(\add_98_3/n303 ) );
  NAND3_X2 \add_98_3/U150  ( .A1(\add_98_3/n202 ), .A2(\add_98_3/n203 ), .A3(
        \add_98_3/n204 ), .ZN(\add_98_3/n201 ) );
  AND2_X4 \add_98_3/U149  ( .A1(\add_98_3/n199 ), .A2(\add_98_3/n200 ), .ZN(
        \add_98_3/n32 ) );
  AND2_X2 \add_98_3/U148  ( .A1(\add_98_3/n201 ), .A2(\add_98_3/n32 ), .ZN(
        \add_98_3/n146 ) );
  NOR2_X2 \add_98_3/U147  ( .A1(\add_98_3/n300 ), .A2(\add_98_3/n219 ), .ZN(
        \add_98_3/n298 ) );
  NAND3_X2 \add_98_3/U146  ( .A1(\add_98_3/n214 ), .A2(\add_98_3/n365 ), .A3(
        \add_98_3/n371 ), .ZN(\add_98_3/n363 ) );
  NOR2_X2 \add_98_3/U145  ( .A1(\add_98_3/n37 ), .A2(\add_98_3/n380 ), .ZN(
        \add_98_3/n362 ) );
  NAND3_X2 \add_98_3/U144  ( .A1(\add_98_3/n362 ), .A2(\add_98_3/n363 ), .A3(
        \add_98_3/n364 ), .ZN(\add_98_3/n360 ) );
  NAND3_X2 \add_98_3/U143  ( .A1(\add_98_3/n330 ), .A2(\add_98_3/n6 ), .A3(
        \add_98_3/n5 ), .ZN(\add_98_3/n329 ) );
  NAND3_X2 \add_98_3/U142  ( .A1(\add_98_3/n22 ), .A2(\add_98_3/n325 ), .A3(
        \add_98_3/n329 ), .ZN(\add_98_3/n327 ) );
  NOR2_X2 \add_98_3/U141  ( .A1(\add_98_3/n79 ), .A2(\add_98_3/n80 ), .ZN(
        \add_98_3/n78 ) );
  NOR2_X2 \add_98_3/U140  ( .A1(\add_98_3/n78 ), .A2(\add_98_3/n36 ), .ZN(
        \add_98_3/n74 ) );
  NOR2_X2 \add_98_3/U139  ( .A1(\add_98_3/n18 ), .A2(\add_98_3/n153 ), .ZN(
        \add_98_3/n154 ) );
  NOR2_X2 \add_98_3/U138  ( .A1(\add_98_3/n237 ), .A2(\add_98_3/n245 ), .ZN(
        \add_98_3/n241 ) );
  NOR2_X2 \add_98_3/U137  ( .A1(\add_98_3/n241 ), .A2(\add_98_3/n242 ), .ZN(
        \add_98_3/n240 ) );
  NOR2_X2 \add_98_3/U136  ( .A1(\add_98_3/n29 ), .A2(\add_98_3/n49 ), .ZN(
        \add_98_3/n48 ) );
  NOR2_X2 \add_98_3/U135  ( .A1(\add_98_3/n48 ), .A2(\add_98_3/n9 ), .ZN(
        \add_98_3/n47 ) );
  NOR2_X2 \add_98_3/U134  ( .A1(\add_98_3/n46 ), .A2(\add_98_3/n47 ), .ZN(
        \add_98_3/n44 ) );
  NOR2_X2 \add_98_3/U133  ( .A1(\add_98_3/n44 ), .A2(\add_98_3/n45 ), .ZN(
        \add_98_3/n41 ) );
  NOR2_X2 \add_98_3/U132  ( .A1(\add_98_3/n29 ), .A2(\add_98_3/n34 ), .ZN(
        \add_98_3/n71 ) );
  NOR2_X2 \add_98_3/U131  ( .A1(\add_98_3/n71 ), .A2(\add_98_3/n72 ), .ZN(
        \add_98_3/n68 ) );
  NOR3_X2 \add_98_3/U130  ( .A1(\add_98_3/n180 ), .A2(\add_98_3/n178 ), .A3(
        \add_98_3/n181 ), .ZN(\add_98_3/n176 ) );
  NOR2_X2 \add_98_3/U129  ( .A1(\add_98_3/n176 ), .A2(\add_98_3/n177 ), .ZN(
        \add_98_3/n173 ) );
  NOR2_X2 \add_98_3/U128  ( .A1(\add_98_3/n60 ), .A2(\add_98_3/n67 ), .ZN(
        \add_98_3/n368 ) );
  NOR2_X2 \add_98_3/U127  ( .A1(\add_98_3/n341 ), .A2(\add_98_3/n342 ), .ZN(
        \add_98_3/n340 ) );
  NAND3_X2 \add_98_3/U126  ( .A1(\add_98_3/n339 ), .A2(\add_98_3/n16 ), .A3(
        \add_98_3/n340 ), .ZN(\add_98_3/n311 ) );
  NOR2_X2 \add_98_3/U125  ( .A1(\add_98_3/n34 ), .A2(\add_98_3/n67 ), .ZN(
        \add_98_3/n64 ) );
  NOR2_X2 \add_98_3/U124  ( .A1(\add_98_3/n20 ), .A2(\add_98_3/n91 ), .ZN(
        \add_98_3/n90 ) );
  NOR2_X2 \add_98_3/U123  ( .A1(\add_98_3/n105 ), .A2(\add_98_3/n101 ), .ZN(
        \add_98_3/n119 ) );
  OR2_X4 \add_98_3/U122  ( .A1(\add_98_3/n137 ), .A2(\add_98_3/n222 ), .ZN(
        \add_98_3/n31 ) );
  AND2_X2 \add_98_3/U121  ( .A1(\add_98_3/n138 ), .A2(\add_98_3/n31 ), .ZN(
        \add_98_3/n80 ) );
  NOR2_X2 \add_98_3/U120  ( .A1(\add_98_3/n252 ), .A2(\add_98_3/n237 ), .ZN(
        \add_98_3/n251 ) );
  NOR2_X2 \add_98_3/U119  ( .A1(\add_98_3/n251 ), .A2(\add_98_3/n35 ), .ZN(
        \add_98_3/n248 ) );
  NOR2_X2 \add_98_3/U118  ( .A1(\add_98_3/n314 ), .A2(\add_98_3/n15 ), .ZN(
        \add_98_3/n320 ) );
  NOR3_X2 \add_98_3/U117  ( .A1(\add_98_3/n135 ), .A2(\add_98_3/n130 ), .A3(
        \add_98_3/n131 ), .ZN(\add_98_3/n128 ) );
  NOR2_X2 \add_98_3/U116  ( .A1(\add_98_3/n128 ), .A2(\add_98_3/n129 ), .ZN(
        \add_98_3/n124 ) );
  NOR2_X2 \add_98_3/U115  ( .A1(\add_98_3/n124 ), .A2(\add_98_3/n125 ), .ZN(
        \add_98_3/n121 ) );
  NOR2_X2 \add_98_3/U114  ( .A1(\add_98_3/n43 ), .A2(\add_98_3/n52 ), .ZN(
        \add_98_3/n380 ) );
  NOR2_X2 \add_98_3/U113  ( .A1(\add_98_3/n147 ), .A2(\add_98_3/n127 ), .ZN(
        \add_98_3/n193 ) );
  NAND3_X2 \add_98_3/U112  ( .A1(\add_98_3/n217 ), .A2(\add_98_3/n218 ), .A3(
        \add_98_3/n373 ), .ZN(\add_98_3/n212 ) );
  AND3_X2 \add_98_3/U111  ( .A1(\add_98_3/n171 ), .A2(\add_98_3/n159 ), .A3(
        \add_98_3/n172 ), .ZN(\add_98_3/n30 ) );
  NAND3_X2 \add_98_3/U110  ( .A1(\add_98_3/n150 ), .A2(\add_98_3/n151 ), .A3(
        \add_98_3/n30 ), .ZN(\add_98_3/n122 ) );
  NOR3_X2 \add_98_3/U109  ( .A1(\add_98_3/n194 ), .A2(\add_98_3/n147 ), .A3(
        \add_98_3/n195 ), .ZN(\add_98_3/n192 ) );
  NOR2_X2 \add_98_3/U108  ( .A1(\add_98_3/n314 ), .A2(\add_98_3/n15 ), .ZN(
        \add_98_3/n330 ) );
  NOR2_X2 \add_98_3/U107  ( .A1(\add_98_3/n46 ), .A2(\add_98_3/n43 ), .ZN(
        \add_98_3/n365 ) );
  AND3_X2 \add_98_3/U106  ( .A1(\add_98_3/n373 ), .A2(\add_98_3/n217 ), .A3(
        \add_98_3/n372 ), .ZN(\add_98_3/n29 ) );
  NAND3_X2 \add_98_3/U105  ( .A1(\add_98_3/n161 ), .A2(\add_98_3/n10 ), .A3(
        \add_98_3/n162 ), .ZN(\add_98_3/n160 ) );
  NAND3_X2 \add_98_3/U104  ( .A1(\add_98_3/n159 ), .A2(\add_98_3/n150 ), .A3(
        \add_98_3/n160 ), .ZN(\add_98_3/n157 ) );
  NOR2_X2 \add_98_3/U103  ( .A1(\add_98_3/n34 ), .A2(\add_98_3/n379 ), .ZN(
        \add_98_3/n378 ) );
  NAND3_X2 \add_98_3/U102  ( .A1(\add_98_3/n3 ), .A2(\add_98_3/n7 ), .A3(
        \add_98_3/n378 ), .ZN(\add_98_3/n49 ) );
  NOR2_X2 \add_98_3/U101  ( .A1(\add_98_3/n20 ), .A2(\add_98_3/n105 ), .ZN(
        \add_98_3/n94 ) );
  OR3_X4 \add_98_3/U100  ( .A1(\add_98_3/n307 ), .A2(\add_98_3/n308 ), .A3(
        \add_98_3/n38 ), .ZN(\add_98_3/n28 ) );
  OR2_X2 \add_98_3/U99  ( .A1(\add_98_3/n28 ), .A2(\add_98_3/n303 ), .ZN(
        \add_98_3/n301 ) );
  NOR2_X2 \add_98_3/U98  ( .A1(\add_98_3/n210 ), .A2(\add_98_3/n211 ), .ZN(
        \add_98_3/n209 ) );
  NAND3_X2 \add_98_3/U97  ( .A1(\add_98_3/n212 ), .A2(\add_98_3/n213 ), .A3(
        \add_98_3/n214 ), .ZN(\add_98_3/n208 ) );
  NAND3_X2 \add_98_3/U96  ( .A1(\add_98_3/n208 ), .A2(\add_98_3/n209 ), .A3(
        \add_98_3/n207 ), .ZN(\add_98_3/n206 ) );
  NAND3_X2 \add_98_3/U95  ( .A1(\add_98_3/n236 ), .A2(\add_98_3/n204 ), .A3(
        \add_98_3/n17 ), .ZN(\add_98_3/n232 ) );
  NAND3_X2 \add_98_3/U94  ( .A1(\add_98_3/n224 ), .A2(\add_98_3/n310 ), .A3(
        \add_98_3/n311 ), .ZN(\add_98_3/n133 ) );
  NOR2_X2 \add_98_3/U93  ( .A1(\add_98_3/n215 ), .A2(\add_98_3/n216 ), .ZN(
        \add_98_3/n288 ) );
  NAND3_X2 \add_98_3/U92  ( .A1(\add_98_3/n162 ), .A2(\add_98_3/n10 ), .A3(
        \add_98_3/n161 ), .ZN(\add_98_3/n170 ) );
  NOR2_X2 \add_98_3/U91  ( .A1(\add_98_3/n313 ), .A2(\add_98_3/n314 ), .ZN(
        \add_98_3/n312 ) );
  NAND3_X2 \add_98_3/U90  ( .A1(\add_98_3/n6 ), .A2(\add_98_3/n11 ), .A3(
        \add_98_3/n312 ), .ZN(\add_98_3/n215 ) );
  NOR3_X2 \add_98_3/U89  ( .A1(\add_98_3/n259 ), .A2(\add_98_3/n211 ), .A3(
        \add_98_3/n210 ), .ZN(\add_98_3/n256 ) );
  NOR2_X2 \add_98_3/U88  ( .A1(\add_98_3/n256 ), .A2(\add_98_3/n129 ), .ZN(
        \add_98_3/n254 ) );
  NOR2_X2 \add_98_3/U87  ( .A1(\add_98_3/n254 ), .A2(\add_98_3/n255 ), .ZN(
        \add_98_3/n237 ) );
  NOR3_X2 \add_98_3/U86  ( .A1(\add_98_3/n219 ), .A2(\add_98_3/n77 ), .A3(
        \add_98_3/n1 ), .ZN(\add_98_3/n297 ) );
  NOR2_X2 \add_98_3/U85  ( .A1(\add_98_3/n345 ), .A2(\add_98_3/n355 ), .ZN(
        \add_98_3/n354 ) );
  NAND3_X2 \add_98_3/U84  ( .A1(\add_98_3/n352 ), .A2(\add_98_3/n353 ), .A3(
        \add_98_3/n354 ), .ZN(\add_98_3/n216 ) );
  NOR3_X2 \add_98_3/U83  ( .A1(\add_98_3/n191 ), .A2(\add_98_3/n192 ), .A3(
        \add_98_3/n193 ), .ZN(\add_98_3/n190 ) );
  NOR2_X2 \add_98_3/U82  ( .A1(\add_98_3/n269 ), .A2(\add_98_3/n258 ), .ZN(
        \add_98_3/n264 ) );
  NOR2_X2 \add_98_3/U81  ( .A1(\add_98_3/n264 ), .A2(\add_98_3/n197 ), .ZN(
        \add_98_3/n263 ) );
  NOR2_X2 \add_98_3/U80  ( .A1(\add_98_3/n118 ), .A2(\add_98_3/n119 ), .ZN(
        \add_98_3/n115 ) );
  NOR3_X2 \add_98_3/U79  ( .A1(\add_98_3/n121 ), .A2(\add_98_3/n122 ), .A3(
        \add_98_3/n123 ), .ZN(\add_98_3/n111 ) );
  NOR2_X2 \add_98_3/U78  ( .A1(\add_98_3/n111 ), .A2(\add_98_3/n112 ), .ZN(
        \add_98_3/n106 ) );
  NOR2_X2 \add_98_3/U77  ( .A1(\add_98_3/n29 ), .A2(\add_98_3/n49 ), .ZN(
        \add_98_3/n53 ) );
  NOR2_X2 \add_98_3/U76  ( .A1(\add_98_3/n53 ), .A2(\add_98_3/n9 ), .ZN(
        \add_98_3/n50 ) );
  NOR2_X2 \add_98_3/U75  ( .A1(\add_98_3/n129 ), .A2(\add_98_3/n147 ), .ZN(
        \add_98_3/n205 ) );
  NOR2_X2 \add_98_3/U74  ( .A1(\add_98_3/n29 ), .A2(\add_98_3/n49 ), .ZN(
        \add_98_3/n356 ) );
  NOR2_X2 \add_98_3/U73  ( .A1(\add_98_3/n356 ), .A2(\add_98_3/n9 ), .ZN(
        \add_98_3/n351 ) );
  NOR2_X2 \add_98_3/U72  ( .A1(\add_98_3/n351 ), .A2(\add_98_3/n216 ), .ZN(
        \add_98_3/n338 ) );
  NOR2_X2 \add_98_3/U71  ( .A1(\add_98_3/n338 ), .A2(\add_98_3/n323 ), .ZN(
        \add_98_3/n335 ) );
  NOR2_X2 \add_98_3/U70  ( .A1(\add_98_3/n92 ), .A2(\add_98_3/n93 ), .ZN(
        \add_98_3/n89 ) );
  NOR2_X2 \add_98_3/U69  ( .A1(\add_98_3/n215 ), .A2(\add_98_3/n216 ), .ZN(
        \add_98_3/n213 ) );
  NOR2_X2 \add_98_3/U68  ( .A1(\add_98_3/n320 ), .A2(\add_98_3/n321 ), .ZN(
        \add_98_3/n319 ) );
  NOR3_X2 \add_98_3/U67  ( .A1(\add_98_3/n318 ), .A2(\add_98_3/n319 ), .A3(
        \add_98_3/n21 ), .ZN(\add_98_3/n317 ) );
  NOR2_X2 \add_98_3/U66  ( .A1(\add_98_3/n308 ), .A2(\add_98_3/n317 ), .ZN(
        \add_98_3/n316 ) );
  NOR2_X2 \add_98_3/U65  ( .A1(\add_98_3/n29 ), .A2(\add_98_3/n49 ), .ZN(
        \add_98_3/n322 ) );
  NAND3_X2 \add_98_3/U64  ( .A1(\add_98_3/n88 ), .A2(\add_98_3/n14 ), .A3(
        \add_98_3/n87 ), .ZN(\add_98_3/n144 ) );
  NOR3_X2 \add_98_3/U63  ( .A1(\add_98_3/n19 ), .A2(\add_98_3/n12 ), .A3(
        \add_98_3/n148 ), .ZN(\add_98_3/n143 ) );
  NOR2_X2 \add_98_3/U62  ( .A1(\add_98_3/n95 ), .A2(\add_98_3/n96 ), .ZN(
        \add_98_3/n84 ) );
  NOR2_X2 \add_98_3/U61  ( .A1(\add_98_3/n89 ), .A2(\add_98_3/n90 ), .ZN(
        \add_98_3/n85 ) );
  NOR4_X2 \add_98_3/U60  ( .A1(\add_98_3/n322 ), .A2(\add_98_3/n323 ), .A3(
        \add_98_3/n9 ), .A4(\add_98_3/n321 ), .ZN(\add_98_3/n318 ) );
  NOR2_X2 \add_98_3/U59  ( .A1(\add_98_3/n262 ), .A2(\add_98_3/n77 ), .ZN(
        \add_98_3/n299 ) );
  NOR2_X2 \add_98_3/U58  ( .A1(\add_98_3/n49 ), .A2(\add_98_3/n297 ), .ZN(
        \add_98_3/n296 ) );
  NOR2_X2 \add_98_3/U57  ( .A1(\add_98_3/n215 ), .A2(\add_98_3/n216 ), .ZN(
        \add_98_3/n294 ) );
  NAND3_X2 \add_98_3/U56  ( .A1(\add_98_3/n294 ), .A2(\add_98_3/n295 ), .A3(
        \add_98_3/n296 ), .ZN(\add_98_3/n134 ) );
  NAND3_X2 \add_98_3/U55  ( .A1(\add_98_3/n87 ), .A2(\add_98_3/n88 ), .A3(
        \add_98_3/n13 ), .ZN(\add_98_3/n86 ) );
  NOR2_X2 \add_98_3/U54  ( .A1(\add_98_3/n211 ), .A2(\add_98_3/n210 ), .ZN(
        \add_98_3/n286 ) );
  NAND3_X2 \add_98_3/U53  ( .A1(\add_98_3/n286 ), .A2(\add_98_3/n134 ), .A3(
        \add_98_3/n260 ), .ZN(\add_98_3/n88 ) );
  NAND3_X1 \add_98_3/U52  ( .A1(cv_q[84]), .A2(rnd_q[84]), .A3(\add_98_3/n243 ), .ZN(\add_98_3/n203 ) );
  OR2_X4 \add_98_3/U51  ( .A1(rnd_q[64]), .A2(cv_q[64]), .ZN(\add_98_3/n374 )
         );
  OR2_X1 \add_98_3/U50  ( .A1(cv_q[81]), .A2(rnd_q[81]), .ZN(\add_98_3/n33 )
         );
  NOR2_X1 \add_98_3/U49  ( .A1(cv_q[81]), .A2(rnd_q[81]), .ZN(\add_98_3/n278 )
         );
  OR2_X4 \add_98_3/U48  ( .A1(rnd_q[82]), .A2(cv_q[82]), .ZN(\add_98_3/n268 )
         );
  NAND2_X1 \add_98_3/U47  ( .A1(cv_q[80]), .A2(rnd_q[80]), .ZN(\add_98_3/n279 ) );
  NOR2_X1 \add_98_3/U46  ( .A1(cv_q[65]), .A2(rnd_q[65]), .ZN(\add_98_3/n137 )
         );
  NOR2_X1 \add_98_3/U45  ( .A1(cv_q[81]), .A2(rnd_q[81]), .ZN(\add_98_3/n275 )
         );
  NOR2_X1 \add_98_3/U44  ( .A1(cv_q[84]), .A2(rnd_q[84]), .ZN(\add_98_3/n252 )
         );
  OR2_X4 \add_98_3/U43  ( .A1(rnd_q[86]), .A2(cv_q[86]), .ZN(\add_98_3/n199 )
         );
  NOR2_X1 \add_98_3/U42  ( .A1(cv_q[84]), .A2(rnd_q[84]), .ZN(\add_98_3/n247 )
         );
  NOR2_X1 \add_98_3/U41  ( .A1(cv_q[85]), .A2(rnd_q[85]), .ZN(\add_98_3/n246 )
         );
  NOR2_X1 \add_98_3/U40  ( .A1(cv_q[85]), .A2(rnd_q[85]), .ZN(\add_98_3/n244 )
         );
  OR2_X4 \add_98_3/U39  ( .A1(rnd_q[83]), .A2(cv_q[83]), .ZN(\add_98_3/n196 )
         );
  NOR2_X1 \add_98_3/U38  ( .A1(cv_q[80]), .A2(rnd_q[80]), .ZN(\add_98_3/n276 )
         );
  OR2_X4 \add_98_3/U37  ( .A1(rnd_q[79]), .A2(cv_q[79]), .ZN(\add_98_3/n302 )
         );
  OR2_X4 \add_98_3/U36  ( .A1(rnd_q[75]), .A2(cv_q[75]), .ZN(\add_98_3/n310 )
         );
  NOR2_X1 \add_98_3/U35  ( .A1(cv_q[76]), .A2(rnd_q[76]), .ZN(\add_98_3/n314 )
         );
  NOR2_X1 \add_98_3/U34  ( .A1(rnd_q[68]), .A2(cv_q[68]), .ZN(\add_98_3/n34 )
         );
  NOR2_X1 \add_98_3/U33  ( .A1(cv_q[73]), .A2(rnd_q[73]), .ZN(\add_98_3/n43 )
         );
  NOR2_X1 \add_98_3/U32  ( .A1(cv_q[72]), .A2(rnd_q[72]), .ZN(\add_98_3/n46 )
         );
  NOR2_X1 \add_98_3/U31  ( .A1(cv_q[78]), .A2(rnd_q[78]), .ZN(\add_98_3/n305 )
         );
  NOR2_X1 \add_98_3/U30  ( .A1(cv_q[74]), .A2(rnd_q[74]), .ZN(\add_98_3/n345 )
         );
  NOR2_X1 \add_98_3/U29  ( .A1(cv_q[77]), .A2(rnd_q[77]), .ZN(\add_98_3/n306 )
         );
  AND2_X4 \add_98_3/U28  ( .A1(\add_98_3/n374 ), .A2(\add_98_3/n222 ), .ZN(N93) );
  AND2_X4 \add_98_3/U27  ( .A1(\add_98_3/n199 ), .A2(\add_98_3/n204 ), .ZN(
        \add_98_3/n26 ) );
  AND2_X4 \add_98_3/U26  ( .A1(\add_98_3/n151 ), .A2(\add_98_3/n101 ), .ZN(
        \add_98_3/n25 ) );
  AND2_X4 \add_98_3/U25  ( .A1(\add_98_3/n159 ), .A2(\add_98_3/n162 ), .ZN(
        \add_98_3/n24 ) );
  AND2_X4 \add_98_3/U24  ( .A1(\add_98_3/n127 ), .A2(\add_98_3/n196 ), .ZN(
        \add_98_3/n23 ) );
  OR2_X4 \add_98_3/U23  ( .A1(\add_98_3/n306 ), .A2(\add_98_3/n324 ), .ZN(
        \add_98_3/n22 ) );
  OR2_X4 \add_98_3/U22  ( .A1(\add_98_3/n305 ), .A2(\add_98_3/n306 ), .ZN(
        \add_98_3/n21 ) );
  AND2_X4 \add_98_3/U21  ( .A1(\add_98_3/n109 ), .A2(\add_98_3/n110 ), .ZN(
        \add_98_3/n20 ) );
  AND2_X4 \add_98_3/U20  ( .A1(\add_98_3/n153 ), .A2(\add_98_3/n151 ), .ZN(
        \add_98_3/n19 ) );
  AND3_X4 \add_98_3/U19  ( .A1(\add_98_3/n30 ), .A2(\add_98_3/n150 ), .A3(
        \add_98_3/n163 ), .ZN(\add_98_3/n18 ) );
  OR2_X4 \add_98_3/U18  ( .A1(\add_98_3/n237 ), .A2(\add_98_3/n231 ), .ZN(
        \add_98_3/n17 ) );
  OR2_X4 \add_98_3/U17  ( .A1(\add_98_3/n345 ), .A2(\add_98_3/n346 ), .ZN(
        \add_98_3/n16 ) );
  AND2_X4 \add_98_3/U16  ( .A1(\add_98_3/n216 ), .A2(\add_98_3/n334 ), .ZN(
        \add_98_3/n15 ) );
  AND2_X4 \add_98_3/U15  ( .A1(\add_98_3/n103 ), .A2(\add_98_3/n104 ), .ZN(
        \add_98_3/n14 ) );
  AND3_X4 \add_98_3/U14  ( .A1(\add_98_3/n103 ), .A2(\add_98_3/n94 ), .A3(
        \add_98_3/n104 ), .ZN(\add_98_3/n13 ) );
  AND2_X4 \add_98_3/U13  ( .A1(\add_98_3/n149 ), .A2(\add_98_3/n104 ), .ZN(
        \add_98_3/n12 ) );
  OR2_X4 \add_98_3/U12  ( .A1(cv_q[78]), .A2(rnd_q[78]), .ZN(\add_98_3/n11 )
         );
  OR2_X4 \add_98_3/U11  ( .A1(\add_98_3/n178 ), .A2(\add_98_3/n179 ), .ZN(
        \add_98_3/n10 ) );
  AND2_X4 \add_98_3/U10  ( .A1(\add_98_3/n366 ), .A2(\add_98_3/n3 ), .ZN(
        \add_98_3/n9 ) );
  OR2_X4 \add_98_3/U9  ( .A1(cv_q[67]), .A2(rnd_q[67]), .ZN(\add_98_3/n8 ) );
  OR2_X4 \add_98_3/U8  ( .A1(cv_q[70]), .A2(rnd_q[70]), .ZN(\add_98_3/n7 ) );
  OR2_X4 \add_98_3/U7  ( .A1(cv_q[77]), .A2(rnd_q[77]), .ZN(\add_98_3/n6 ) );
  OR3_X4 \add_98_3/U6  ( .A1(\add_98_3/n322 ), .A2(\add_98_3/n9 ), .A3(
        \add_98_3/n323 ), .ZN(\add_98_3/n5 ) );
  OR2_X4 \add_98_3/U5  ( .A1(cv_q[66]), .A2(rnd_q[66]), .ZN(\add_98_3/n4 ) );
  OR2_X4 \add_98_3/U4  ( .A1(cv_q[71]), .A2(rnd_q[71]), .ZN(\add_98_3/n3 ) );
  OR2_X4 \add_98_3/U3  ( .A1(cv_q[65]), .A2(rnd_q[65]), .ZN(\add_98_3/n2 ) );
  AND3_X4 \add_98_3/U2  ( .A1(\add_98_3/n4 ), .A2(\add_98_3/n8 ), .A3(
        \add_98_3/n2 ), .ZN(\add_98_3/n1 ) );
  INV_X4 \add_98_5/U424  ( .A(rnd_q[0]), .ZN(\add_98_5/n391 ) );
  INV_X4 \add_98_5/U423  ( .A(cv_q[0]), .ZN(\add_98_5/n392 ) );
  NAND2_X2 \add_98_5/U422  ( .A1(\add_98_5/n391 ), .A2(\add_98_5/n392 ), .ZN(
        \add_98_5/n381 ) );
  NAND2_X2 \add_98_5/U421  ( .A1(rnd_q[0]), .A2(cv_q[0]), .ZN(\add_98_5/n221 )
         );
  INV_X4 \add_98_5/U420  ( .A(\add_98_5/n352 ), .ZN(\add_98_5/n390 ) );
  NAND2_X2 \add_98_5/U419  ( .A1(rnd_q[10]), .A2(cv_q[10]), .ZN(
        \add_98_5/n351 ) );
  NAND2_X2 \add_98_5/U418  ( .A1(\add_98_5/n390 ), .A2(\add_98_5/n351 ), .ZN(
        \add_98_5/n368 ) );
  NAND2_X2 \add_98_5/U417  ( .A1(rnd_q[8]), .A2(cv_q[8]), .ZN(\add_98_5/n53 )
         );
  INV_X4 \add_98_5/U416  ( .A(rnd_q[4]), .ZN(\add_98_5/n387 ) );
  INV_X4 \add_98_5/U415  ( .A(cv_q[4]), .ZN(\add_98_5/n388 ) );
  INV_X4 \add_98_5/U414  ( .A(\add_98_5/n50 ), .ZN(\add_98_5/n378 ) );
  NAND2_X2 \add_98_5/U413  ( .A1(rnd_q[1]), .A2(cv_q[1]), .ZN(\add_98_5/n384 )
         );
  NAND2_X2 \add_98_5/U412  ( .A1(\add_98_5/n384 ), .A2(\add_98_5/n221 ), .ZN(
        \add_98_5/n383 ) );
  NAND2_X2 \add_98_5/U411  ( .A1(\add_98_5/n1 ), .A2(\add_98_5/n383 ), .ZN(
        \add_98_5/n380 ) );
  NAND2_X2 \add_98_5/U410  ( .A1(cv_q[2]), .A2(rnd_q[2]), .ZN(\add_98_5/n382 )
         );
  NAND2_X2 \add_98_5/U409  ( .A1(rnd_q[3]), .A2(cv_q[3]), .ZN(\add_98_5/n215 )
         );
  INV_X4 \add_98_5/U408  ( .A(\add_98_5/n33 ), .ZN(\add_98_5/n379 ) );
  NAND2_X2 \add_98_5/U407  ( .A1(rnd_q[7]), .A2(cv_q[7]), .ZN(\add_98_5/n57 )
         );
  NAND2_X2 \add_98_5/U406  ( .A1(rnd_q[6]), .A2(cv_q[6]), .ZN(\add_98_5/n377 )
         );
  NAND2_X2 \add_98_5/U405  ( .A1(rnd_q[4]), .A2(cv_q[4]), .ZN(\add_98_5/n67 )
         );
  NAND2_X2 \add_98_5/U404  ( .A1(rnd_q[5]), .A2(cv_q[5]), .ZN(\add_98_5/n64 )
         );
  NAND2_X2 \add_98_5/U403  ( .A1(\add_98_5/n67 ), .A2(\add_98_5/n64 ), .ZN(
        \add_98_5/n376 ) );
  NAND2_X2 \add_98_5/U402  ( .A1(\add_98_5/n375 ), .A2(\add_98_5/n376 ), .ZN(
        \add_98_5/n374 ) );
  NAND2_X2 \add_98_5/U401  ( .A1(\add_98_5/n38 ), .A2(\add_98_5/n374 ), .ZN(
        \add_98_5/n373 ) );
  NAND2_X2 \add_98_5/U400  ( .A1(\add_98_5/n19 ), .A2(\add_98_5/n372 ), .ZN(
        \add_98_5/n371 ) );
  XNOR2_X2 \add_98_5/U399  ( .A(\add_98_5/n368 ), .B(\add_98_5/n367 ), .ZN(
        N167) );
  NAND2_X2 \add_98_5/U398  ( .A1(\add_98_5/n367 ), .A2(\add_98_5/n390 ), .ZN(
        \add_98_5/n366 ) );
  NAND2_X2 \add_98_5/U397  ( .A1(\add_98_5/n366 ), .A2(\add_98_5/n351 ), .ZN(
        \add_98_5/n364 ) );
  NAND2_X2 \add_98_5/U396  ( .A1(rnd_q[11]), .A2(cv_q[11]), .ZN(
        \add_98_5/n350 ) );
  NAND2_X2 \add_98_5/U395  ( .A1(\add_98_5/n350 ), .A2(\add_98_5/n315 ), .ZN(
        \add_98_5/n365 ) );
  XNOR2_X2 \add_98_5/U394  ( .A(\add_98_5/n364 ), .B(\add_98_5/n365 ), .ZN(
        N168) );
  INV_X4 \add_98_5/U393  ( .A(\add_98_5/n44 ), .ZN(\add_98_5/n359 ) );
  INV_X4 \add_98_5/U392  ( .A(\add_98_5/n47 ), .ZN(\add_98_5/n360 ) );
  INV_X4 \add_98_5/U391  ( .A(\add_98_5/n315 ), .ZN(\add_98_5/n362 ) );
  NAND2_X2 \add_98_5/U390  ( .A1(\add_98_5/n354 ), .A2(\add_98_5/n355 ), .ZN(
        \add_98_5/n346 ) );
  NAND2_X2 \add_98_5/U389  ( .A1(cv_q[9]), .A2(rnd_q[9]), .ZN(\add_98_5/n353 )
         );
  INV_X4 \add_98_5/U388  ( .A(\add_98_5/n351 ), .ZN(\add_98_5/n348 ) );
  INV_X4 \add_98_5/U387  ( .A(\add_98_5/n350 ), .ZN(\add_98_5/n349 ) );
  NAND2_X2 \add_98_5/U386  ( .A1(\add_98_5/n316 ), .A2(\add_98_5/n315 ), .ZN(
        \add_98_5/n341 ) );
  INV_X4 \add_98_5/U385  ( .A(\add_98_5/n341 ), .ZN(\add_98_5/n328 ) );
  NAND2_X2 \add_98_5/U384  ( .A1(rnd_q[12]), .A2(cv_q[12]), .ZN(
        \add_98_5/n329 ) );
  INV_X4 \add_98_5/U383  ( .A(\add_98_5/n329 ), .ZN(\add_98_5/n344 ) );
  XNOR2_X2 \add_98_5/U382  ( .A(\add_98_5/n342 ), .B(\add_98_5/n343 ), .ZN(
        N169) );
  NAND2_X2 \add_98_5/U381  ( .A1(\add_98_5/n337 ), .A2(\add_98_5/n6 ), .ZN(
        \add_98_5/n340 ) );
  NAND2_X2 \add_98_5/U380  ( .A1(\add_98_5/n340 ), .A2(\add_98_5/n329 ), .ZN(
        \add_98_5/n338 ) );
  NAND2_X2 \add_98_5/U379  ( .A1(rnd_q[13]), .A2(cv_q[13]), .ZN(
        \add_98_5/n330 ) );
  NAND2_X2 \add_98_5/U378  ( .A1(\add_98_5/n330 ), .A2(\add_98_5/n4 ), .ZN(
        \add_98_5/n339 ) );
  XNOR2_X2 \add_98_5/U377  ( .A(\add_98_5/n338 ), .B(\add_98_5/n339 ), .ZN(
        N170) );
  NAND2_X2 \add_98_5/U376  ( .A1(rnd_q[14]), .A2(cv_q[14]), .ZN(
        \add_98_5/n331 ) );
  NAND2_X2 \add_98_5/U375  ( .A1(\add_98_5/n9 ), .A2(\add_98_5/n331 ), .ZN(
        \add_98_5/n335 ) );
  XNOR2_X2 \add_98_5/U374  ( .A(\add_98_5/n334 ), .B(\add_98_5/n335 ), .ZN(
        N171) );
  INV_X4 \add_98_5/U373  ( .A(rnd_q[15]), .ZN(\add_98_5/n332 ) );
  INV_X4 \add_98_5/U372  ( .A(cv_q[15]), .ZN(\add_98_5/n333 ) );
  NAND2_X2 \add_98_5/U371  ( .A1(\add_98_5/n332 ), .A2(\add_98_5/n333 ), .ZN(
        \add_98_5/n306 ) );
  INV_X4 \add_98_5/U370  ( .A(\add_98_5/n306 ), .ZN(\add_98_5/n318 ) );
  INV_X4 \add_98_5/U369  ( .A(\add_98_5/n331 ), .ZN(\add_98_5/n312 ) );
  NAND2_X2 \add_98_5/U368  ( .A1(\add_98_5/n329 ), .A2(\add_98_5/n330 ), .ZN(
        \add_98_5/n326 ) );
  XNOR2_X2 \add_98_5/U367  ( .A(\add_98_5/n320 ), .B(\add_98_5/n321 ), .ZN(
        N172) );
  NAND2_X2 \add_98_5/U366  ( .A1(rnd_q[16]), .A2(cv_q[16]), .ZN(
        \add_98_5/n287 ) );
  NAND2_X2 \add_98_5/U365  ( .A1(\add_98_5/n287 ), .A2(\add_98_5/n289 ), .ZN(
        \add_98_5/n290 ) );
  INV_X4 \add_98_5/U364  ( .A(\add_98_5/n213 ), .ZN(\add_98_5/n314 ) );
  INV_X4 \add_98_5/U363  ( .A(\add_98_5/n132 ), .ZN(\add_98_5/n210 ) );
  NAND2_X2 \add_98_5/U362  ( .A1(cv_q[13]), .A2(rnd_q[13]), .ZN(
        \add_98_5/n313 ) );
  NAND2_X2 \add_98_5/U361  ( .A1(rnd_q[12]), .A2(cv_q[12]), .ZN(
        \add_98_5/n308 ) );
  NAND2_X2 \add_98_5/U360  ( .A1(\add_98_5/n305 ), .A2(\add_98_5/n306 ), .ZN(
        \add_98_5/n131 ) );
  INV_X4 \add_98_5/U359  ( .A(\add_98_5/n131 ), .ZN(\add_98_5/n209 ) );
  NAND2_X2 \add_98_5/U358  ( .A1(rnd_q[1]), .A2(cv_q[1]), .ZN(\add_98_5/n137 )
         );
  INV_X4 \add_98_5/U357  ( .A(\add_98_5/n137 ), .ZN(\add_98_5/n262 ) );
  INV_X4 \add_98_5/U356  ( .A(\add_98_5/n215 ), .ZN(\add_98_5/n78 ) );
  NAND2_X2 \add_98_5/U355  ( .A1(\add_98_5/n303 ), .A2(\add_98_5/n304 ), .ZN(
        \add_98_5/n300 ) );
  NAND2_X2 \add_98_5/U354  ( .A1(rnd_q[5]), .A2(cv_q[5]), .ZN(\add_98_5/n296 )
         );
  NAND2_X2 \add_98_5/U353  ( .A1(\add_98_5/n67 ), .A2(\add_98_5/n296 ), .ZN(
        \add_98_5/n295 ) );
  NAND2_X2 \add_98_5/U352  ( .A1(\add_98_5/n225 ), .A2(\add_98_5/n295 ), .ZN(
        \add_98_5/n294 ) );
  NAND2_X2 \add_98_5/U351  ( .A1(\add_98_5/n38 ), .A2(\add_98_5/n294 ), .ZN(
        \add_98_5/n292 ) );
  NAND3_X2 \add_98_5/U350  ( .A1(\add_98_5/n292 ), .A2(\add_98_5/n3 ), .A3(
        \add_98_5/n293 ), .ZN(\add_98_5/n260 ) );
  INV_X4 \add_98_5/U349  ( .A(\add_98_5/n260 ), .ZN(\add_98_5/n134 ) );
  XNOR2_X2 \add_98_5/U348  ( .A(\add_98_5/n290 ), .B(\add_98_5/n89 ), .ZN(N173) );
  INV_X4 \add_98_5/U347  ( .A(\add_98_5/n281 ), .ZN(\add_98_5/n289 ) );
  NAND2_X2 \add_98_5/U346  ( .A1(\add_98_5/n89 ), .A2(\add_98_5/n289 ), .ZN(
        \add_98_5/n288 ) );
  NAND2_X2 \add_98_5/U345  ( .A1(\add_98_5/n287 ), .A2(\add_98_5/n288 ), .ZN(
        \add_98_5/n285 ) );
  NAND2_X2 \add_98_5/U344  ( .A1(rnd_q[17]), .A2(cv_q[17]), .ZN(
        \add_98_5/n282 ) );
  NAND2_X2 \add_98_5/U343  ( .A1(\add_98_5/n39 ), .A2(\add_98_5/n282 ), .ZN(
        \add_98_5/n286 ) );
  XNOR2_X2 \add_98_5/U342  ( .A(\add_98_5/n285 ), .B(\add_98_5/n286 ), .ZN(
        N174) );
  NAND2_X2 \add_98_5/U341  ( .A1(cv_q[16]), .A2(rnd_q[16]), .ZN(
        \add_98_5/n284 ) );
  NAND2_X2 \add_98_5/U340  ( .A1(\add_98_5/n31 ), .A2(\add_98_5/n282 ), .ZN(
        \add_98_5/n270 ) );
  INV_X4 \add_98_5/U339  ( .A(\add_98_5/n270 ), .ZN(\add_98_5/n278 ) );
  NAND2_X2 \add_98_5/U338  ( .A1(\add_98_5/n273 ), .A2(\add_98_5/n89 ), .ZN(
        \add_98_5/n279 ) );
  NAND2_X2 \add_98_5/U337  ( .A1(\add_98_5/n278 ), .A2(\add_98_5/n279 ), .ZN(
        \add_98_5/n274 ) );
  NAND2_X2 \add_98_5/U336  ( .A1(rnd_q[18]), .A2(cv_q[18]), .ZN(
        \add_98_5/n269 ) );
  INV_X4 \add_98_5/U335  ( .A(rnd_q[18]), .ZN(\add_98_5/n276 ) );
  INV_X4 \add_98_5/U334  ( .A(cv_q[18]), .ZN(\add_98_5/n277 ) );
  NAND2_X2 \add_98_5/U333  ( .A1(\add_98_5/n276 ), .A2(\add_98_5/n277 ), .ZN(
        \add_98_5/n271 ) );
  NAND2_X2 \add_98_5/U332  ( .A1(\add_98_5/n269 ), .A2(\add_98_5/n271 ), .ZN(
        \add_98_5/n275 ) );
  XNOR2_X2 \add_98_5/U331  ( .A(\add_98_5/n274 ), .B(\add_98_5/n275 ), .ZN(
        N175) );
  INV_X4 \add_98_5/U330  ( .A(\add_98_5/n89 ), .ZN(\add_98_5/n272 ) );
  NAND2_X2 \add_98_5/U329  ( .A1(\add_98_5/n273 ), .A2(\add_98_5/n271 ), .ZN(
        \add_98_5/n258 ) );
  NAND2_X2 \add_98_5/U328  ( .A1(\add_98_5/n270 ), .A2(\add_98_5/n271 ), .ZN(
        \add_98_5/n268 ) );
  NAND2_X2 \add_98_5/U327  ( .A1(\add_98_5/n268 ), .A2(\add_98_5/n269 ), .ZN(
        \add_98_5/n196 ) );
  NAND2_X2 \add_98_5/U326  ( .A1(rnd_q[19]), .A2(cv_q[19]), .ZN(
        \add_98_5/n126 ) );
  INV_X4 \add_98_5/U325  ( .A(rnd_q[19]), .ZN(\add_98_5/n265 ) );
  INV_X4 \add_98_5/U324  ( .A(cv_q[19]), .ZN(\add_98_5/n266 ) );
  NAND2_X2 \add_98_5/U323  ( .A1(\add_98_5/n265 ), .A2(\add_98_5/n266 ), .ZN(
        \add_98_5/n195 ) );
  XNOR2_X2 \add_98_5/U322  ( .A(\add_98_5/n264 ), .B(\add_98_5/n25 ), .ZN(N176) );
  INV_X4 \add_98_5/U321  ( .A(\add_98_5/n221 ), .ZN(\add_98_5/n263 ) );
  XNOR2_X2 \add_98_5/U320  ( .A(\add_98_5/n221 ), .B(\add_98_5/n261 ), .ZN(
        N158) );
  INV_X4 \add_98_5/U319  ( .A(\add_98_5/n258 ), .ZN(\add_98_5/n257 ) );
  NAND2_X2 \add_98_5/U318  ( .A1(\add_98_5/n257 ), .A2(\add_98_5/n195 ), .ZN(
        \add_98_5/n128 ) );
  NAND2_X2 \add_98_5/U317  ( .A1(\add_98_5/n196 ), .A2(\add_98_5/n195 ), .ZN(
        \add_98_5/n125 ) );
  NAND2_X2 \add_98_5/U316  ( .A1(\add_98_5/n125 ), .A2(\add_98_5/n126 ), .ZN(
        \add_98_5/n255 ) );
  XNOR2_X2 \add_98_5/U315  ( .A(\add_98_5/n235 ), .B(\add_98_5/n253 ), .ZN(
        N177) );
  NAND2_X2 \add_98_5/U314  ( .A1(rnd_q[21]), .A2(cv_q[21]), .ZN(
        \add_98_5/n201 ) );
  INV_X4 \add_98_5/U313  ( .A(\add_98_5/n201 ), .ZN(\add_98_5/n250 ) );
  XNOR2_X2 \add_98_5/U312  ( .A(\add_98_5/n248 ), .B(\add_98_5/n249 ), .ZN(
        N178) );
  INV_X4 \add_98_5/U311  ( .A(\add_98_5/n236 ), .ZN(\add_98_5/n245 ) );
  INV_X4 \add_98_5/U310  ( .A(\add_98_5/n244 ), .ZN(\add_98_5/n243 ) );
  NAND2_X2 \add_98_5/U309  ( .A1(\add_98_5/n202 ), .A2(\add_98_5/n201 ), .ZN(
        \add_98_5/n242 ) );
  INV_X4 \add_98_5/U308  ( .A(rnd_q[22]), .ZN(\add_98_5/n239 ) );
  INV_X4 \add_98_5/U307  ( .A(cv_q[22]), .ZN(\add_98_5/n240 ) );
  NAND2_X2 \add_98_5/U306  ( .A1(\add_98_5/n239 ), .A2(\add_98_5/n240 ), .ZN(
        \add_98_5/n198 ) );
  NAND2_X2 \add_98_5/U305  ( .A1(rnd_q[22]), .A2(cv_q[22]), .ZN(
        \add_98_5/n203 ) );
  XNOR2_X2 \add_98_5/U304  ( .A(\add_98_5/n238 ), .B(\add_98_5/n28 ), .ZN(N179) );
  NAND2_X2 \add_98_5/U303  ( .A1(\add_98_5/n202 ), .A2(\add_98_5/n201 ), .ZN(
        \add_98_5/n237 ) );
  NAND2_X2 \add_98_5/U302  ( .A1(\add_98_5/n237 ), .A2(\add_98_5/n198 ), .ZN(
        \add_98_5/n234 ) );
  NAND2_X2 \add_98_5/U301  ( .A1(\add_98_5/n236 ), .A2(\add_98_5/n198 ), .ZN(
        \add_98_5/n229 ) );
  INV_X4 \add_98_5/U300  ( .A(rnd_q[23]), .ZN(\add_98_5/n232 ) );
  INV_X4 \add_98_5/U299  ( .A(cv_q[23]), .ZN(\add_98_5/n233 ) );
  NAND2_X2 \add_98_5/U298  ( .A1(\add_98_5/n232 ), .A2(\add_98_5/n233 ), .ZN(
        \add_98_5/n199 ) );
  NAND2_X2 \add_98_5/U297  ( .A1(rnd_q[23]), .A2(cv_q[23]), .ZN(
        \add_98_5/n151 ) );
  NAND2_X2 \add_98_5/U296  ( .A1(\add_98_5/n199 ), .A2(\add_98_5/n151 ), .ZN(
        \add_98_5/n231 ) );
  XNOR2_X2 \add_98_5/U295  ( .A(\add_98_5/n230 ), .B(\add_98_5/n231 ), .ZN(
        N180) );
  INV_X4 \add_98_5/U294  ( .A(\add_98_5/n229 ), .ZN(\add_98_5/n228 ) );
  NAND2_X2 \add_98_5/U293  ( .A1(\add_98_5/n228 ), .A2(\add_98_5/n199 ), .ZN(
        \add_98_5/n146 ) );
  NAND2_X2 \add_98_5/U292  ( .A1(rnd_q[5]), .A2(cv_q[5]), .ZN(\add_98_5/n227 )
         );
  NAND2_X2 \add_98_5/U291  ( .A1(\add_98_5/n67 ), .A2(\add_98_5/n227 ), .ZN(
        \add_98_5/n226 ) );
  NAND2_X2 \add_98_5/U290  ( .A1(\add_98_5/n225 ), .A2(\add_98_5/n226 ), .ZN(
        \add_98_5/n224 ) );
  NAND2_X2 \add_98_5/U289  ( .A1(\add_98_5/n38 ), .A2(\add_98_5/n224 ), .ZN(
        \add_98_5/n222 ) );
  INV_X4 \add_98_5/U288  ( .A(\add_98_5/n214 ), .ZN(\add_98_5/n223 ) );
  NAND4_X2 \add_98_5/U287  ( .A1(\add_98_5/n222 ), .A2(\add_98_5/n3 ), .A3(
        \add_98_5/n314 ), .A4(\add_98_5/n223 ), .ZN(\add_98_5/n206 ) );
  NAND2_X2 \add_98_5/U286  ( .A1(rnd_q[1]), .A2(cv_q[1]), .ZN(\add_98_5/n220 )
         );
  NAND2_X2 \add_98_5/U285  ( .A1(\add_98_5/n220 ), .A2(\add_98_5/n221 ), .ZN(
        \add_98_5/n219 ) );
  NAND2_X2 \add_98_5/U284  ( .A1(\add_98_5/n1 ), .A2(\add_98_5/n219 ), .ZN(
        \add_98_5/n216 ) );
  INV_X4 \add_98_5/U283  ( .A(\add_98_5/n218 ), .ZN(\add_98_5/n217 ) );
  NAND2_X2 \add_98_5/U282  ( .A1(\add_98_5/n204 ), .A2(\add_98_5/n205 ), .ZN(
        \add_98_5/n188 ) );
  INV_X4 \add_98_5/U281  ( .A(\add_98_5/n145 ), .ZN(\add_98_5/n197 ) );
  NAND2_X2 \add_98_5/U280  ( .A1(\add_98_5/n197 ), .A2(\add_98_5/n151 ), .ZN(
        \add_98_5/n190 ) );
  INV_X4 \add_98_5/U279  ( .A(\add_98_5/n196 ), .ZN(\add_98_5/n193 ) );
  INV_X4 \add_98_5/U278  ( .A(\add_98_5/n195 ), .ZN(\add_98_5/n194 ) );
  NAND2_X2 \add_98_5/U277  ( .A1(\add_98_5/n188 ), .A2(\add_98_5/n189 ), .ZN(
        \add_98_5/n162 ) );
  NAND2_X2 \add_98_5/U276  ( .A1(rnd_q[24]), .A2(cv_q[24]), .ZN(
        \add_98_5/n186 ) );
  NAND2_X2 \add_98_5/U275  ( .A1(\add_98_5/n186 ), .A2(\add_98_5/n171 ), .ZN(
        \add_98_5/n187 ) );
  XNOR2_X2 \add_98_5/U274  ( .A(\add_98_5/n162 ), .B(\add_98_5/n187 ), .ZN(
        N181) );
  INV_X4 \add_98_5/U273  ( .A(\add_98_5/n180 ), .ZN(\add_98_5/n171 ) );
  NAND2_X2 \add_98_5/U272  ( .A1(\add_98_5/n171 ), .A2(\add_98_5/n162 ), .ZN(
        \add_98_5/n185 ) );
  NAND2_X2 \add_98_5/U271  ( .A1(\add_98_5/n185 ), .A2(\add_98_5/n186 ), .ZN(
        \add_98_5/n181 ) );
  NAND2_X2 \add_98_5/U270  ( .A1(rnd_q[25]), .A2(cv_q[25]), .ZN(
        \add_98_5/n160 ) );
  INV_X4 \add_98_5/U269  ( .A(rnd_q[25]), .ZN(\add_98_5/n183 ) );
  INV_X4 \add_98_5/U268  ( .A(cv_q[25]), .ZN(\add_98_5/n184 ) );
  NAND2_X2 \add_98_5/U267  ( .A1(\add_98_5/n183 ), .A2(\add_98_5/n184 ), .ZN(
        \add_98_5/n170 ) );
  NAND2_X2 \add_98_5/U266  ( .A1(\add_98_5/n160 ), .A2(\add_98_5/n170 ), .ZN(
        \add_98_5/n182 ) );
  XNOR2_X2 \add_98_5/U265  ( .A(\add_98_5/n181 ), .B(\add_98_5/n182 ), .ZN(
        N182) );
  INV_X4 \add_98_5/U264  ( .A(\add_98_5/n162 ), .ZN(\add_98_5/n179 ) );
  INV_X4 \add_98_5/U263  ( .A(\add_98_5/n170 ), .ZN(\add_98_5/n177 ) );
  NAND2_X2 \add_98_5/U262  ( .A1(cv_q[24]), .A2(rnd_q[24]), .ZN(
        \add_98_5/n178 ) );
  NAND2_X2 \add_98_5/U261  ( .A1(\add_98_5/n8 ), .A2(\add_98_5/n160 ), .ZN(
        \add_98_5/n176 ) );
  INV_X4 \add_98_5/U260  ( .A(rnd_q[26]), .ZN(\add_98_5/n173 ) );
  INV_X4 \add_98_5/U259  ( .A(cv_q[26]), .ZN(\add_98_5/n174 ) );
  NAND2_X2 \add_98_5/U258  ( .A1(\add_98_5/n173 ), .A2(\add_98_5/n174 ), .ZN(
        \add_98_5/n158 ) );
  NAND2_X2 \add_98_5/U257  ( .A1(rnd_q[26]), .A2(cv_q[26]), .ZN(
        \add_98_5/n161 ) );
  XNOR2_X2 \add_98_5/U256  ( .A(\add_98_5/n172 ), .B(\add_98_5/n27 ), .ZN(N183) );
  NAND2_X2 \add_98_5/U255  ( .A1(\add_98_5/n34 ), .A2(\add_98_5/n162 ), .ZN(
        \add_98_5/n167 ) );
  NAND2_X2 \add_98_5/U254  ( .A1(\add_98_5/n169 ), .A2(\add_98_5/n158 ), .ZN(
        \add_98_5/n168 ) );
  NAND2_X2 \add_98_5/U253  ( .A1(\add_98_5/n167 ), .A2(\add_98_5/n168 ), .ZN(
        \add_98_5/n163 ) );
  INV_X4 \add_98_5/U252  ( .A(rnd_q[27]), .ZN(\add_98_5/n165 ) );
  INV_X4 \add_98_5/U251  ( .A(cv_q[27]), .ZN(\add_98_5/n166 ) );
  NAND2_X2 \add_98_5/U250  ( .A1(\add_98_5/n165 ), .A2(\add_98_5/n166 ), .ZN(
        \add_98_5/n149 ) );
  NAND2_X2 \add_98_5/U249  ( .A1(rnd_q[27]), .A2(cv_q[27]), .ZN(
        \add_98_5/n157 ) );
  NAND2_X2 \add_98_5/U248  ( .A1(\add_98_5/n149 ), .A2(\add_98_5/n157 ), .ZN(
        \add_98_5/n164 ) );
  XNOR2_X2 \add_98_5/U247  ( .A(\add_98_5/n163 ), .B(\add_98_5/n164 ), .ZN(
        N184) );
  NAND2_X2 \add_98_5/U246  ( .A1(\add_98_5/n156 ), .A2(\add_98_5/n157 ), .ZN(
        \add_98_5/n152 ) );
  INV_X4 \add_98_5/U245  ( .A(rnd_q[28]), .ZN(\add_98_5/n154 ) );
  INV_X4 \add_98_5/U244  ( .A(cv_q[28]), .ZN(\add_98_5/n155 ) );
  NAND2_X2 \add_98_5/U243  ( .A1(\add_98_5/n154 ), .A2(\add_98_5/n155 ), .ZN(
        \add_98_5/n150 ) );
  NAND2_X2 \add_98_5/U242  ( .A1(rnd_q[28]), .A2(cv_q[28]), .ZN(
        \add_98_5/n102 ) );
  XNOR2_X2 \add_98_5/U241  ( .A(\add_98_5/n153 ), .B(\add_98_5/n29 ), .ZN(N185) );
  INV_X4 \add_98_5/U240  ( .A(\add_98_5/n151 ), .ZN(\add_98_5/n148 ) );
  INV_X4 \add_98_5/U239  ( .A(\add_98_5/n121 ), .ZN(\add_98_5/n105 ) );
  INV_X4 \add_98_5/U238  ( .A(\add_98_5/n102 ), .ZN(\add_98_5/n147 ) );
  INV_X4 \add_98_5/U237  ( .A(\add_98_5/n146 ), .ZN(\add_98_5/n104 ) );
  INV_X4 \add_98_5/U236  ( .A(\add_98_5/n128 ), .ZN(\add_98_5/n88 ) );
  NAND2_X2 \add_98_5/U235  ( .A1(\add_98_5/n125 ), .A2(\add_98_5/n126 ), .ZN(
        \add_98_5/n103 ) );
  NAND2_X2 \add_98_5/U234  ( .A1(\add_98_5/n103 ), .A2(\add_98_5/n13 ), .ZN(
        \add_98_5/n144 ) );
  NAND2_X2 \add_98_5/U233  ( .A1(\add_98_5/n145 ), .A2(\add_98_5/n105 ), .ZN(
        \add_98_5/n94 ) );
  NAND4_X2 \add_98_5/U232  ( .A1(\add_98_5/n142 ), .A2(\add_98_5/n143 ), .A3(
        \add_98_5/n144 ), .A4(\add_98_5/n94 ), .ZN(\add_98_5/n138 ) );
  NAND2_X2 \add_98_5/U231  ( .A1(rnd_q[29]), .A2(cv_q[29]), .ZN(\add_98_5/n92 ) );
  INV_X4 \add_98_5/U230  ( .A(rnd_q[29]), .ZN(\add_98_5/n140 ) );
  INV_X4 \add_98_5/U229  ( .A(cv_q[29]), .ZN(\add_98_5/n141 ) );
  NAND2_X2 \add_98_5/U228  ( .A1(\add_98_5/n140 ), .A2(\add_98_5/n141 ), .ZN(
        \add_98_5/n118 ) );
  NAND2_X2 \add_98_5/U227  ( .A1(\add_98_5/n92 ), .A2(\add_98_5/n118 ), .ZN(
        \add_98_5/n139 ) );
  XNOR2_X2 \add_98_5/U226  ( .A(\add_98_5/n138 ), .B(\add_98_5/n139 ), .ZN(
        N186) );
  XNOR2_X2 \add_98_5/U225  ( .A(\add_98_5/n81 ), .B(\add_98_5/n135 ), .ZN(N159) );
  INV_X4 \add_98_5/U224  ( .A(\add_98_5/n133 ), .ZN(\add_98_5/n129 ) );
  NAND2_X2 \add_98_5/U223  ( .A1(\add_98_5/n131 ), .A2(\add_98_5/n132 ), .ZN(
        \add_98_5/n130 ) );
  NAND2_X2 \add_98_5/U222  ( .A1(\add_98_5/n125 ), .A2(\add_98_5/n126 ), .ZN(
        \add_98_5/n124 ) );
  NAND2_X2 \add_98_5/U221  ( .A1(\add_98_5/n104 ), .A2(\add_98_5/n118 ), .ZN(
        \add_98_5/n122 ) );
  NAND2_X2 \add_98_5/U220  ( .A1(\add_98_5/n21 ), .A2(\add_98_5/n118 ), .ZN(
        \add_98_5/n114 ) );
  INV_X4 \add_98_5/U219  ( .A(\add_98_5/n94 ), .ZN(\add_98_5/n119 ) );
  NAND2_X2 \add_98_5/U218  ( .A1(\add_98_5/n119 ), .A2(\add_98_5/n118 ), .ZN(
        \add_98_5/n115 ) );
  INV_X4 \add_98_5/U217  ( .A(\add_98_5/n118 ), .ZN(\add_98_5/n106 ) );
  NAND2_X2 \add_98_5/U216  ( .A1(\add_98_5/n11 ), .A2(\add_98_5/n118 ), .ZN(
        \add_98_5/n117 ) );
  NAND4_X2 \add_98_5/U215  ( .A1(\add_98_5/n114 ), .A2(\add_98_5/n115 ), .A3(
        \add_98_5/n116 ), .A4(\add_98_5/n117 ), .ZN(\add_98_5/n113 ) );
  INV_X4 \add_98_5/U214  ( .A(rnd_q[30]), .ZN(\add_98_5/n110 ) );
  INV_X4 \add_98_5/U213  ( .A(cv_q[30]), .ZN(\add_98_5/n111 ) );
  NAND2_X2 \add_98_5/U212  ( .A1(rnd_q[30]), .A2(cv_q[30]), .ZN(
        \add_98_5/n101 ) );
  INV_X4 \add_98_5/U211  ( .A(\add_98_5/n101 ), .ZN(\add_98_5/n109 ) );
  XNOR2_X2 \add_98_5/U210  ( .A(\add_98_5/n107 ), .B(\add_98_5/n108 ), .ZN(
        N187) );
  NAND2_X2 \add_98_5/U209  ( .A1(\add_98_5/n12 ), .A2(\add_98_5/n103 ), .ZN(
        \add_98_5/n84 ) );
  NAND2_X2 \add_98_5/U208  ( .A1(\add_98_5/n95 ), .A2(\add_98_5/n147 ), .ZN(
        \add_98_5/n100 ) );
  NAND2_X2 \add_98_5/U207  ( .A1(\add_98_5/n100 ), .A2(\add_98_5/n101 ), .ZN(
        \add_98_5/n96 ) );
  NAND2_X2 \add_98_5/U206  ( .A1(\add_98_5/n21 ), .A2(\add_98_5/n95 ), .ZN(
        \add_98_5/n98 ) );
  NAND2_X2 \add_98_5/U205  ( .A1(\add_98_5/n11 ), .A2(\add_98_5/n95 ), .ZN(
        \add_98_5/n99 ) );
  NAND2_X2 \add_98_5/U204  ( .A1(\add_98_5/n98 ), .A2(\add_98_5/n99 ), .ZN(
        \add_98_5/n97 ) );
  INV_X4 \add_98_5/U203  ( .A(\add_98_5/n95 ), .ZN(\add_98_5/n93 ) );
  NAND4_X2 \add_98_5/U202  ( .A1(\add_98_5/n84 ), .A2(\add_98_5/n85 ), .A3(
        \add_98_5/n86 ), .A4(\add_98_5/n87 ), .ZN(\add_98_5/n82 ) );
  XNOR2_X2 \add_98_5/U201  ( .A(rnd_q[31]), .B(cv_q[31]), .ZN(\add_98_5/n83 )
         );
  XNOR2_X2 \add_98_5/U200  ( .A(\add_98_5/n82 ), .B(\add_98_5/n83 ), .ZN(N188)
         );
  XNOR2_X2 \add_98_5/U199  ( .A(\add_98_5/n75 ), .B(\add_98_5/n76 ), .ZN(N160)
         );
  INV_X4 \add_98_5/U198  ( .A(\add_98_5/n67 ), .ZN(\add_98_5/n73 ) );
  XNOR2_X2 \add_98_5/U197  ( .A(\add_98_5/n33 ), .B(\add_98_5/n74 ), .ZN(N161)
         );
  INV_X4 \add_98_5/U196  ( .A(\add_98_5/n64 ), .ZN(\add_98_5/n71 ) );
  XNOR2_X2 \add_98_5/U195  ( .A(\add_98_5/n69 ), .B(\add_98_5/n70 ), .ZN(N162)
         );
  NAND2_X2 \add_98_5/U194  ( .A1(rnd_q[6]), .A2(cv_q[6]), .ZN(\add_98_5/n59 )
         );
  NAND2_X2 \add_98_5/U193  ( .A1(\add_98_5/n59 ), .A2(\add_98_5/n5 ), .ZN(
        \add_98_5/n62 ) );
  NAND2_X2 \add_98_5/U192  ( .A1(\add_98_5/n33 ), .A2(\add_98_5/n67 ), .ZN(
        \add_98_5/n66 ) );
  NAND2_X2 \add_98_5/U191  ( .A1(\add_98_5/n65 ), .A2(\add_98_5/n66 ), .ZN(
        \add_98_5/n63 ) );
  NAND2_X2 \add_98_5/U190  ( .A1(\add_98_5/n63 ), .A2(\add_98_5/n64 ), .ZN(
        \add_98_5/n60 ) );
  XNOR2_X2 \add_98_5/U189  ( .A(\add_98_5/n62 ), .B(\add_98_5/n60 ), .ZN(N163)
         );
  NAND2_X2 \add_98_5/U188  ( .A1(\add_98_5/n60 ), .A2(\add_98_5/n5 ), .ZN(
        \add_98_5/n58 ) );
  NAND2_X2 \add_98_5/U187  ( .A1(\add_98_5/n58 ), .A2(\add_98_5/n59 ), .ZN(
        \add_98_5/n55 ) );
  NAND2_X2 \add_98_5/U186  ( .A1(\add_98_5/n57 ), .A2(\add_98_5/n3 ), .ZN(
        \add_98_5/n56 ) );
  XNOR2_X2 \add_98_5/U185  ( .A(\add_98_5/n55 ), .B(\add_98_5/n56 ), .ZN(N164)
         );
  INV_X4 \add_98_5/U184  ( .A(\add_98_5/n53 ), .ZN(\add_98_5/n46 ) );
  XNOR2_X2 \add_98_5/U183  ( .A(\add_98_5/n51 ), .B(\add_98_5/n52 ), .ZN(N165)
         );
  XNOR2_X2 \add_98_5/U182  ( .A(\add_98_5/n42 ), .B(\add_98_5/n43 ), .ZN(N166)
         );
  NAND2_X2 \add_98_5/U181  ( .A1(\add_98_5/n260 ), .A2(\add_98_5/n133 ), .ZN(
        \add_98_5/n259 ) );
  NOR2_X2 \add_98_5/U180  ( .A1(\add_98_5/n20 ), .A2(\add_98_5/n109 ), .ZN(
        \add_98_5/n108 ) );
  NOR2_X2 \add_98_5/U179  ( .A1(\add_98_5/n14 ), .A2(\add_98_5/n73 ), .ZN(
        \add_98_5/n74 ) );
  NOR2_X2 \add_98_5/U178  ( .A1(\add_98_5/n262 ), .A2(\add_98_5/n136 ), .ZN(
        \add_98_5/n261 ) );
  AND2_X2 \add_98_5/U177  ( .A1(cv_q[8]), .A2(rnd_q[8]), .ZN(\add_98_5/n354 )
         );
  NOR2_X2 \add_98_5/U176  ( .A1(cv_q[9]), .A2(rnd_q[9]), .ZN(\add_98_5/n356 )
         );
  NOR2_X2 \add_98_5/U175  ( .A1(cv_q[10]), .A2(rnd_q[10]), .ZN(\add_98_5/n357 ) );
  NOR2_X2 \add_98_5/U174  ( .A1(\add_98_5/n356 ), .A2(\add_98_5/n357 ), .ZN(
        \add_98_5/n355 ) );
  NOR2_X2 \add_98_5/U173  ( .A1(\add_98_5/n47 ), .A2(\add_98_5/n46 ), .ZN(
        \add_98_5/n52 ) );
  NOR2_X2 \add_98_5/U172  ( .A1(\add_98_5/n77 ), .A2(\add_98_5/n78 ), .ZN(
        \add_98_5/n76 ) );
  AND2_X2 \add_98_5/U171  ( .A1(rnd_q[2]), .A2(cv_q[2]), .ZN(\add_98_5/n41 )
         );
  AND2_X2 \add_98_5/U170  ( .A1(rnd_q[9]), .A2(cv_q[9]), .ZN(\add_98_5/n40 )
         );
  OR2_X2 \add_98_5/U169  ( .A1(cv_q[17]), .A2(rnd_q[17]), .ZN(\add_98_5/n39 )
         );
  NOR2_X2 \add_98_5/U168  ( .A1(cv_q[17]), .A2(rnd_q[17]), .ZN(\add_98_5/n280 ) );
  NOR2_X2 \add_98_5/U167  ( .A1(\add_98_5/n280 ), .A2(\add_98_5/n281 ), .ZN(
        \add_98_5/n273 ) );
  NOR2_X2 \add_98_5/U166  ( .A1(cv_q[5]), .A2(rnd_q[5]), .ZN(\add_98_5/n297 )
         );
  NOR2_X2 \add_98_5/U165  ( .A1(cv_q[6]), .A2(rnd_q[6]), .ZN(\add_98_5/n298 )
         );
  NOR2_X2 \add_98_5/U164  ( .A1(\add_98_5/n297 ), .A2(\add_98_5/n298 ), .ZN(
        \add_98_5/n225 ) );
  NOR2_X2 \add_98_5/U163  ( .A1(\add_98_5/n309 ), .A2(\add_98_5/n313 ), .ZN(
        \add_98_5/n311 ) );
  NOR2_X2 \add_98_5/U162  ( .A1(\add_98_5/n22 ), .A2(\add_98_5/n252 ), .ZN(
        \add_98_5/n253 ) );
  NOR2_X2 \add_98_5/U161  ( .A1(\add_98_5/n41 ), .A2(\add_98_5/n80 ), .ZN(
        \add_98_5/n135 ) );
  NOR2_X2 \add_98_5/U160  ( .A1(\add_98_5/n344 ), .A2(\add_98_5/n319 ), .ZN(
        \add_98_5/n343 ) );
  NOR2_X2 \add_98_5/U159  ( .A1(\add_98_5/n244 ), .A2(\add_98_5/n250 ), .ZN(
        \add_98_5/n249 ) );
  NOR2_X2 \add_98_5/U158  ( .A1(\add_98_5/n40 ), .A2(\add_98_5/n44 ), .ZN(
        \add_98_5/n43 ) );
  NOR2_X2 \add_98_5/U157  ( .A1(\add_98_5/n71 ), .A2(\add_98_5/n68 ), .ZN(
        \add_98_5/n70 ) );
  NOR2_X2 \add_98_5/U156  ( .A1(\add_98_5/n318 ), .A2(\add_98_5/n15 ), .ZN(
        \add_98_5/n320 ) );
  AND2_X2 \add_98_5/U155  ( .A1(\add_98_5/n57 ), .A2(\add_98_5/n377 ), .ZN(
        \add_98_5/n38 ) );
  NOR2_X2 \add_98_5/U154  ( .A1(cv_q[5]), .A2(rnd_q[5]), .ZN(\add_98_5/n386 )
         );
  NOR2_X2 \add_98_5/U153  ( .A1(cv_q[21]), .A2(rnd_q[21]), .ZN(\add_98_5/n244 ) );
  NOR2_X2 \add_98_5/U152  ( .A1(cv_q[17]), .A2(rnd_q[17]), .ZN(\add_98_5/n283 ) );
  NOR2_X2 \add_98_5/U151  ( .A1(cv_q[3]), .A2(rnd_q[3]), .ZN(\add_98_5/n77 )
         );
  NOR2_X2 \add_98_5/U150  ( .A1(cv_q[2]), .A2(rnd_q[2]), .ZN(\add_98_5/n80 )
         );
  NOR2_X2 \add_98_5/U149  ( .A1(cv_q[1]), .A2(rnd_q[1]), .ZN(\add_98_5/n136 )
         );
  NOR2_X2 \add_98_5/U148  ( .A1(cv_q[20]), .A2(rnd_q[20]), .ZN(\add_98_5/n252 ) );
  NAND3_X2 \add_98_5/U147  ( .A1(cv_q[20]), .A2(rnd_q[20]), .A3(
        \add_98_5/n243 ), .ZN(\add_98_5/n202 ) );
  NOR2_X2 \add_98_5/U146  ( .A1(cv_q[16]), .A2(rnd_q[16]), .ZN(\add_98_5/n281 ) );
  NOR2_X2 \add_98_5/U145  ( .A1(cv_q[6]), .A2(rnd_q[6]), .ZN(\add_98_5/n61 )
         );
  NOR2_X2 \add_98_5/U144  ( .A1(cv_q[24]), .A2(rnd_q[24]), .ZN(\add_98_5/n180 ) );
  NOR2_X2 \add_98_5/U143  ( .A1(cv_q[5]), .A2(rnd_q[5]), .ZN(\add_98_5/n68 )
         );
  NOR2_X2 \add_98_5/U142  ( .A1(\add_98_5/n77 ), .A2(\add_98_5/n382 ), .ZN(
        \add_98_5/n218 ) );
  NOR2_X2 \add_98_5/U141  ( .A1(cv_q[14]), .A2(rnd_q[14]), .ZN(\add_98_5/n309 ) );
  NOR3_X2 \add_98_5/U140  ( .A1(\add_98_5/n308 ), .A2(\add_98_5/n309 ), .A3(
        \add_98_5/n310 ), .ZN(\add_98_5/n307 ) );
  NOR2_X2 \add_98_5/U139  ( .A1(cv_q[20]), .A2(rnd_q[20]), .ZN(\add_98_5/n247 ) );
  NOR2_X2 \add_98_5/U138  ( .A1(cv_q[21]), .A2(rnd_q[21]), .ZN(\add_98_5/n246 ) );
  NOR2_X2 \add_98_5/U137  ( .A1(\add_98_5/n246 ), .A2(\add_98_5/n247 ), .ZN(
        \add_98_5/n236 ) );
  NOR2_X2 \add_98_5/U136  ( .A1(cv_q[10]), .A2(rnd_q[10]), .ZN(\add_98_5/n352 ) );
  NOR2_X2 \add_98_5/U135  ( .A1(cv_q[8]), .A2(rnd_q[8]), .ZN(\add_98_5/n47 )
         );
  NOR2_X2 \add_98_5/U134  ( .A1(cv_q[9]), .A2(rnd_q[9]), .ZN(\add_98_5/n44 )
         );
  NOR2_X2 \add_98_5/U133  ( .A1(cv_q[12]), .A2(rnd_q[12]), .ZN(\add_98_5/n319 ) );
  NOR2_X2 \add_98_5/U132  ( .A1(cv_q[13]), .A2(rnd_q[13]), .ZN(\add_98_5/n310 ) );
  NAND3_X2 \add_98_5/U131  ( .A1(\add_98_5/n201 ), .A2(\add_98_5/n202 ), .A3(
        \add_98_5/n203 ), .ZN(\add_98_5/n200 ) );
  AND2_X4 \add_98_5/U130  ( .A1(\add_98_5/n198 ), .A2(\add_98_5/n199 ), .ZN(
        \add_98_5/n37 ) );
  AND2_X2 \add_98_5/U129  ( .A1(\add_98_5/n200 ), .A2(\add_98_5/n37 ), .ZN(
        \add_98_5/n145 ) );
  NOR2_X2 \add_98_5/U128  ( .A1(\add_98_5/n18 ), .A2(\add_98_5/n152 ), .ZN(
        \add_98_5/n153 ) );
  NOR2_X2 \add_98_5/U127  ( .A1(\add_98_5/n263 ), .A2(\add_98_5/n218 ), .ZN(
        \add_98_5/n303 ) );
  NOR2_X2 \add_98_5/U126  ( .A1(\add_98_5/n96 ), .A2(\add_98_5/n97 ), .ZN(
        \add_98_5/n85 ) );
  OR2_X4 \add_98_5/U125  ( .A1(\add_98_5/n106 ), .A2(\add_98_5/n102 ), .ZN(
        \add_98_5/n36 ) );
  AND2_X2 \add_98_5/U124  ( .A1(\add_98_5/n92 ), .A2(\add_98_5/n36 ), .ZN(
        \add_98_5/n116 ) );
  NAND3_X2 \add_98_5/U123  ( .A1(\add_98_5/n378 ), .A2(\add_98_5/n372 ), .A3(
        \add_98_5/n379 ), .ZN(\add_98_5/n370 ) );
  NOR2_X2 \add_98_5/U122  ( .A1(\add_98_5/n40 ), .A2(\add_98_5/n389 ), .ZN(
        \add_98_5/n369 ) );
  NAND3_X2 \add_98_5/U121  ( .A1(\add_98_5/n369 ), .A2(\add_98_5/n370 ), .A3(
        \add_98_5/n371 ), .ZN(\add_98_5/n367 ) );
  NAND3_X2 \add_98_5/U120  ( .A1(\add_98_5/n337 ), .A2(\add_98_5/n4 ), .A3(
        \add_98_5/n6 ), .ZN(\add_98_5/n336 ) );
  NAND3_X2 \add_98_5/U119  ( .A1(\add_98_5/n26 ), .A2(\add_98_5/n330 ), .A3(
        \add_98_5/n336 ), .ZN(\add_98_5/n334 ) );
  NOR2_X2 \add_98_5/U118  ( .A1(\add_98_5/n80 ), .A2(\add_98_5/n81 ), .ZN(
        \add_98_5/n79 ) );
  NOR2_X2 \add_98_5/U117  ( .A1(\add_98_5/n79 ), .A2(\add_98_5/n41 ), .ZN(
        \add_98_5/n75 ) );
  NOR2_X2 \add_98_5/U116  ( .A1(\add_98_5/n235 ), .A2(\add_98_5/n245 ), .ZN(
        \add_98_5/n241 ) );
  NOR2_X2 \add_98_5/U115  ( .A1(\add_98_5/n241 ), .A2(\add_98_5/n242 ), .ZN(
        \add_98_5/n238 ) );
  NOR2_X2 \add_98_5/U114  ( .A1(\add_98_5/n33 ), .A2(\add_98_5/n50 ), .ZN(
        \add_98_5/n49 ) );
  NOR2_X2 \add_98_5/U113  ( .A1(\add_98_5/n49 ), .A2(\add_98_5/n19 ), .ZN(
        \add_98_5/n48 ) );
  NOR2_X2 \add_98_5/U112  ( .A1(\add_98_5/n47 ), .A2(\add_98_5/n48 ), .ZN(
        \add_98_5/n45 ) );
  NOR2_X2 \add_98_5/U111  ( .A1(\add_98_5/n45 ), .A2(\add_98_5/n46 ), .ZN(
        \add_98_5/n42 ) );
  NOR2_X2 \add_98_5/U110  ( .A1(\add_98_5/n252 ), .A2(\add_98_5/n235 ), .ZN(
        \add_98_5/n251 ) );
  NOR2_X2 \add_98_5/U109  ( .A1(\add_98_5/n251 ), .A2(\add_98_5/n22 ), .ZN(
        \add_98_5/n248 ) );
  NOR2_X2 \add_98_5/U108  ( .A1(\add_98_5/n33 ), .A2(\add_98_5/n14 ), .ZN(
        \add_98_5/n72 ) );
  NOR2_X2 \add_98_5/U107  ( .A1(\add_98_5/n72 ), .A2(\add_98_5/n73 ), .ZN(
        \add_98_5/n69 ) );
  NOR2_X2 \add_98_5/U106  ( .A1(\add_98_5/n61 ), .A2(\add_98_5/n68 ), .ZN(
        \add_98_5/n375 ) );
  NOR2_X2 \add_98_5/U105  ( .A1(\add_98_5/n348 ), .A2(\add_98_5/n349 ), .ZN(
        \add_98_5/n347 ) );
  NAND3_X2 \add_98_5/U104  ( .A1(\add_98_5/n346 ), .A2(\add_98_5/n16 ), .A3(
        \add_98_5/n347 ), .ZN(\add_98_5/n316 ) );
  NOR2_X2 \add_98_5/U103  ( .A1(\add_98_5/n14 ), .A2(\add_98_5/n68 ), .ZN(
        \add_98_5/n65 ) );
  NAND3_X2 \add_98_5/U102  ( .A1(\add_98_5/n314 ), .A2(\add_98_5/n315 ), .A3(
        \add_98_5/n316 ), .ZN(\add_98_5/n132 ) );
  NOR2_X2 \add_98_5/U101  ( .A1(\add_98_5/n20 ), .A2(\add_98_5/n92 ), .ZN(
        \add_98_5/n91 ) );
  NOR2_X2 \add_98_5/U100  ( .A1(\add_98_5/n319 ), .A2(\add_98_5/n23 ), .ZN(
        \add_98_5/n325 ) );
  NAND3_X2 \add_98_5/U99  ( .A1(\add_98_5/n160 ), .A2(\add_98_5/n8 ), .A3(
        \add_98_5/n161 ), .ZN(\add_98_5/n159 ) );
  NAND3_X2 \add_98_5/U98  ( .A1(\add_98_5/n158 ), .A2(\add_98_5/n149 ), .A3(
        \add_98_5/n159 ), .ZN(\add_98_5/n156 ) );
  NOR2_X2 \add_98_5/U97  ( .A1(\add_98_5/n44 ), .A2(\add_98_5/n53 ), .ZN(
        \add_98_5/n389 ) );
  NAND3_X2 \add_98_5/U96  ( .A1(\add_98_5/n215 ), .A2(\add_98_5/n216 ), .A3(
        \add_98_5/n217 ), .ZN(\add_98_5/n211 ) );
  NOR3_X2 \add_98_5/U95  ( .A1(\add_98_5/n134 ), .A2(\add_98_5/n129 ), .A3(
        \add_98_5/n130 ), .ZN(\add_98_5/n127 ) );
  NOR2_X2 \add_98_5/U94  ( .A1(\add_98_5/n127 ), .A2(\add_98_5/n128 ), .ZN(
        \add_98_5/n123 ) );
  NOR2_X2 \add_98_5/U93  ( .A1(\add_98_5/n123 ), .A2(\add_98_5/n124 ), .ZN(
        \add_98_5/n120 ) );
  NOR3_X2 \add_98_5/U92  ( .A1(\add_98_5/n179 ), .A2(\add_98_5/n177 ), .A3(
        \add_98_5/n180 ), .ZN(\add_98_5/n175 ) );
  NOR2_X2 \add_98_5/U91  ( .A1(\add_98_5/n175 ), .A2(\add_98_5/n176 ), .ZN(
        \add_98_5/n172 ) );
  OR2_X4 \add_98_5/U90  ( .A1(\add_98_5/n136 ), .A2(\add_98_5/n221 ), .ZN(
        \add_98_5/n35 ) );
  AND2_X2 \add_98_5/U89  ( .A1(\add_98_5/n137 ), .A2(\add_98_5/n35 ), .ZN(
        \add_98_5/n81 ) );
  AND3_X2 \add_98_5/U88  ( .A1(\add_98_5/n170 ), .A2(\add_98_5/n158 ), .A3(
        \add_98_5/n171 ), .ZN(\add_98_5/n34 ) );
  NAND3_X2 \add_98_5/U87  ( .A1(\add_98_5/n149 ), .A2(\add_98_5/n150 ), .A3(
        \add_98_5/n34 ), .ZN(\add_98_5/n121 ) );
  NOR2_X2 \add_98_5/U86  ( .A1(\add_98_5/n319 ), .A2(\add_98_5/n23 ), .ZN(
        \add_98_5/n337 ) );
  NOR2_X2 \add_98_5/U85  ( .A1(\add_98_5/n47 ), .A2(\add_98_5/n44 ), .ZN(
        \add_98_5/n372 ) );
  AND3_X2 \add_98_5/U84  ( .A1(\add_98_5/n217 ), .A2(\add_98_5/n215 ), .A3(
        \add_98_5/n380 ), .ZN(\add_98_5/n33 ) );
  NOR2_X2 \add_98_5/U83  ( .A1(\add_98_5/n14 ), .A2(\add_98_5/n386 ), .ZN(
        \add_98_5/n385 ) );
  NAND3_X2 \add_98_5/U82  ( .A1(\add_98_5/n3 ), .A2(\add_98_5/n5 ), .A3(
        \add_98_5/n385 ), .ZN(\add_98_5/n50 ) );
  NOR3_X2 \add_98_5/U81  ( .A1(\add_98_5/n120 ), .A2(\add_98_5/n121 ), .A3(
        \add_98_5/n122 ), .ZN(\add_98_5/n112 ) );
  NOR2_X2 \add_98_5/U80  ( .A1(\add_98_5/n112 ), .A2(\add_98_5/n113 ), .ZN(
        \add_98_5/n107 ) );
  NOR2_X2 \add_98_5/U79  ( .A1(\add_98_5/n20 ), .A2(\add_98_5/n106 ), .ZN(
        \add_98_5/n95 ) );
  NAND3_X2 \add_98_5/U78  ( .A1(\add_98_5/n234 ), .A2(\add_98_5/n203 ), .A3(
        \add_98_5/n17 ), .ZN(\add_98_5/n230 ) );
  NOR2_X2 \add_98_5/U77  ( .A1(\add_98_5/n213 ), .A2(\add_98_5/n214 ), .ZN(
        \add_98_5/n293 ) );
  NAND3_X2 \add_98_5/U76  ( .A1(\add_98_5/n161 ), .A2(\add_98_5/n8 ), .A3(
        \add_98_5/n160 ), .ZN(\add_98_5/n169 ) );
  NOR2_X2 \add_98_5/U75  ( .A1(\add_98_5/n146 ), .A2(\add_98_5/n126 ), .ZN(
        \add_98_5/n192 ) );
  NOR2_X2 \add_98_5/U74  ( .A1(\add_98_5/n209 ), .A2(\add_98_5/n210 ), .ZN(
        \add_98_5/n208 ) );
  NAND3_X2 \add_98_5/U73  ( .A1(\add_98_5/n211 ), .A2(\add_98_5/n212 ), .A3(
        \add_98_5/n378 ), .ZN(\add_98_5/n207 ) );
  NAND3_X2 \add_98_5/U72  ( .A1(\add_98_5/n207 ), .A2(\add_98_5/n208 ), .A3(
        \add_98_5/n206 ), .ZN(\add_98_5/n205 ) );
  NOR3_X2 \add_98_5/U71  ( .A1(\add_98_5/n259 ), .A2(\add_98_5/n210 ), .A3(
        \add_98_5/n209 ), .ZN(\add_98_5/n256 ) );
  NOR2_X2 \add_98_5/U70  ( .A1(\add_98_5/n256 ), .A2(\add_98_5/n128 ), .ZN(
        \add_98_5/n254 ) );
  NOR2_X2 \add_98_5/U69  ( .A1(\add_98_5/n254 ), .A2(\add_98_5/n255 ), .ZN(
        \add_98_5/n235 ) );
  NOR3_X2 \add_98_5/U68  ( .A1(\add_98_5/n218 ), .A2(\add_98_5/n78 ), .A3(
        \add_98_5/n1 ), .ZN(\add_98_5/n302 ) );
  NOR2_X2 \add_98_5/U67  ( .A1(\add_98_5/n318 ), .A2(\add_98_5/n319 ), .ZN(
        \add_98_5/n317 ) );
  NAND3_X2 \add_98_5/U66  ( .A1(\add_98_5/n4 ), .A2(\add_98_5/n9 ), .A3(
        \add_98_5/n317 ), .ZN(\add_98_5/n213 ) );
  NOR3_X2 \add_98_5/U65  ( .A1(\add_98_5/n193 ), .A2(\add_98_5/n146 ), .A3(
        \add_98_5/n194 ), .ZN(\add_98_5/n191 ) );
  OR3_X4 \add_98_5/U64  ( .A1(\add_98_5/n311 ), .A2(\add_98_5/n312 ), .A3(
        \add_98_5/n15 ), .ZN(\add_98_5/n32 ) );
  OR2_X2 \add_98_5/U63  ( .A1(\add_98_5/n32 ), .A2(\add_98_5/n307 ), .ZN(
        \add_98_5/n305 ) );
  NOR2_X2 \add_98_5/U62  ( .A1(\add_98_5/n352 ), .A2(\add_98_5/n362 ), .ZN(
        \add_98_5/n361 ) );
  NAND3_X2 \add_98_5/U61  ( .A1(\add_98_5/n359 ), .A2(\add_98_5/n360 ), .A3(
        \add_98_5/n361 ), .ZN(\add_98_5/n214 ) );
  NOR2_X2 \add_98_5/U60  ( .A1(\add_98_5/n262 ), .A2(\add_98_5/n78 ), .ZN(
        \add_98_5/n304 ) );
  NOR2_X2 \add_98_5/U59  ( .A1(\add_98_5/n325 ), .A2(\add_98_5/n326 ), .ZN(
        \add_98_5/n324 ) );
  NOR3_X2 \add_98_5/U58  ( .A1(\add_98_5/n323 ), .A2(\add_98_5/n324 ), .A3(
        \add_98_5/n24 ), .ZN(\add_98_5/n322 ) );
  NOR2_X2 \add_98_5/U57  ( .A1(\add_98_5/n312 ), .A2(\add_98_5/n322 ), .ZN(
        \add_98_5/n321 ) );
  NOR2_X2 \add_98_5/U56  ( .A1(\add_98_5/n33 ), .A2(\add_98_5/n50 ), .ZN(
        \add_98_5/n54 ) );
  NOR2_X2 \add_98_5/U55  ( .A1(\add_98_5/n54 ), .A2(\add_98_5/n19 ), .ZN(
        \add_98_5/n51 ) );
  NOR2_X2 \add_98_5/U54  ( .A1(\add_98_5/n272 ), .A2(\add_98_5/n258 ), .ZN(
        \add_98_5/n267 ) );
  NOR2_X2 \add_98_5/U53  ( .A1(\add_98_5/n267 ), .A2(\add_98_5/n196 ), .ZN(
        \add_98_5/n264 ) );
  NOR2_X2 \add_98_5/U52  ( .A1(\add_98_5/n33 ), .A2(\add_98_5/n50 ), .ZN(
        \add_98_5/n363 ) );
  NOR2_X2 \add_98_5/U51  ( .A1(\add_98_5/n363 ), .A2(\add_98_5/n19 ), .ZN(
        \add_98_5/n358 ) );
  NOR2_X2 \add_98_5/U50  ( .A1(\add_98_5/n358 ), .A2(\add_98_5/n214 ), .ZN(
        \add_98_5/n345 ) );
  NOR2_X2 \add_98_5/U49  ( .A1(\add_98_5/n345 ), .A2(\add_98_5/n328 ), .ZN(
        \add_98_5/n342 ) );
  NOR2_X2 \add_98_5/U48  ( .A1(\add_98_5/n93 ), .A2(\add_98_5/n94 ), .ZN(
        \add_98_5/n90 ) );
  NOR2_X2 \add_98_5/U47  ( .A1(\add_98_5/n213 ), .A2(\add_98_5/n214 ), .ZN(
        \add_98_5/n212 ) );
  NOR2_X2 \add_98_5/U46  ( .A1(\add_98_5/n33 ), .A2(\add_98_5/n50 ), .ZN(
        \add_98_5/n327 ) );
  NAND3_X2 \add_98_5/U45  ( .A1(\add_98_5/n89 ), .A2(\add_98_5/n13 ), .A3(
        \add_98_5/n88 ), .ZN(\add_98_5/n143 ) );
  NOR3_X2 \add_98_5/U44  ( .A1(\add_98_5/n11 ), .A2(\add_98_5/n21 ), .A3(
        \add_98_5/n147 ), .ZN(\add_98_5/n142 ) );
  NAND3_X2 \add_98_5/U43  ( .A1(\add_98_5/n88 ), .A2(\add_98_5/n89 ), .A3(
        \add_98_5/n12 ), .ZN(\add_98_5/n87 ) );
  NOR2_X2 \add_98_5/U42  ( .A1(\add_98_5/n90 ), .A2(\add_98_5/n91 ), .ZN(
        \add_98_5/n86 ) );
  NOR4_X2 \add_98_5/U41  ( .A1(\add_98_5/n327 ), .A2(\add_98_5/n328 ), .A3(
        \add_98_5/n19 ), .A4(\add_98_5/n326 ), .ZN(\add_98_5/n323 ) );
  NOR2_X2 \add_98_5/U40  ( .A1(\add_98_5/n50 ), .A2(\add_98_5/n302 ), .ZN(
        \add_98_5/n301 ) );
  NOR2_X2 \add_98_5/U39  ( .A1(\add_98_5/n213 ), .A2(\add_98_5/n214 ), .ZN(
        \add_98_5/n299 ) );
  NAND3_X2 \add_98_5/U38  ( .A1(\add_98_5/n299 ), .A2(\add_98_5/n300 ), .A3(
        \add_98_5/n301 ), .ZN(\add_98_5/n133 ) );
  NOR2_X2 \add_98_5/U37  ( .A1(\add_98_5/n128 ), .A2(\add_98_5/n146 ), .ZN(
        \add_98_5/n204 ) );
  NOR3_X2 \add_98_5/U36  ( .A1(\add_98_5/n190 ), .A2(\add_98_5/n191 ), .A3(
        \add_98_5/n192 ), .ZN(\add_98_5/n189 ) );
  NOR2_X2 \add_98_5/U35  ( .A1(\add_98_5/n210 ), .A2(\add_98_5/n209 ), .ZN(
        \add_98_5/n291 ) );
  NAND3_X2 \add_98_5/U34  ( .A1(\add_98_5/n291 ), .A2(\add_98_5/n133 ), .A3(
        \add_98_5/n260 ), .ZN(\add_98_5/n89 ) );
  OR2_X4 \add_98_5/U33  ( .A1(rnd_q[11]), .A2(cv_q[11]), .ZN(\add_98_5/n315 )
         );
  OR2_X4 \add_98_5/U32  ( .A1(\add_98_5/n283 ), .A2(\add_98_5/n284 ), .ZN(
        \add_98_5/n31 ) );
  AND2_X4 \add_98_5/U31  ( .A1(\add_98_5/n381 ), .A2(\add_98_5/n221 ), .ZN(
        N157) );
  AND2_X4 \add_98_5/U30  ( .A1(\add_98_5/n150 ), .A2(\add_98_5/n102 ), .ZN(
        \add_98_5/n29 ) );
  AND2_X4 \add_98_5/U29  ( .A1(\add_98_5/n198 ), .A2(\add_98_5/n203 ), .ZN(
        \add_98_5/n28 ) );
  AND2_X4 \add_98_5/U28  ( .A1(\add_98_5/n158 ), .A2(\add_98_5/n161 ), .ZN(
        \add_98_5/n27 ) );
  OR2_X4 \add_98_5/U27  ( .A1(\add_98_5/n310 ), .A2(\add_98_5/n329 ), .ZN(
        \add_98_5/n26 ) );
  AND2_X4 \add_98_5/U26  ( .A1(\add_98_5/n126 ), .A2(\add_98_5/n195 ), .ZN(
        \add_98_5/n25 ) );
  OR2_X4 \add_98_5/U25  ( .A1(\add_98_5/n309 ), .A2(\add_98_5/n310 ), .ZN(
        \add_98_5/n24 ) );
  AND2_X4 \add_98_5/U24  ( .A1(\add_98_5/n214 ), .A2(\add_98_5/n341 ), .ZN(
        \add_98_5/n23 ) );
  AND2_X4 \add_98_5/U23  ( .A1(rnd_q[20]), .A2(cv_q[20]), .ZN(\add_98_5/n22 )
         );
  AND2_X4 \add_98_5/U22  ( .A1(\add_98_5/n148 ), .A2(\add_98_5/n105 ), .ZN(
        \add_98_5/n21 ) );
  AND2_X4 \add_98_5/U21  ( .A1(\add_98_5/n110 ), .A2(\add_98_5/n111 ), .ZN(
        \add_98_5/n20 ) );
  AND2_X4 \add_98_5/U20  ( .A1(\add_98_5/n373 ), .A2(\add_98_5/n3 ), .ZN(
        \add_98_5/n19 ) );
  AND3_X4 \add_98_5/U19  ( .A1(\add_98_5/n34 ), .A2(\add_98_5/n149 ), .A3(
        \add_98_5/n162 ), .ZN(\add_98_5/n18 ) );
  OR2_X4 \add_98_5/U18  ( .A1(\add_98_5/n235 ), .A2(\add_98_5/n229 ), .ZN(
        \add_98_5/n17 ) );
  OR2_X4 \add_98_5/U17  ( .A1(\add_98_5/n352 ), .A2(\add_98_5/n353 ), .ZN(
        \add_98_5/n16 ) );
  AND2_X4 \add_98_5/U16  ( .A1(rnd_q[15]), .A2(cv_q[15]), .ZN(\add_98_5/n15 )
         );
  AND2_X4 \add_98_5/U15  ( .A1(\add_98_5/n387 ), .A2(\add_98_5/n388 ), .ZN(
        \add_98_5/n14 ) );
  AND2_X4 \add_98_5/U14  ( .A1(\add_98_5/n104 ), .A2(\add_98_5/n105 ), .ZN(
        \add_98_5/n13 ) );
  AND3_X4 \add_98_5/U13  ( .A1(\add_98_5/n104 ), .A2(\add_98_5/n95 ), .A3(
        \add_98_5/n105 ), .ZN(\add_98_5/n12 ) );
  AND2_X4 \add_98_5/U12  ( .A1(\add_98_5/n152 ), .A2(\add_98_5/n150 ), .ZN(
        \add_98_5/n11 ) );
  OR2_X4 \add_98_5/U11  ( .A1(cv_q[3]), .A2(rnd_q[3]), .ZN(\add_98_5/n10 ) );
  OR2_X4 \add_98_5/U10  ( .A1(cv_q[14]), .A2(rnd_q[14]), .ZN(\add_98_5/n9 ) );
  OR2_X4 \add_98_5/U9  ( .A1(\add_98_5/n177 ), .A2(\add_98_5/n178 ), .ZN(
        \add_98_5/n8 ) );
  OR2_X4 \add_98_5/U8  ( .A1(cv_q[2]), .A2(rnd_q[2]), .ZN(\add_98_5/n7 ) );
  OR3_X4 \add_98_5/U7  ( .A1(\add_98_5/n327 ), .A2(\add_98_5/n19 ), .A3(
        \add_98_5/n328 ), .ZN(\add_98_5/n6 ) );
  OR2_X4 \add_98_5/U6  ( .A1(cv_q[6]), .A2(rnd_q[6]), .ZN(\add_98_5/n5 ) );
  OR2_X4 \add_98_5/U5  ( .A1(cv_q[13]), .A2(rnd_q[13]), .ZN(\add_98_5/n4 ) );
  OR2_X4 \add_98_5/U4  ( .A1(cv_q[7]), .A2(rnd_q[7]), .ZN(\add_98_5/n3 ) );
  OR2_X4 \add_98_5/U3  ( .A1(cv_q[1]), .A2(rnd_q[1]), .ZN(\add_98_5/n2 ) );
  AND3_X4 \add_98_5/U2  ( .A1(\add_98_5/n7 ), .A2(\add_98_5/n10 ), .A3(
        \add_98_5/n2 ), .ZN(\add_98_5/n1 ) );
  INV_X4 \add_98/U426  ( .A(rnd_q[128]), .ZN(\add_98/n393 ) );
  INV_X4 \add_98/U425  ( .A(cv_q[128]), .ZN(\add_98/n394 ) );
  NAND2_X2 \add_98/U424  ( .A1(\add_98/n393 ), .A2(\add_98/n394 ), .ZN(
        \add_98/n383 ) );
  NAND2_X2 \add_98/U423  ( .A1(rnd_q[128]), .A2(cv_q[128]), .ZN(\add_98/n220 )
         );
  INV_X4 \add_98/U422  ( .A(\add_98/n351 ), .ZN(\add_98/n392 ) );
  NAND2_X2 \add_98/U421  ( .A1(rnd_q[138]), .A2(cv_q[138]), .ZN(\add_98/n350 )
         );
  NAND2_X2 \add_98/U420  ( .A1(\add_98/n392 ), .A2(\add_98/n350 ), .ZN(
        \add_98/n369 ) );
  NAND2_X2 \add_98/U419  ( .A1(rnd_q[136]), .A2(cv_q[136]), .ZN(\add_98/n53 )
         );
  INV_X4 \add_98/U418  ( .A(rnd_q[132]), .ZN(\add_98/n389 ) );
  INV_X4 \add_98/U417  ( .A(cv_q[132]), .ZN(\add_98/n390 ) );
  INV_X4 \add_98/U416  ( .A(\add_98/n50 ), .ZN(\add_98/n379 ) );
  NAND2_X2 \add_98/U415  ( .A1(rnd_q[129]), .A2(cv_q[129]), .ZN(\add_98/n386 )
         );
  NAND2_X2 \add_98/U414  ( .A1(\add_98/n386 ), .A2(\add_98/n220 ), .ZN(
        \add_98/n385 ) );
  NAND2_X2 \add_98/U413  ( .A1(\add_98/n1 ), .A2(\add_98/n385 ), .ZN(
        \add_98/n381 ) );
  NAND2_X2 \add_98/U412  ( .A1(cv_q[130]), .A2(rnd_q[130]), .ZN(\add_98/n384 )
         );
  INV_X4 \add_98/U411  ( .A(\add_98/n217 ), .ZN(\add_98/n382 ) );
  NAND2_X2 \add_98/U410  ( .A1(rnd_q[131]), .A2(cv_q[131]), .ZN(\add_98/n215 )
         );
  INV_X4 \add_98/U409  ( .A(\add_98/n35 ), .ZN(\add_98/n380 ) );
  NAND2_X2 \add_98/U408  ( .A1(rnd_q[135]), .A2(cv_q[135]), .ZN(\add_98/n57 )
         );
  NAND2_X2 \add_98/U407  ( .A1(rnd_q[134]), .A2(cv_q[134]), .ZN(\add_98/n378 )
         );
  NAND2_X2 \add_98/U406  ( .A1(rnd_q[132]), .A2(cv_q[132]), .ZN(\add_98/n67 )
         );
  NAND2_X2 \add_98/U405  ( .A1(rnd_q[133]), .A2(cv_q[133]), .ZN(\add_98/n64 )
         );
  NAND2_X2 \add_98/U404  ( .A1(\add_98/n67 ), .A2(\add_98/n64 ), .ZN(
        \add_98/n377 ) );
  NAND2_X2 \add_98/U403  ( .A1(\add_98/n376 ), .A2(\add_98/n377 ), .ZN(
        \add_98/n375 ) );
  NAND2_X2 \add_98/U402  ( .A1(\add_98/n22 ), .A2(\add_98/n375 ), .ZN(
        \add_98/n374 ) );
  NAND2_X2 \add_98/U401  ( .A1(\add_98/n19 ), .A2(\add_98/n373 ), .ZN(
        \add_98/n372 ) );
  XNOR2_X2 \add_98/U400  ( .A(\add_98/n369 ), .B(\add_98/n368 ), .ZN(N39) );
  NAND2_X2 \add_98/U399  ( .A1(\add_98/n368 ), .A2(\add_98/n392 ), .ZN(
        \add_98/n367 ) );
  NAND2_X2 \add_98/U398  ( .A1(\add_98/n367 ), .A2(\add_98/n350 ), .ZN(
        \add_98/n363 ) );
  NAND2_X2 \add_98/U397  ( .A1(rnd_q[139]), .A2(cv_q[139]), .ZN(\add_98/n349 )
         );
  INV_X4 \add_98/U396  ( .A(rnd_q[139]), .ZN(\add_98/n365 ) );
  INV_X4 \add_98/U395  ( .A(cv_q[139]), .ZN(\add_98/n366 ) );
  NAND2_X2 \add_98/U394  ( .A1(\add_98/n365 ), .A2(\add_98/n366 ), .ZN(
        \add_98/n314 ) );
  NAND2_X2 \add_98/U393  ( .A1(\add_98/n349 ), .A2(\add_98/n314 ), .ZN(
        \add_98/n364 ) );
  XNOR2_X2 \add_98/U392  ( .A(\add_98/n363 ), .B(\add_98/n364 ), .ZN(N40) );
  INV_X4 \add_98/U391  ( .A(\add_98/n44 ), .ZN(\add_98/n358 ) );
  INV_X4 \add_98/U390  ( .A(\add_98/n47 ), .ZN(\add_98/n359 ) );
  INV_X4 \add_98/U389  ( .A(\add_98/n314 ), .ZN(\add_98/n361 ) );
  NAND2_X2 \add_98/U388  ( .A1(\add_98/n353 ), .A2(\add_98/n354 ), .ZN(
        \add_98/n345 ) );
  NAND2_X2 \add_98/U387  ( .A1(cv_q[137]), .A2(rnd_q[137]), .ZN(\add_98/n352 )
         );
  INV_X4 \add_98/U386  ( .A(\add_98/n350 ), .ZN(\add_98/n347 ) );
  INV_X4 \add_98/U385  ( .A(\add_98/n349 ), .ZN(\add_98/n348 ) );
  NAND2_X2 \add_98/U384  ( .A1(\add_98/n315 ), .A2(\add_98/n314 ), .ZN(
        \add_98/n340 ) );
  INV_X4 \add_98/U383  ( .A(\add_98/n340 ), .ZN(\add_98/n327 ) );
  NAND2_X2 \add_98/U382  ( .A1(rnd_q[140]), .A2(cv_q[140]), .ZN(\add_98/n328 )
         );
  INV_X4 \add_98/U381  ( .A(\add_98/n328 ), .ZN(\add_98/n343 ) );
  XNOR2_X2 \add_98/U380  ( .A(\add_98/n341 ), .B(\add_98/n342 ), .ZN(N41) );
  NAND2_X2 \add_98/U379  ( .A1(\add_98/n336 ), .A2(\add_98/n6 ), .ZN(
        \add_98/n339 ) );
  NAND2_X2 \add_98/U378  ( .A1(\add_98/n339 ), .A2(\add_98/n328 ), .ZN(
        \add_98/n337 ) );
  NAND2_X2 \add_98/U377  ( .A1(rnd_q[141]), .A2(cv_q[141]), .ZN(\add_98/n329 )
         );
  NAND2_X2 \add_98/U376  ( .A1(\add_98/n329 ), .A2(\add_98/n4 ), .ZN(
        \add_98/n338 ) );
  XNOR2_X2 \add_98/U375  ( .A(\add_98/n337 ), .B(\add_98/n338 ), .ZN(N42) );
  NAND2_X2 \add_98/U374  ( .A1(rnd_q[142]), .A2(cv_q[142]), .ZN(\add_98/n330 )
         );
  NAND2_X2 \add_98/U373  ( .A1(\add_98/n9 ), .A2(\add_98/n330 ), .ZN(
        \add_98/n334 ) );
  XNOR2_X2 \add_98/U372  ( .A(\add_98/n333 ), .B(\add_98/n334 ), .ZN(N43) );
  INV_X4 \add_98/U371  ( .A(rnd_q[143]), .ZN(\add_98/n331 ) );
  INV_X4 \add_98/U370  ( .A(cv_q[143]), .ZN(\add_98/n332 ) );
  NAND2_X2 \add_98/U369  ( .A1(\add_98/n331 ), .A2(\add_98/n332 ), .ZN(
        \add_98/n305 ) );
  INV_X4 \add_98/U368  ( .A(\add_98/n305 ), .ZN(\add_98/n317 ) );
  INV_X4 \add_98/U367  ( .A(\add_98/n330 ), .ZN(\add_98/n311 ) );
  NAND2_X2 \add_98/U366  ( .A1(\add_98/n328 ), .A2(\add_98/n329 ), .ZN(
        \add_98/n325 ) );
  XNOR2_X2 \add_98/U365  ( .A(\add_98/n319 ), .B(\add_98/n320 ), .ZN(N44) );
  NAND2_X2 \add_98/U364  ( .A1(rnd_q[144]), .A2(cv_q[144]), .ZN(\add_98/n285 )
         );
  NAND2_X2 \add_98/U363  ( .A1(\add_98/n285 ), .A2(\add_98/n287 ), .ZN(
        \add_98/n288 ) );
  INV_X4 \add_98/U362  ( .A(\add_98/n213 ), .ZN(\add_98/n313 ) );
  INV_X4 \add_98/U361  ( .A(\add_98/n132 ), .ZN(\add_98/n210 ) );
  NAND2_X2 \add_98/U360  ( .A1(cv_q[141]), .A2(rnd_q[141]), .ZN(\add_98/n312 )
         );
  NAND2_X2 \add_98/U359  ( .A1(rnd_q[140]), .A2(cv_q[140]), .ZN(\add_98/n307 )
         );
  NAND2_X2 \add_98/U358  ( .A1(\add_98/n304 ), .A2(\add_98/n305 ), .ZN(
        \add_98/n131 ) );
  INV_X4 \add_98/U357  ( .A(\add_98/n131 ), .ZN(\add_98/n209 ) );
  INV_X4 \add_98/U356  ( .A(\add_98/n220 ), .ZN(\add_98/n303 ) );
  NAND2_X2 \add_98/U355  ( .A1(rnd_q[129]), .A2(cv_q[129]), .ZN(\add_98/n137 )
         );
  INV_X4 \add_98/U354  ( .A(\add_98/n137 ), .ZN(\add_98/n261 ) );
  INV_X4 \add_98/U353  ( .A(\add_98/n215 ), .ZN(\add_98/n78 ) );
  NAND2_X2 \add_98/U352  ( .A1(\add_98/n301 ), .A2(\add_98/n302 ), .ZN(
        \add_98/n298 ) );
  NAND2_X2 \add_98/U351  ( .A1(rnd_q[133]), .A2(cv_q[133]), .ZN(\add_98/n294 )
         );
  NAND2_X2 \add_98/U350  ( .A1(\add_98/n67 ), .A2(\add_98/n294 ), .ZN(
        \add_98/n293 ) );
  NAND2_X2 \add_98/U349  ( .A1(\add_98/n224 ), .A2(\add_98/n293 ), .ZN(
        \add_98/n292 ) );
  NAND2_X2 \add_98/U348  ( .A1(\add_98/n22 ), .A2(\add_98/n292 ), .ZN(
        \add_98/n290 ) );
  NAND3_X2 \add_98/U347  ( .A1(\add_98/n290 ), .A2(\add_98/n3 ), .A3(
        \add_98/n291 ), .ZN(\add_98/n259 ) );
  INV_X4 \add_98/U346  ( .A(\add_98/n259 ), .ZN(\add_98/n134 ) );
  XNOR2_X2 \add_98/U345  ( .A(\add_98/n288 ), .B(\add_98/n89 ), .ZN(N45) );
  INV_X4 \add_98/U344  ( .A(\add_98/n279 ), .ZN(\add_98/n287 ) );
  NAND2_X2 \add_98/U343  ( .A1(\add_98/n89 ), .A2(\add_98/n287 ), .ZN(
        \add_98/n286 ) );
  NAND2_X2 \add_98/U342  ( .A1(\add_98/n285 ), .A2(\add_98/n286 ), .ZN(
        \add_98/n283 ) );
  NAND2_X2 \add_98/U341  ( .A1(rnd_q[145]), .A2(cv_q[145]), .ZN(\add_98/n280 )
         );
  NAND2_X2 \add_98/U340  ( .A1(\add_98/n41 ), .A2(\add_98/n280 ), .ZN(
        \add_98/n284 ) );
  XNOR2_X2 \add_98/U339  ( .A(\add_98/n283 ), .B(\add_98/n284 ), .ZN(N46) );
  NAND2_X2 \add_98/U338  ( .A1(cv_q[144]), .A2(rnd_q[144]), .ZN(\add_98/n282 )
         );
  NAND2_X2 \add_98/U337  ( .A1(\add_98/n40 ), .A2(\add_98/n280 ), .ZN(
        \add_98/n268 ) );
  INV_X4 \add_98/U336  ( .A(\add_98/n268 ), .ZN(\add_98/n276 ) );
  NAND2_X2 \add_98/U335  ( .A1(\add_98/n271 ), .A2(\add_98/n89 ), .ZN(
        \add_98/n277 ) );
  NAND2_X2 \add_98/U334  ( .A1(\add_98/n276 ), .A2(\add_98/n277 ), .ZN(
        \add_98/n272 ) );
  NAND2_X2 \add_98/U333  ( .A1(rnd_q[146]), .A2(cv_q[146]), .ZN(\add_98/n267 )
         );
  INV_X4 \add_98/U332  ( .A(rnd_q[146]), .ZN(\add_98/n274 ) );
  INV_X4 \add_98/U331  ( .A(cv_q[146]), .ZN(\add_98/n275 ) );
  NAND2_X2 \add_98/U330  ( .A1(\add_98/n274 ), .A2(\add_98/n275 ), .ZN(
        \add_98/n269 ) );
  NAND2_X2 \add_98/U329  ( .A1(\add_98/n267 ), .A2(\add_98/n269 ), .ZN(
        \add_98/n273 ) );
  XNOR2_X2 \add_98/U328  ( .A(\add_98/n272 ), .B(\add_98/n273 ), .ZN(N47) );
  INV_X4 \add_98/U327  ( .A(\add_98/n89 ), .ZN(\add_98/n270 ) );
  NAND2_X2 \add_98/U326  ( .A1(\add_98/n271 ), .A2(\add_98/n269 ), .ZN(
        \add_98/n257 ) );
  NAND2_X2 \add_98/U325  ( .A1(\add_98/n268 ), .A2(\add_98/n269 ), .ZN(
        \add_98/n266 ) );
  NAND2_X2 \add_98/U324  ( .A1(\add_98/n266 ), .A2(\add_98/n267 ), .ZN(
        \add_98/n196 ) );
  NAND2_X2 \add_98/U323  ( .A1(rnd_q[147]), .A2(cv_q[147]), .ZN(\add_98/n126 )
         );
  INV_X4 \add_98/U322  ( .A(rnd_q[147]), .ZN(\add_98/n263 ) );
  INV_X4 \add_98/U321  ( .A(cv_q[147]), .ZN(\add_98/n264 ) );
  NAND2_X2 \add_98/U320  ( .A1(\add_98/n263 ), .A2(\add_98/n264 ), .ZN(
        \add_98/n195 ) );
  XNOR2_X2 \add_98/U319  ( .A(\add_98/n262 ), .B(\add_98/n28 ), .ZN(N48) );
  XNOR2_X2 \add_98/U318  ( .A(\add_98/n220 ), .B(\add_98/n260 ), .ZN(N30) );
  INV_X4 \add_98/U317  ( .A(\add_98/n257 ), .ZN(\add_98/n256 ) );
  NAND2_X2 \add_98/U316  ( .A1(\add_98/n256 ), .A2(\add_98/n195 ), .ZN(
        \add_98/n128 ) );
  NAND2_X2 \add_98/U315  ( .A1(\add_98/n196 ), .A2(\add_98/n195 ), .ZN(
        \add_98/n125 ) );
  NAND2_X2 \add_98/U314  ( .A1(\add_98/n125 ), .A2(\add_98/n126 ), .ZN(
        \add_98/n254 ) );
  XNOR2_X2 \add_98/U313  ( .A(\add_98/n234 ), .B(\add_98/n252 ), .ZN(N49) );
  NAND2_X2 \add_98/U312  ( .A1(rnd_q[149]), .A2(cv_q[149]), .ZN(\add_98/n201 )
         );
  INV_X4 \add_98/U311  ( .A(\add_98/n201 ), .ZN(\add_98/n249 ) );
  XNOR2_X2 \add_98/U310  ( .A(\add_98/n247 ), .B(\add_98/n248 ), .ZN(N50) );
  INV_X4 \add_98/U309  ( .A(\add_98/n235 ), .ZN(\add_98/n244 ) );
  INV_X4 \add_98/U308  ( .A(\add_98/n243 ), .ZN(\add_98/n242 ) );
  NAND2_X2 \add_98/U307  ( .A1(\add_98/n202 ), .A2(\add_98/n201 ), .ZN(
        \add_98/n241 ) );
  INV_X4 \add_98/U306  ( .A(rnd_q[150]), .ZN(\add_98/n238 ) );
  INV_X4 \add_98/U305  ( .A(cv_q[150]), .ZN(\add_98/n239 ) );
  NAND2_X2 \add_98/U304  ( .A1(\add_98/n238 ), .A2(\add_98/n239 ), .ZN(
        \add_98/n198 ) );
  NAND2_X2 \add_98/U303  ( .A1(rnd_q[150]), .A2(cv_q[150]), .ZN(\add_98/n203 )
         );
  XNOR2_X2 \add_98/U302  ( .A(\add_98/n237 ), .B(\add_98/n31 ), .ZN(N51) );
  NAND2_X2 \add_98/U301  ( .A1(\add_98/n202 ), .A2(\add_98/n201 ), .ZN(
        \add_98/n236 ) );
  NAND2_X2 \add_98/U300  ( .A1(\add_98/n236 ), .A2(\add_98/n198 ), .ZN(
        \add_98/n233 ) );
  NAND2_X2 \add_98/U299  ( .A1(\add_98/n235 ), .A2(\add_98/n198 ), .ZN(
        \add_98/n228 ) );
  INV_X4 \add_98/U298  ( .A(rnd_q[151]), .ZN(\add_98/n231 ) );
  INV_X4 \add_98/U297  ( .A(cv_q[151]), .ZN(\add_98/n232 ) );
  NAND2_X2 \add_98/U296  ( .A1(\add_98/n231 ), .A2(\add_98/n232 ), .ZN(
        \add_98/n199 ) );
  NAND2_X2 \add_98/U295  ( .A1(rnd_q[151]), .A2(cv_q[151]), .ZN(\add_98/n151 )
         );
  NAND2_X2 \add_98/U294  ( .A1(\add_98/n199 ), .A2(\add_98/n151 ), .ZN(
        \add_98/n230 ) );
  XNOR2_X2 \add_98/U293  ( .A(\add_98/n229 ), .B(\add_98/n230 ), .ZN(N52) );
  INV_X4 \add_98/U292  ( .A(\add_98/n228 ), .ZN(\add_98/n227 ) );
  NAND2_X2 \add_98/U291  ( .A1(\add_98/n227 ), .A2(\add_98/n199 ), .ZN(
        \add_98/n146 ) );
  NAND2_X2 \add_98/U290  ( .A1(rnd_q[133]), .A2(cv_q[133]), .ZN(\add_98/n226 )
         );
  NAND2_X2 \add_98/U289  ( .A1(\add_98/n67 ), .A2(\add_98/n226 ), .ZN(
        \add_98/n225 ) );
  NAND2_X2 \add_98/U288  ( .A1(\add_98/n224 ), .A2(\add_98/n225 ), .ZN(
        \add_98/n223 ) );
  NAND2_X2 \add_98/U287  ( .A1(\add_98/n22 ), .A2(\add_98/n223 ), .ZN(
        \add_98/n221 ) );
  INV_X4 \add_98/U286  ( .A(\add_98/n214 ), .ZN(\add_98/n222 ) );
  NAND4_X2 \add_98/U285  ( .A1(\add_98/n221 ), .A2(\add_98/n3 ), .A3(
        \add_98/n313 ), .A4(\add_98/n222 ), .ZN(\add_98/n206 ) );
  NAND2_X2 \add_98/U284  ( .A1(rnd_q[129]), .A2(cv_q[129]), .ZN(\add_98/n219 )
         );
  NAND2_X2 \add_98/U283  ( .A1(\add_98/n219 ), .A2(\add_98/n220 ), .ZN(
        \add_98/n218 ) );
  NAND2_X2 \add_98/U282  ( .A1(\add_98/n1 ), .A2(\add_98/n218 ), .ZN(
        \add_98/n216 ) );
  NAND2_X2 \add_98/U281  ( .A1(\add_98/n204 ), .A2(\add_98/n205 ), .ZN(
        \add_98/n188 ) );
  INV_X4 \add_98/U280  ( .A(\add_98/n145 ), .ZN(\add_98/n197 ) );
  NAND2_X2 \add_98/U279  ( .A1(\add_98/n197 ), .A2(\add_98/n151 ), .ZN(
        \add_98/n190 ) );
  INV_X4 \add_98/U278  ( .A(\add_98/n196 ), .ZN(\add_98/n193 ) );
  INV_X4 \add_98/U277  ( .A(\add_98/n195 ), .ZN(\add_98/n194 ) );
  NAND2_X2 \add_98/U276  ( .A1(\add_98/n188 ), .A2(\add_98/n189 ), .ZN(
        \add_98/n162 ) );
  NAND2_X2 \add_98/U275  ( .A1(rnd_q[152]), .A2(cv_q[152]), .ZN(\add_98/n186 )
         );
  NAND2_X2 \add_98/U274  ( .A1(\add_98/n186 ), .A2(\add_98/n171 ), .ZN(
        \add_98/n187 ) );
  XNOR2_X2 \add_98/U273  ( .A(\add_98/n162 ), .B(\add_98/n187 ), .ZN(N53) );
  INV_X4 \add_98/U272  ( .A(\add_98/n180 ), .ZN(\add_98/n171 ) );
  NAND2_X2 \add_98/U271  ( .A1(\add_98/n171 ), .A2(\add_98/n162 ), .ZN(
        \add_98/n185 ) );
  NAND2_X2 \add_98/U270  ( .A1(\add_98/n185 ), .A2(\add_98/n186 ), .ZN(
        \add_98/n181 ) );
  NAND2_X2 \add_98/U269  ( .A1(rnd_q[153]), .A2(cv_q[153]), .ZN(\add_98/n160 )
         );
  INV_X4 \add_98/U268  ( .A(rnd_q[153]), .ZN(\add_98/n183 ) );
  INV_X4 \add_98/U267  ( .A(cv_q[153]), .ZN(\add_98/n184 ) );
  NAND2_X2 \add_98/U266  ( .A1(\add_98/n183 ), .A2(\add_98/n184 ), .ZN(
        \add_98/n170 ) );
  NAND2_X2 \add_98/U265  ( .A1(\add_98/n160 ), .A2(\add_98/n170 ), .ZN(
        \add_98/n182 ) );
  XNOR2_X2 \add_98/U264  ( .A(\add_98/n181 ), .B(\add_98/n182 ), .ZN(N54) );
  INV_X4 \add_98/U263  ( .A(\add_98/n162 ), .ZN(\add_98/n179 ) );
  INV_X4 \add_98/U262  ( .A(\add_98/n170 ), .ZN(\add_98/n177 ) );
  NAND2_X2 \add_98/U261  ( .A1(cv_q[152]), .A2(rnd_q[152]), .ZN(\add_98/n178 )
         );
  NAND2_X2 \add_98/U260  ( .A1(\add_98/n8 ), .A2(\add_98/n160 ), .ZN(
        \add_98/n176 ) );
  INV_X4 \add_98/U259  ( .A(rnd_q[154]), .ZN(\add_98/n173 ) );
  INV_X4 \add_98/U258  ( .A(cv_q[154]), .ZN(\add_98/n174 ) );
  NAND2_X2 \add_98/U257  ( .A1(\add_98/n173 ), .A2(\add_98/n174 ), .ZN(
        \add_98/n158 ) );
  NAND2_X2 \add_98/U256  ( .A1(rnd_q[154]), .A2(cv_q[154]), .ZN(\add_98/n161 )
         );
  XNOR2_X2 \add_98/U255  ( .A(\add_98/n172 ), .B(\add_98/n30 ), .ZN(N55) );
  NAND2_X2 \add_98/U254  ( .A1(\add_98/n36 ), .A2(\add_98/n162 ), .ZN(
        \add_98/n167 ) );
  NAND2_X2 \add_98/U253  ( .A1(\add_98/n169 ), .A2(\add_98/n158 ), .ZN(
        \add_98/n168 ) );
  NAND2_X2 \add_98/U252  ( .A1(\add_98/n167 ), .A2(\add_98/n168 ), .ZN(
        \add_98/n163 ) );
  INV_X4 \add_98/U251  ( .A(rnd_q[155]), .ZN(\add_98/n165 ) );
  INV_X4 \add_98/U250  ( .A(cv_q[155]), .ZN(\add_98/n166 ) );
  NAND2_X2 \add_98/U249  ( .A1(\add_98/n165 ), .A2(\add_98/n166 ), .ZN(
        \add_98/n149 ) );
  NAND2_X2 \add_98/U248  ( .A1(rnd_q[155]), .A2(cv_q[155]), .ZN(\add_98/n157 )
         );
  NAND2_X2 \add_98/U247  ( .A1(\add_98/n149 ), .A2(\add_98/n157 ), .ZN(
        \add_98/n164 ) );
  XNOR2_X2 \add_98/U246  ( .A(\add_98/n163 ), .B(\add_98/n164 ), .ZN(N56) );
  NAND2_X2 \add_98/U245  ( .A1(\add_98/n156 ), .A2(\add_98/n157 ), .ZN(
        \add_98/n152 ) );
  INV_X4 \add_98/U244  ( .A(rnd_q[156]), .ZN(\add_98/n154 ) );
  INV_X4 \add_98/U243  ( .A(cv_q[156]), .ZN(\add_98/n155 ) );
  NAND2_X2 \add_98/U242  ( .A1(\add_98/n154 ), .A2(\add_98/n155 ), .ZN(
        \add_98/n150 ) );
  NAND2_X2 \add_98/U241  ( .A1(rnd_q[156]), .A2(cv_q[156]), .ZN(\add_98/n102 )
         );
  XNOR2_X2 \add_98/U240  ( .A(\add_98/n153 ), .B(\add_98/n32 ), .ZN(N57) );
  INV_X4 \add_98/U239  ( .A(\add_98/n151 ), .ZN(\add_98/n148 ) );
  INV_X4 \add_98/U238  ( .A(\add_98/n121 ), .ZN(\add_98/n105 ) );
  INV_X4 \add_98/U237  ( .A(\add_98/n102 ), .ZN(\add_98/n147 ) );
  INV_X4 \add_98/U236  ( .A(\add_98/n146 ), .ZN(\add_98/n104 ) );
  INV_X4 \add_98/U235  ( .A(\add_98/n128 ), .ZN(\add_98/n88 ) );
  NAND2_X2 \add_98/U234  ( .A1(\add_98/n125 ), .A2(\add_98/n126 ), .ZN(
        \add_98/n103 ) );
  NAND2_X2 \add_98/U233  ( .A1(\add_98/n103 ), .A2(\add_98/n13 ), .ZN(
        \add_98/n144 ) );
  NAND2_X2 \add_98/U232  ( .A1(\add_98/n145 ), .A2(\add_98/n105 ), .ZN(
        \add_98/n94 ) );
  NAND4_X2 \add_98/U231  ( .A1(\add_98/n142 ), .A2(\add_98/n143 ), .A3(
        \add_98/n144 ), .A4(\add_98/n94 ), .ZN(\add_98/n138 ) );
  NAND2_X2 \add_98/U230  ( .A1(rnd_q[157]), .A2(cv_q[157]), .ZN(\add_98/n92 )
         );
  INV_X4 \add_98/U229  ( .A(rnd_q[157]), .ZN(\add_98/n140 ) );
  INV_X4 \add_98/U228  ( .A(cv_q[157]), .ZN(\add_98/n141 ) );
  NAND2_X2 \add_98/U227  ( .A1(\add_98/n140 ), .A2(\add_98/n141 ), .ZN(
        \add_98/n118 ) );
  NAND2_X2 \add_98/U226  ( .A1(\add_98/n92 ), .A2(\add_98/n118 ), .ZN(
        \add_98/n139 ) );
  XNOR2_X2 \add_98/U225  ( .A(\add_98/n138 ), .B(\add_98/n139 ), .ZN(N58) );
  XNOR2_X2 \add_98/U224  ( .A(\add_98/n81 ), .B(\add_98/n135 ), .ZN(N31) );
  INV_X4 \add_98/U223  ( .A(\add_98/n133 ), .ZN(\add_98/n129 ) );
  NAND2_X2 \add_98/U222  ( .A1(\add_98/n131 ), .A2(\add_98/n132 ), .ZN(
        \add_98/n130 ) );
  NAND2_X2 \add_98/U221  ( .A1(\add_98/n125 ), .A2(\add_98/n126 ), .ZN(
        \add_98/n124 ) );
  NAND2_X2 \add_98/U220  ( .A1(\add_98/n104 ), .A2(\add_98/n118 ), .ZN(
        \add_98/n122 ) );
  NAND2_X2 \add_98/U219  ( .A1(\add_98/n21 ), .A2(\add_98/n118 ), .ZN(
        \add_98/n114 ) );
  INV_X4 \add_98/U218  ( .A(\add_98/n94 ), .ZN(\add_98/n119 ) );
  NAND2_X2 \add_98/U217  ( .A1(\add_98/n119 ), .A2(\add_98/n118 ), .ZN(
        \add_98/n115 ) );
  INV_X4 \add_98/U216  ( .A(\add_98/n118 ), .ZN(\add_98/n106 ) );
  NAND2_X2 \add_98/U215  ( .A1(\add_98/n11 ), .A2(\add_98/n118 ), .ZN(
        \add_98/n117 ) );
  NAND4_X2 \add_98/U214  ( .A1(\add_98/n114 ), .A2(\add_98/n115 ), .A3(
        \add_98/n116 ), .A4(\add_98/n117 ), .ZN(\add_98/n113 ) );
  INV_X4 \add_98/U213  ( .A(rnd_q[158]), .ZN(\add_98/n110 ) );
  INV_X4 \add_98/U212  ( .A(cv_q[158]), .ZN(\add_98/n111 ) );
  NAND2_X2 \add_98/U211  ( .A1(rnd_q[158]), .A2(cv_q[158]), .ZN(\add_98/n101 )
         );
  INV_X4 \add_98/U210  ( .A(\add_98/n101 ), .ZN(\add_98/n109 ) );
  XNOR2_X2 \add_98/U209  ( .A(\add_98/n107 ), .B(\add_98/n108 ), .ZN(N59) );
  NAND2_X2 \add_98/U208  ( .A1(\add_98/n12 ), .A2(\add_98/n103 ), .ZN(
        \add_98/n84 ) );
  NAND2_X2 \add_98/U207  ( .A1(\add_98/n95 ), .A2(\add_98/n147 ), .ZN(
        \add_98/n100 ) );
  NAND2_X2 \add_98/U206  ( .A1(\add_98/n100 ), .A2(\add_98/n101 ), .ZN(
        \add_98/n96 ) );
  NAND2_X2 \add_98/U205  ( .A1(\add_98/n21 ), .A2(\add_98/n95 ), .ZN(
        \add_98/n98 ) );
  NAND2_X2 \add_98/U204  ( .A1(\add_98/n11 ), .A2(\add_98/n95 ), .ZN(
        \add_98/n99 ) );
  NAND2_X2 \add_98/U203  ( .A1(\add_98/n98 ), .A2(\add_98/n99 ), .ZN(
        \add_98/n97 ) );
  INV_X4 \add_98/U202  ( .A(\add_98/n95 ), .ZN(\add_98/n93 ) );
  NAND4_X2 \add_98/U201  ( .A1(\add_98/n84 ), .A2(\add_98/n85 ), .A3(
        \add_98/n86 ), .A4(\add_98/n87 ), .ZN(\add_98/n82 ) );
  XNOR2_X2 \add_98/U200  ( .A(rnd_q[159]), .B(cv_q[159]), .ZN(\add_98/n83 ) );
  XNOR2_X2 \add_98/U199  ( .A(\add_98/n82 ), .B(\add_98/n83 ), .ZN(N60) );
  XNOR2_X2 \add_98/U198  ( .A(\add_98/n75 ), .B(\add_98/n76 ), .ZN(N32) );
  INV_X4 \add_98/U197  ( .A(\add_98/n67 ), .ZN(\add_98/n73 ) );
  XNOR2_X2 \add_98/U196  ( .A(\add_98/n35 ), .B(\add_98/n74 ), .ZN(N33) );
  INV_X4 \add_98/U195  ( .A(\add_98/n64 ), .ZN(\add_98/n71 ) );
  XNOR2_X2 \add_98/U194  ( .A(\add_98/n69 ), .B(\add_98/n70 ), .ZN(N34) );
  NAND2_X2 \add_98/U193  ( .A1(rnd_q[134]), .A2(cv_q[134]), .ZN(\add_98/n59 )
         );
  NAND2_X2 \add_98/U192  ( .A1(\add_98/n59 ), .A2(\add_98/n5 ), .ZN(
        \add_98/n62 ) );
  NAND2_X2 \add_98/U191  ( .A1(\add_98/n35 ), .A2(\add_98/n67 ), .ZN(
        \add_98/n66 ) );
  NAND2_X2 \add_98/U190  ( .A1(\add_98/n65 ), .A2(\add_98/n66 ), .ZN(
        \add_98/n63 ) );
  NAND2_X2 \add_98/U189  ( .A1(\add_98/n63 ), .A2(\add_98/n64 ), .ZN(
        \add_98/n60 ) );
  XNOR2_X2 \add_98/U188  ( .A(\add_98/n62 ), .B(\add_98/n60 ), .ZN(N35) );
  NAND2_X2 \add_98/U187  ( .A1(\add_98/n60 ), .A2(\add_98/n5 ), .ZN(
        \add_98/n58 ) );
  NAND2_X2 \add_98/U186  ( .A1(\add_98/n58 ), .A2(\add_98/n59 ), .ZN(
        \add_98/n55 ) );
  NAND2_X2 \add_98/U185  ( .A1(\add_98/n57 ), .A2(\add_98/n3 ), .ZN(
        \add_98/n56 ) );
  XNOR2_X2 \add_98/U184  ( .A(\add_98/n55 ), .B(\add_98/n56 ), .ZN(N36) );
  INV_X4 \add_98/U183  ( .A(\add_98/n53 ), .ZN(\add_98/n46 ) );
  XNOR2_X2 \add_98/U182  ( .A(\add_98/n51 ), .B(\add_98/n52 ), .ZN(N37) );
  XNOR2_X2 \add_98/U181  ( .A(\add_98/n42 ), .B(\add_98/n43 ), .ZN(N38) );
  NAND2_X2 \add_98/U180  ( .A1(\add_98/n259 ), .A2(\add_98/n133 ), .ZN(
        \add_98/n258 ) );
  OR2_X2 \add_98/U179  ( .A1(cv_q[145]), .A2(rnd_q[145]), .ZN(\add_98/n41 ) );
  NOR2_X2 \add_98/U178  ( .A1(\add_98/n20 ), .A2(\add_98/n109 ), .ZN(
        \add_98/n108 ) );
  NOR2_X2 \add_98/U177  ( .A1(\add_98/n243 ), .A2(\add_98/n249 ), .ZN(
        \add_98/n248 ) );
  NOR2_X2 \add_98/U176  ( .A1(\add_98/n317 ), .A2(\add_98/n15 ), .ZN(
        \add_98/n319 ) );
  NOR2_X2 \add_98/U175  ( .A1(\add_98/n23 ), .A2(\add_98/n44 ), .ZN(
        \add_98/n43 ) );
  NOR2_X2 \add_98/U174  ( .A1(\add_98/n71 ), .A2(\add_98/n68 ), .ZN(
        \add_98/n70 ) );
  NOR2_X2 \add_98/U173  ( .A1(\add_98/n14 ), .A2(\add_98/n73 ), .ZN(
        \add_98/n74 ) );
  NOR2_X2 \add_98/U172  ( .A1(\add_98/n77 ), .A2(\add_98/n78 ), .ZN(
        \add_98/n76 ) );
  AND2_X2 \add_98/U171  ( .A1(cv_q[136]), .A2(rnd_q[136]), .ZN(\add_98/n353 )
         );
  NOR2_X2 \add_98/U170  ( .A1(\add_98/n24 ), .A2(\add_98/n251 ), .ZN(
        \add_98/n252 ) );
  NOR2_X2 \add_98/U169  ( .A1(\add_98/n47 ), .A2(\add_98/n46 ), .ZN(
        \add_98/n52 ) );
  NOR2_X2 \add_98/U168  ( .A1(\add_98/n26 ), .A2(\add_98/n80 ), .ZN(
        \add_98/n135 ) );
  NOR2_X2 \add_98/U167  ( .A1(\add_98/n261 ), .A2(\add_98/n136 ), .ZN(
        \add_98/n260 ) );
  NOR2_X2 \add_98/U166  ( .A1(cv_q[145]), .A2(rnd_q[145]), .ZN(\add_98/n278 )
         );
  NOR2_X2 \add_98/U165  ( .A1(\add_98/n278 ), .A2(\add_98/n279 ), .ZN(
        \add_98/n271 ) );
  NOR2_X2 \add_98/U164  ( .A1(cv_q[137]), .A2(rnd_q[137]), .ZN(\add_98/n355 )
         );
  NOR2_X2 \add_98/U163  ( .A1(cv_q[138]), .A2(rnd_q[138]), .ZN(\add_98/n356 )
         );
  NOR2_X2 \add_98/U162  ( .A1(\add_98/n355 ), .A2(\add_98/n356 ), .ZN(
        \add_98/n354 ) );
  NOR2_X2 \add_98/U161  ( .A1(cv_q[145]), .A2(rnd_q[145]), .ZN(\add_98/n281 )
         );
  NOR2_X2 \add_98/U160  ( .A1(\add_98/n308 ), .A2(\add_98/n312 ), .ZN(
        \add_98/n310 ) );
  NOR2_X2 \add_98/U159  ( .A1(cv_q[148]), .A2(rnd_q[148]), .ZN(\add_98/n246 )
         );
  NOR2_X2 \add_98/U158  ( .A1(cv_q[149]), .A2(rnd_q[149]), .ZN(\add_98/n245 )
         );
  NOR2_X2 \add_98/U157  ( .A1(\add_98/n245 ), .A2(\add_98/n246 ), .ZN(
        \add_98/n235 ) );
  NOR2_X2 \add_98/U156  ( .A1(cv_q[133]), .A2(rnd_q[133]), .ZN(\add_98/n295 )
         );
  NOR2_X2 \add_98/U155  ( .A1(cv_q[134]), .A2(rnd_q[134]), .ZN(\add_98/n296 )
         );
  NOR2_X2 \add_98/U154  ( .A1(\add_98/n295 ), .A2(\add_98/n296 ), .ZN(
        \add_98/n224 ) );
  NOR2_X2 \add_98/U153  ( .A1(cv_q[133]), .A2(rnd_q[133]), .ZN(\add_98/n388 )
         );
  NOR2_X2 \add_98/U152  ( .A1(\add_98/n343 ), .A2(\add_98/n318 ), .ZN(
        \add_98/n342 ) );
  NOR2_X2 \add_98/U151  ( .A1(cv_q[149]), .A2(rnd_q[149]), .ZN(\add_98/n243 )
         );
  OR2_X2 \add_98/U150  ( .A1(\add_98/n281 ), .A2(\add_98/n282 ), .ZN(
        \add_98/n40 ) );
  NAND3_X2 \add_98/U149  ( .A1(cv_q[148]), .A2(rnd_q[148]), .A3(\add_98/n242 ), 
        .ZN(\add_98/n202 ) );
  NOR2_X2 \add_98/U148  ( .A1(cv_q[130]), .A2(rnd_q[130]), .ZN(\add_98/n80 )
         );
  NOR2_X2 \add_98/U147  ( .A1(cv_q[131]), .A2(rnd_q[131]), .ZN(\add_98/n77 )
         );
  NOR2_X2 \add_98/U146  ( .A1(cv_q[129]), .A2(rnd_q[129]), .ZN(\add_98/n136 )
         );
  NOR2_X2 \add_98/U145  ( .A1(cv_q[148]), .A2(rnd_q[148]), .ZN(\add_98/n251 )
         );
  NOR2_X2 \add_98/U144  ( .A1(cv_q[144]), .A2(rnd_q[144]), .ZN(\add_98/n279 )
         );
  NOR2_X2 \add_98/U143  ( .A1(cv_q[134]), .A2(rnd_q[134]), .ZN(\add_98/n61 )
         );
  NOR2_X2 \add_98/U142  ( .A1(cv_q[152]), .A2(rnd_q[152]), .ZN(\add_98/n180 )
         );
  NOR2_X2 \add_98/U141  ( .A1(cv_q[133]), .A2(rnd_q[133]), .ZN(\add_98/n68 )
         );
  NOR2_X2 \add_98/U140  ( .A1(\add_98/n77 ), .A2(\add_98/n384 ), .ZN(
        \add_98/n217 ) );
  NOR2_X2 \add_98/U139  ( .A1(cv_q[142]), .A2(rnd_q[142]), .ZN(\add_98/n308 )
         );
  NOR3_X2 \add_98/U138  ( .A1(\add_98/n307 ), .A2(\add_98/n308 ), .A3(
        \add_98/n309 ), .ZN(\add_98/n306 ) );
  NOR2_X2 \add_98/U137  ( .A1(cv_q[138]), .A2(rnd_q[138]), .ZN(\add_98/n351 )
         );
  NOR2_X2 \add_98/U136  ( .A1(cv_q[136]), .A2(rnd_q[136]), .ZN(\add_98/n47 )
         );
  NOR2_X2 \add_98/U135  ( .A1(cv_q[137]), .A2(rnd_q[137]), .ZN(\add_98/n44 )
         );
  NOR2_X2 \add_98/U134  ( .A1(cv_q[140]), .A2(rnd_q[140]), .ZN(\add_98/n318 )
         );
  NOR2_X2 \add_98/U133  ( .A1(cv_q[141]), .A2(rnd_q[141]), .ZN(\add_98/n309 )
         );
  NOR2_X2 \add_98/U132  ( .A1(\add_98/n18 ), .A2(\add_98/n152 ), .ZN(
        \add_98/n153 ) );
  NOR2_X2 \add_98/U131  ( .A1(\add_98/n347 ), .A2(\add_98/n348 ), .ZN(
        \add_98/n346 ) );
  NAND3_X2 \add_98/U130  ( .A1(\add_98/n345 ), .A2(\add_98/n16 ), .A3(
        \add_98/n346 ), .ZN(\add_98/n315 ) );
  NOR2_X2 \add_98/U129  ( .A1(\add_98/n303 ), .A2(\add_98/n217 ), .ZN(
        \add_98/n301 ) );
  NAND3_X2 \add_98/U128  ( .A1(\add_98/n379 ), .A2(\add_98/n373 ), .A3(
        \add_98/n380 ), .ZN(\add_98/n371 ) );
  NOR2_X2 \add_98/U127  ( .A1(\add_98/n23 ), .A2(\add_98/n391 ), .ZN(
        \add_98/n370 ) );
  NAND3_X2 \add_98/U126  ( .A1(\add_98/n370 ), .A2(\add_98/n371 ), .A3(
        \add_98/n372 ), .ZN(\add_98/n368 ) );
  NOR2_X2 \add_98/U125  ( .A1(\add_98/n96 ), .A2(\add_98/n97 ), .ZN(
        \add_98/n85 ) );
  OR2_X4 \add_98/U124  ( .A1(\add_98/n106 ), .A2(\add_98/n102 ), .ZN(
        \add_98/n39 ) );
  AND2_X2 \add_98/U123  ( .A1(\add_98/n92 ), .A2(\add_98/n39 ), .ZN(
        \add_98/n116 ) );
  NAND3_X2 \add_98/U122  ( .A1(\add_98/n336 ), .A2(\add_98/n4 ), .A3(
        \add_98/n6 ), .ZN(\add_98/n335 ) );
  NAND3_X2 \add_98/U121  ( .A1(\add_98/n29 ), .A2(\add_98/n329 ), .A3(
        \add_98/n335 ), .ZN(\add_98/n333 ) );
  NOR2_X2 \add_98/U120  ( .A1(\add_98/n80 ), .A2(\add_98/n81 ), .ZN(
        \add_98/n79 ) );
  NOR2_X2 \add_98/U119  ( .A1(\add_98/n79 ), .A2(\add_98/n26 ), .ZN(
        \add_98/n75 ) );
  NOR2_X2 \add_98/U118  ( .A1(\add_98/n35 ), .A2(\add_98/n50 ), .ZN(
        \add_98/n49 ) );
  NOR2_X2 \add_98/U117  ( .A1(\add_98/n49 ), .A2(\add_98/n19 ), .ZN(
        \add_98/n48 ) );
  NOR2_X2 \add_98/U116  ( .A1(\add_98/n47 ), .A2(\add_98/n48 ), .ZN(
        \add_98/n45 ) );
  NOR2_X2 \add_98/U115  ( .A1(\add_98/n45 ), .A2(\add_98/n46 ), .ZN(
        \add_98/n42 ) );
  NOR2_X2 \add_98/U114  ( .A1(\add_98/n251 ), .A2(\add_98/n234 ), .ZN(
        \add_98/n250 ) );
  NOR2_X2 \add_98/U113  ( .A1(\add_98/n250 ), .A2(\add_98/n24 ), .ZN(
        \add_98/n247 ) );
  NOR2_X2 \add_98/U112  ( .A1(\add_98/n35 ), .A2(\add_98/n14 ), .ZN(
        \add_98/n72 ) );
  NOR2_X2 \add_98/U111  ( .A1(\add_98/n72 ), .A2(\add_98/n73 ), .ZN(
        \add_98/n69 ) );
  NOR3_X2 \add_98/U110  ( .A1(\add_98/n179 ), .A2(\add_98/n177 ), .A3(
        \add_98/n180 ), .ZN(\add_98/n175 ) );
  NOR2_X2 \add_98/U109  ( .A1(\add_98/n175 ), .A2(\add_98/n176 ), .ZN(
        \add_98/n172 ) );
  NOR2_X2 \add_98/U108  ( .A1(\add_98/n61 ), .A2(\add_98/n68 ), .ZN(
        \add_98/n376 ) );
  NAND3_X2 \add_98/U107  ( .A1(\add_98/n313 ), .A2(\add_98/n314 ), .A3(
        \add_98/n315 ), .ZN(\add_98/n132 ) );
  NOR2_X2 \add_98/U106  ( .A1(\add_98/n234 ), .A2(\add_98/n244 ), .ZN(
        \add_98/n240 ) );
  NOR2_X2 \add_98/U105  ( .A1(\add_98/n240 ), .A2(\add_98/n241 ), .ZN(
        \add_98/n237 ) );
  NOR3_X2 \add_98/U104  ( .A1(\add_98/n134 ), .A2(\add_98/n129 ), .A3(
        \add_98/n130 ), .ZN(\add_98/n127 ) );
  NOR2_X2 \add_98/U103  ( .A1(\add_98/n127 ), .A2(\add_98/n128 ), .ZN(
        \add_98/n123 ) );
  NOR2_X2 \add_98/U102  ( .A1(\add_98/n123 ), .A2(\add_98/n124 ), .ZN(
        \add_98/n120 ) );
  NAND3_X2 \add_98/U101  ( .A1(\add_98/n201 ), .A2(\add_98/n202 ), .A3(
        \add_98/n203 ), .ZN(\add_98/n200 ) );
  AND2_X4 \add_98/U100  ( .A1(\add_98/n198 ), .A2(\add_98/n199 ), .ZN(
        \add_98/n38 ) );
  AND2_X2 \add_98/U99  ( .A1(\add_98/n200 ), .A2(\add_98/n38 ), .ZN(
        \add_98/n145 ) );
  NOR2_X2 \add_98/U98  ( .A1(\add_98/n318 ), .A2(\add_98/n25 ), .ZN(
        \add_98/n324 ) );
  NOR2_X2 \add_98/U97  ( .A1(\add_98/n44 ), .A2(\add_98/n53 ), .ZN(
        \add_98/n391 ) );
  NOR2_X2 \add_98/U96  ( .A1(\add_98/n20 ), .A2(\add_98/n92 ), .ZN(
        \add_98/n91 ) );
  NOR2_X2 \add_98/U95  ( .A1(\add_98/n146 ), .A2(\add_98/n126 ), .ZN(
        \add_98/n192 ) );
  OR2_X4 \add_98/U94  ( .A1(\add_98/n136 ), .A2(\add_98/n220 ), .ZN(
        \add_98/n37 ) );
  AND2_X2 \add_98/U93  ( .A1(\add_98/n137 ), .A2(\add_98/n37 ), .ZN(
        \add_98/n81 ) );
  AND3_X2 \add_98/U92  ( .A1(\add_98/n170 ), .A2(\add_98/n158 ), .A3(
        \add_98/n171 ), .ZN(\add_98/n36 ) );
  NAND3_X2 \add_98/U91  ( .A1(\add_98/n149 ), .A2(\add_98/n150 ), .A3(
        \add_98/n36 ), .ZN(\add_98/n121 ) );
  NOR3_X2 \add_98/U90  ( .A1(\add_98/n193 ), .A2(\add_98/n146 ), .A3(
        \add_98/n194 ), .ZN(\add_98/n191 ) );
  NOR2_X2 \add_98/U89  ( .A1(\add_98/n318 ), .A2(\add_98/n25 ), .ZN(
        \add_98/n336 ) );
  NOR2_X2 \add_98/U88  ( .A1(\add_98/n47 ), .A2(\add_98/n44 ), .ZN(
        \add_98/n373 ) );
  NOR2_X2 \add_98/U87  ( .A1(\add_98/n14 ), .A2(\add_98/n68 ), .ZN(
        \add_98/n65 ) );
  NAND3_X2 \add_98/U86  ( .A1(\add_98/n215 ), .A2(\add_98/n216 ), .A3(
        \add_98/n382 ), .ZN(\add_98/n211 ) );
  AND3_X2 \add_98/U85  ( .A1(\add_98/n382 ), .A2(\add_98/n215 ), .A3(
        \add_98/n381 ), .ZN(\add_98/n35 ) );
  NAND3_X2 \add_98/U84  ( .A1(\add_98/n160 ), .A2(\add_98/n8 ), .A3(
        \add_98/n161 ), .ZN(\add_98/n159 ) );
  NAND3_X2 \add_98/U83  ( .A1(\add_98/n158 ), .A2(\add_98/n149 ), .A3(
        \add_98/n159 ), .ZN(\add_98/n156 ) );
  NOR2_X2 \add_98/U82  ( .A1(\add_98/n14 ), .A2(\add_98/n388 ), .ZN(
        \add_98/n387 ) );
  NAND3_X2 \add_98/U81  ( .A1(\add_98/n3 ), .A2(\add_98/n5 ), .A3(
        \add_98/n387 ), .ZN(\add_98/n50 ) );
  NOR3_X2 \add_98/U80  ( .A1(\add_98/n120 ), .A2(\add_98/n121 ), .A3(
        \add_98/n122 ), .ZN(\add_98/n112 ) );
  NOR2_X2 \add_98/U79  ( .A1(\add_98/n112 ), .A2(\add_98/n113 ), .ZN(
        \add_98/n107 ) );
  NOR2_X2 \add_98/U78  ( .A1(\add_98/n20 ), .A2(\add_98/n106 ), .ZN(
        \add_98/n95 ) );
  NOR2_X2 \add_98/U77  ( .A1(\add_98/n209 ), .A2(\add_98/n210 ), .ZN(
        \add_98/n208 ) );
  NAND3_X2 \add_98/U76  ( .A1(\add_98/n211 ), .A2(\add_98/n212 ), .A3(
        \add_98/n379 ), .ZN(\add_98/n207 ) );
  NAND3_X2 \add_98/U75  ( .A1(\add_98/n207 ), .A2(\add_98/n208 ), .A3(
        \add_98/n206 ), .ZN(\add_98/n205 ) );
  NAND3_X2 \add_98/U74  ( .A1(\add_98/n233 ), .A2(\add_98/n203 ), .A3(
        \add_98/n17 ), .ZN(\add_98/n229 ) );
  NOR2_X2 \add_98/U73  ( .A1(\add_98/n213 ), .A2(\add_98/n214 ), .ZN(
        \add_98/n291 ) );
  NAND3_X2 \add_98/U72  ( .A1(\add_98/n161 ), .A2(\add_98/n8 ), .A3(
        \add_98/n160 ), .ZN(\add_98/n169 ) );
  NOR3_X2 \add_98/U71  ( .A1(\add_98/n258 ), .A2(\add_98/n210 ), .A3(
        \add_98/n209 ), .ZN(\add_98/n255 ) );
  NOR2_X2 \add_98/U70  ( .A1(\add_98/n255 ), .A2(\add_98/n128 ), .ZN(
        \add_98/n253 ) );
  NOR2_X2 \add_98/U69  ( .A1(\add_98/n253 ), .A2(\add_98/n254 ), .ZN(
        \add_98/n234 ) );
  NOR3_X2 \add_98/U68  ( .A1(\add_98/n217 ), .A2(\add_98/n78 ), .A3(
        \add_98/n1 ), .ZN(\add_98/n300 ) );
  NOR2_X2 \add_98/U67  ( .A1(\add_98/n317 ), .A2(\add_98/n318 ), .ZN(
        \add_98/n316 ) );
  NAND3_X2 \add_98/U66  ( .A1(\add_98/n4 ), .A2(\add_98/n9 ), .A3(
        \add_98/n316 ), .ZN(\add_98/n213 ) );
  OR3_X4 \add_98/U65  ( .A1(\add_98/n310 ), .A2(\add_98/n311 ), .A3(
        \add_98/n15 ), .ZN(\add_98/n34 ) );
  OR2_X2 \add_98/U64  ( .A1(\add_98/n34 ), .A2(\add_98/n306 ), .ZN(
        \add_98/n304 ) );
  NOR2_X2 \add_98/U63  ( .A1(\add_98/n351 ), .A2(\add_98/n361 ), .ZN(
        \add_98/n360 ) );
  NAND3_X2 \add_98/U62  ( .A1(\add_98/n358 ), .A2(\add_98/n359 ), .A3(
        \add_98/n360 ), .ZN(\add_98/n214 ) );
  NOR3_X2 \add_98/U61  ( .A1(\add_98/n190 ), .A2(\add_98/n191 ), .A3(
        \add_98/n192 ), .ZN(\add_98/n189 ) );
  NOR2_X2 \add_98/U60  ( .A1(\add_98/n270 ), .A2(\add_98/n257 ), .ZN(
        \add_98/n265 ) );
  NOR2_X2 \add_98/U59  ( .A1(\add_98/n265 ), .A2(\add_98/n196 ), .ZN(
        \add_98/n262 ) );
  NOR2_X2 \add_98/U58  ( .A1(\add_98/n35 ), .A2(\add_98/n50 ), .ZN(
        \add_98/n54 ) );
  NOR2_X2 \add_98/U57  ( .A1(\add_98/n54 ), .A2(\add_98/n19 ), .ZN(
        \add_98/n51 ) );
  NOR2_X2 \add_98/U56  ( .A1(\add_98/n128 ), .A2(\add_98/n146 ), .ZN(
        \add_98/n204 ) );
  NOR2_X2 \add_98/U55  ( .A1(\add_98/n35 ), .A2(\add_98/n50 ), .ZN(
        \add_98/n362 ) );
  NOR2_X2 \add_98/U54  ( .A1(\add_98/n362 ), .A2(\add_98/n19 ), .ZN(
        \add_98/n357 ) );
  NOR2_X2 \add_98/U53  ( .A1(\add_98/n357 ), .A2(\add_98/n214 ), .ZN(
        \add_98/n344 ) );
  NOR2_X2 \add_98/U52  ( .A1(\add_98/n344 ), .A2(\add_98/n327 ), .ZN(
        \add_98/n341 ) );
  NOR2_X2 \add_98/U51  ( .A1(\add_98/n93 ), .A2(\add_98/n94 ), .ZN(
        \add_98/n90 ) );
  NOR2_X2 \add_98/U50  ( .A1(\add_98/n213 ), .A2(\add_98/n214 ), .ZN(
        \add_98/n212 ) );
  NOR2_X2 \add_98/U49  ( .A1(\add_98/n324 ), .A2(\add_98/n325 ), .ZN(
        \add_98/n323 ) );
  NOR3_X2 \add_98/U48  ( .A1(\add_98/n322 ), .A2(\add_98/n323 ), .A3(
        \add_98/n27 ), .ZN(\add_98/n321 ) );
  NOR2_X2 \add_98/U47  ( .A1(\add_98/n311 ), .A2(\add_98/n321 ), .ZN(
        \add_98/n320 ) );
  NOR2_X2 \add_98/U46  ( .A1(\add_98/n35 ), .A2(\add_98/n50 ), .ZN(
        \add_98/n326 ) );
  NAND3_X2 \add_98/U45  ( .A1(\add_98/n89 ), .A2(\add_98/n13 ), .A3(
        \add_98/n88 ), .ZN(\add_98/n143 ) );
  NOR3_X2 \add_98/U44  ( .A1(\add_98/n11 ), .A2(\add_98/n21 ), .A3(
        \add_98/n147 ), .ZN(\add_98/n142 ) );
  NAND3_X2 \add_98/U43  ( .A1(\add_98/n88 ), .A2(\add_98/n89 ), .A3(
        \add_98/n12 ), .ZN(\add_98/n87 ) );
  NOR2_X2 \add_98/U42  ( .A1(\add_98/n90 ), .A2(\add_98/n91 ), .ZN(
        \add_98/n86 ) );
  NOR4_X2 \add_98/U41  ( .A1(\add_98/n326 ), .A2(\add_98/n327 ), .A3(
        \add_98/n19 ), .A4(\add_98/n325 ), .ZN(\add_98/n322 ) );
  NOR2_X2 \add_98/U40  ( .A1(\add_98/n261 ), .A2(\add_98/n78 ), .ZN(
        \add_98/n302 ) );
  NOR2_X2 \add_98/U39  ( .A1(\add_98/n50 ), .A2(\add_98/n300 ), .ZN(
        \add_98/n299 ) );
  NOR2_X2 \add_98/U38  ( .A1(\add_98/n213 ), .A2(\add_98/n214 ), .ZN(
        \add_98/n297 ) );
  NAND3_X2 \add_98/U37  ( .A1(\add_98/n297 ), .A2(\add_98/n298 ), .A3(
        \add_98/n299 ), .ZN(\add_98/n133 ) );
  NOR2_X2 \add_98/U36  ( .A1(\add_98/n210 ), .A2(\add_98/n209 ), .ZN(
        \add_98/n289 ) );
  NAND3_X2 \add_98/U35  ( .A1(\add_98/n289 ), .A2(\add_98/n133 ), .A3(
        \add_98/n259 ), .ZN(\add_98/n89 ) );
  AND2_X4 \add_98/U34  ( .A1(\add_98/n383 ), .A2(\add_98/n220 ), .ZN(N29) );
  AND2_X4 \add_98/U33  ( .A1(\add_98/n150 ), .A2(\add_98/n102 ), .ZN(
        \add_98/n32 ) );
  AND2_X4 \add_98/U32  ( .A1(\add_98/n198 ), .A2(\add_98/n203 ), .ZN(
        \add_98/n31 ) );
  AND2_X4 \add_98/U31  ( .A1(\add_98/n158 ), .A2(\add_98/n161 ), .ZN(
        \add_98/n30 ) );
  OR2_X4 \add_98/U30  ( .A1(\add_98/n309 ), .A2(\add_98/n328 ), .ZN(
        \add_98/n29 ) );
  AND2_X4 \add_98/U29  ( .A1(\add_98/n126 ), .A2(\add_98/n195 ), .ZN(
        \add_98/n28 ) );
  OR2_X4 \add_98/U28  ( .A1(\add_98/n308 ), .A2(\add_98/n309 ), .ZN(
        \add_98/n27 ) );
  AND2_X4 \add_98/U27  ( .A1(rnd_q[130]), .A2(cv_q[130]), .ZN(\add_98/n26 ) );
  AND2_X4 \add_98/U26  ( .A1(\add_98/n214 ), .A2(\add_98/n340 ), .ZN(
        \add_98/n25 ) );
  AND2_X4 \add_98/U25  ( .A1(rnd_q[148]), .A2(cv_q[148]), .ZN(\add_98/n24 ) );
  AND2_X4 \add_98/U24  ( .A1(rnd_q[137]), .A2(cv_q[137]), .ZN(\add_98/n23 ) );
  AND2_X4 \add_98/U23  ( .A1(\add_98/n57 ), .A2(\add_98/n378 ), .ZN(
        \add_98/n22 ) );
  AND2_X4 \add_98/U22  ( .A1(\add_98/n148 ), .A2(\add_98/n105 ), .ZN(
        \add_98/n21 ) );
  AND2_X4 \add_98/U21  ( .A1(\add_98/n110 ), .A2(\add_98/n111 ), .ZN(
        \add_98/n20 ) );
  AND2_X4 \add_98/U20  ( .A1(\add_98/n374 ), .A2(\add_98/n3 ), .ZN(
        \add_98/n19 ) );
  AND3_X4 \add_98/U19  ( .A1(\add_98/n36 ), .A2(\add_98/n149 ), .A3(
        \add_98/n162 ), .ZN(\add_98/n18 ) );
  OR2_X4 \add_98/U18  ( .A1(\add_98/n234 ), .A2(\add_98/n228 ), .ZN(
        \add_98/n17 ) );
  OR2_X4 \add_98/U17  ( .A1(\add_98/n351 ), .A2(\add_98/n352 ), .ZN(
        \add_98/n16 ) );
  AND2_X4 \add_98/U16  ( .A1(rnd_q[143]), .A2(cv_q[143]), .ZN(\add_98/n15 ) );
  AND2_X4 \add_98/U15  ( .A1(\add_98/n389 ), .A2(\add_98/n390 ), .ZN(
        \add_98/n14 ) );
  AND2_X4 \add_98/U14  ( .A1(\add_98/n104 ), .A2(\add_98/n105 ), .ZN(
        \add_98/n13 ) );
  AND3_X4 \add_98/U13  ( .A1(\add_98/n104 ), .A2(\add_98/n95 ), .A3(
        \add_98/n105 ), .ZN(\add_98/n12 ) );
  AND2_X4 \add_98/U12  ( .A1(\add_98/n152 ), .A2(\add_98/n150 ), .ZN(
        \add_98/n11 ) );
  OR2_X4 \add_98/U11  ( .A1(cv_q[130]), .A2(rnd_q[130]), .ZN(\add_98/n10 ) );
  OR2_X4 \add_98/U10  ( .A1(cv_q[142]), .A2(rnd_q[142]), .ZN(\add_98/n9 ) );
  OR2_X4 \add_98/U9  ( .A1(\add_98/n177 ), .A2(\add_98/n178 ), .ZN(\add_98/n8 ) );
  OR2_X4 \add_98/U8  ( .A1(cv_q[131]), .A2(rnd_q[131]), .ZN(\add_98/n7 ) );
  OR3_X4 \add_98/U7  ( .A1(\add_98/n326 ), .A2(\add_98/n19 ), .A3(
        \add_98/n327 ), .ZN(\add_98/n6 ) );
  OR2_X4 \add_98/U6  ( .A1(cv_q[134]), .A2(rnd_q[134]), .ZN(\add_98/n5 ) );
  OR2_X4 \add_98/U5  ( .A1(cv_q[141]), .A2(rnd_q[141]), .ZN(\add_98/n4 ) );
  OR2_X4 \add_98/U4  ( .A1(cv_q[135]), .A2(rnd_q[135]), .ZN(\add_98/n3 ) );
  OR2_X4 \add_98/U3  ( .A1(cv_q[129]), .A2(rnd_q[129]), .ZN(\add_98/n2 ) );
  AND3_X4 \add_98/U2  ( .A1(\add_98/n10 ), .A2(\add_98/n7 ), .A3(\add_98/n2 ), 
        .ZN(\add_98/n1 ) );
  NAND2_X2 \add_98_4/U421  ( .A1(rnd_q[32]), .A2(cv_q[32]), .ZN(
        \add_98_4/n221 ) );
  INV_X4 \add_98_4/U420  ( .A(\add_98_4/n352 ), .ZN(\add_98_4/n389 ) );
  NAND2_X2 \add_98_4/U419  ( .A1(rnd_q[42]), .A2(cv_q[42]), .ZN(
        \add_98_4/n351 ) );
  NAND2_X2 \add_98_4/U418  ( .A1(\add_98_4/n389 ), .A2(\add_98_4/n351 ), .ZN(
        \add_98_4/n368 ) );
  NAND2_X2 \add_98_4/U417  ( .A1(rnd_q[40]), .A2(cv_q[40]), .ZN(\add_98_4/n52 ) );
  INV_X4 \add_98_4/U416  ( .A(\add_98_4/n49 ), .ZN(\add_98_4/n378 ) );
  NAND2_X2 \add_98_4/U415  ( .A1(rnd_q[33]), .A2(cv_q[33]), .ZN(
        \add_98_4/n385 ) );
  NAND2_X2 \add_98_4/U414  ( .A1(\add_98_4/n385 ), .A2(\add_98_4/n221 ), .ZN(
        \add_98_4/n384 ) );
  NAND2_X2 \add_98_4/U413  ( .A1(\add_98_4/n1 ), .A2(\add_98_4/n384 ), .ZN(
        \add_98_4/n380 ) );
  NAND2_X2 \add_98_4/U412  ( .A1(cv_q[34]), .A2(rnd_q[34]), .ZN(
        \add_98_4/n383 ) );
  INV_X4 \add_98_4/U411  ( .A(\add_98_4/n218 ), .ZN(\add_98_4/n381 ) );
  NAND2_X2 \add_98_4/U410  ( .A1(rnd_q[35]), .A2(cv_q[35]), .ZN(
        \add_98_4/n216 ) );
  INV_X4 \add_98_4/U409  ( .A(\add_98_4/n30 ), .ZN(\add_98_4/n379 ) );
  NAND2_X2 \add_98_4/U408  ( .A1(rnd_q[39]), .A2(cv_q[39]), .ZN(\add_98_4/n56 ) );
  NAND2_X2 \add_98_4/U407  ( .A1(rnd_q[38]), .A2(cv_q[38]), .ZN(
        \add_98_4/n377 ) );
  NAND2_X2 \add_98_4/U406  ( .A1(rnd_q[36]), .A2(cv_q[36]), .ZN(\add_98_4/n66 ) );
  NAND2_X2 \add_98_4/U405  ( .A1(rnd_q[37]), .A2(cv_q[37]), .ZN(\add_98_4/n63 ) );
  NAND2_X2 \add_98_4/U404  ( .A1(\add_98_4/n66 ), .A2(\add_98_4/n63 ), .ZN(
        \add_98_4/n376 ) );
  NAND2_X2 \add_98_4/U403  ( .A1(\add_98_4/n375 ), .A2(\add_98_4/n376 ), .ZN(
        \add_98_4/n374 ) );
  NAND2_X2 \add_98_4/U402  ( .A1(\add_98_4/n35 ), .A2(\add_98_4/n374 ), .ZN(
        \add_98_4/n373 ) );
  NAND2_X2 \add_98_4/U401  ( .A1(\add_98_4/n19 ), .A2(\add_98_4/n372 ), .ZN(
        \add_98_4/n371 ) );
  XNOR2_X2 \add_98_4/U400  ( .A(\add_98_4/n368 ), .B(\add_98_4/n367 ), .ZN(
        N135) );
  NAND2_X2 \add_98_4/U399  ( .A1(\add_98_4/n367 ), .A2(\add_98_4/n389 ), .ZN(
        \add_98_4/n366 ) );
  NAND2_X2 \add_98_4/U398  ( .A1(\add_98_4/n366 ), .A2(\add_98_4/n351 ), .ZN(
        \add_98_4/n364 ) );
  NAND2_X2 \add_98_4/U397  ( .A1(rnd_q[43]), .A2(cv_q[43]), .ZN(
        \add_98_4/n350 ) );
  NAND2_X2 \add_98_4/U396  ( .A1(\add_98_4/n350 ), .A2(\add_98_4/n315 ), .ZN(
        \add_98_4/n365 ) );
  XNOR2_X2 \add_98_4/U395  ( .A(\add_98_4/n364 ), .B(\add_98_4/n365 ), .ZN(
        N136) );
  INV_X4 \add_98_4/U394  ( .A(\add_98_4/n43 ), .ZN(\add_98_4/n359 ) );
  INV_X4 \add_98_4/U393  ( .A(\add_98_4/n46 ), .ZN(\add_98_4/n360 ) );
  INV_X4 \add_98_4/U392  ( .A(\add_98_4/n315 ), .ZN(\add_98_4/n362 ) );
  NAND2_X2 \add_98_4/U391  ( .A1(\add_98_4/n354 ), .A2(\add_98_4/n355 ), .ZN(
        \add_98_4/n346 ) );
  NAND2_X2 \add_98_4/U390  ( .A1(cv_q[41]), .A2(rnd_q[41]), .ZN(
        \add_98_4/n353 ) );
  INV_X4 \add_98_4/U389  ( .A(\add_98_4/n351 ), .ZN(\add_98_4/n348 ) );
  INV_X4 \add_98_4/U388  ( .A(\add_98_4/n350 ), .ZN(\add_98_4/n349 ) );
  NAND2_X2 \add_98_4/U387  ( .A1(\add_98_4/n316 ), .A2(\add_98_4/n315 ), .ZN(
        \add_98_4/n341 ) );
  INV_X4 \add_98_4/U386  ( .A(\add_98_4/n341 ), .ZN(\add_98_4/n328 ) );
  NAND2_X2 \add_98_4/U385  ( .A1(rnd_q[44]), .A2(cv_q[44]), .ZN(
        \add_98_4/n329 ) );
  INV_X4 \add_98_4/U384  ( .A(\add_98_4/n329 ), .ZN(\add_98_4/n344 ) );
  XNOR2_X2 \add_98_4/U383  ( .A(\add_98_4/n342 ), .B(\add_98_4/n343 ), .ZN(
        N137) );
  NAND2_X2 \add_98_4/U382  ( .A1(\add_98_4/n337 ), .A2(\add_98_4/n7 ), .ZN(
        \add_98_4/n340 ) );
  NAND2_X2 \add_98_4/U381  ( .A1(\add_98_4/n340 ), .A2(\add_98_4/n329 ), .ZN(
        \add_98_4/n338 ) );
  NAND2_X2 \add_98_4/U380  ( .A1(rnd_q[45]), .A2(cv_q[45]), .ZN(
        \add_98_4/n330 ) );
  NAND2_X2 \add_98_4/U379  ( .A1(\add_98_4/n330 ), .A2(\add_98_4/n4 ), .ZN(
        \add_98_4/n339 ) );
  XNOR2_X2 \add_98_4/U378  ( .A(\add_98_4/n338 ), .B(\add_98_4/n339 ), .ZN(
        N138) );
  NAND2_X2 \add_98_4/U377  ( .A1(rnd_q[46]), .A2(cv_q[46]), .ZN(
        \add_98_4/n331 ) );
  NAND2_X2 \add_98_4/U376  ( .A1(\add_98_4/n10 ), .A2(\add_98_4/n331 ), .ZN(
        \add_98_4/n335 ) );
  XNOR2_X2 \add_98_4/U375  ( .A(\add_98_4/n334 ), .B(\add_98_4/n335 ), .ZN(
        N139) );
  INV_X4 \add_98_4/U374  ( .A(rnd_q[47]), .ZN(\add_98_4/n332 ) );
  INV_X4 \add_98_4/U373  ( .A(cv_q[47]), .ZN(\add_98_4/n333 ) );
  NAND2_X2 \add_98_4/U372  ( .A1(\add_98_4/n332 ), .A2(\add_98_4/n333 ), .ZN(
        \add_98_4/n306 ) );
  INV_X4 \add_98_4/U371  ( .A(\add_98_4/n306 ), .ZN(\add_98_4/n318 ) );
  INV_X4 \add_98_4/U370  ( .A(\add_98_4/n331 ), .ZN(\add_98_4/n312 ) );
  NAND2_X2 \add_98_4/U369  ( .A1(\add_98_4/n329 ), .A2(\add_98_4/n330 ), .ZN(
        \add_98_4/n326 ) );
  XNOR2_X2 \add_98_4/U368  ( .A(\add_98_4/n320 ), .B(\add_98_4/n321 ), .ZN(
        N140) );
  NAND2_X2 \add_98_4/U367  ( .A1(rnd_q[48]), .A2(cv_q[48]), .ZN(
        \add_98_4/n287 ) );
  NAND2_X2 \add_98_4/U366  ( .A1(\add_98_4/n287 ), .A2(\add_98_4/n289 ), .ZN(
        \add_98_4/n290 ) );
  INV_X4 \add_98_4/U365  ( .A(\add_98_4/n214 ), .ZN(\add_98_4/n314 ) );
  INV_X4 \add_98_4/U364  ( .A(\add_98_4/n133 ), .ZN(\add_98_4/n211 ) );
  NAND2_X2 \add_98_4/U363  ( .A1(cv_q[45]), .A2(rnd_q[45]), .ZN(
        \add_98_4/n313 ) );
  NAND2_X2 \add_98_4/U362  ( .A1(rnd_q[44]), .A2(cv_q[44]), .ZN(
        \add_98_4/n308 ) );
  NAND2_X2 \add_98_4/U361  ( .A1(\add_98_4/n305 ), .A2(\add_98_4/n306 ), .ZN(
        \add_98_4/n132 ) );
  INV_X4 \add_98_4/U360  ( .A(\add_98_4/n132 ), .ZN(\add_98_4/n210 ) );
  NAND2_X2 \add_98_4/U359  ( .A1(rnd_q[33]), .A2(cv_q[33]), .ZN(
        \add_98_4/n138 ) );
  INV_X4 \add_98_4/U358  ( .A(\add_98_4/n138 ), .ZN(\add_98_4/n262 ) );
  INV_X4 \add_98_4/U357  ( .A(\add_98_4/n216 ), .ZN(\add_98_4/n77 ) );
  NAND2_X2 \add_98_4/U356  ( .A1(\add_98_4/n303 ), .A2(\add_98_4/n304 ), .ZN(
        \add_98_4/n300 ) );
  NAND2_X2 \add_98_4/U355  ( .A1(rnd_q[37]), .A2(cv_q[37]), .ZN(
        \add_98_4/n296 ) );
  NAND2_X2 \add_98_4/U354  ( .A1(\add_98_4/n66 ), .A2(\add_98_4/n296 ), .ZN(
        \add_98_4/n295 ) );
  NAND2_X2 \add_98_4/U353  ( .A1(\add_98_4/n225 ), .A2(\add_98_4/n295 ), .ZN(
        \add_98_4/n294 ) );
  NAND2_X2 \add_98_4/U352  ( .A1(\add_98_4/n35 ), .A2(\add_98_4/n294 ), .ZN(
        \add_98_4/n292 ) );
  NAND3_X2 \add_98_4/U351  ( .A1(\add_98_4/n292 ), .A2(\add_98_4/n3 ), .A3(
        \add_98_4/n293 ), .ZN(\add_98_4/n260 ) );
  INV_X4 \add_98_4/U350  ( .A(\add_98_4/n260 ), .ZN(\add_98_4/n135 ) );
  XNOR2_X2 \add_98_4/U349  ( .A(\add_98_4/n290 ), .B(\add_98_4/n88 ), .ZN(N141) );
  INV_X4 \add_98_4/U348  ( .A(\add_98_4/n281 ), .ZN(\add_98_4/n289 ) );
  NAND2_X2 \add_98_4/U347  ( .A1(\add_98_4/n88 ), .A2(\add_98_4/n289 ), .ZN(
        \add_98_4/n288 ) );
  NAND2_X2 \add_98_4/U346  ( .A1(\add_98_4/n287 ), .A2(\add_98_4/n288 ), .ZN(
        \add_98_4/n285 ) );
  NAND2_X2 \add_98_4/U345  ( .A1(rnd_q[49]), .A2(cv_q[49]), .ZN(
        \add_98_4/n282 ) );
  NAND2_X2 \add_98_4/U344  ( .A1(\add_98_4/n37 ), .A2(\add_98_4/n282 ), .ZN(
        \add_98_4/n286 ) );
  XNOR2_X2 \add_98_4/U343  ( .A(\add_98_4/n285 ), .B(\add_98_4/n286 ), .ZN(
        N142) );
  NAND2_X2 \add_98_4/U342  ( .A1(cv_q[48]), .A2(rnd_q[48]), .ZN(
        \add_98_4/n284 ) );
  NAND2_X2 \add_98_4/U341  ( .A1(\add_98_4/n34 ), .A2(\add_98_4/n282 ), .ZN(
        \add_98_4/n270 ) );
  INV_X4 \add_98_4/U340  ( .A(\add_98_4/n270 ), .ZN(\add_98_4/n278 ) );
  NAND2_X2 \add_98_4/U339  ( .A1(\add_98_4/n273 ), .A2(\add_98_4/n88 ), .ZN(
        \add_98_4/n279 ) );
  NAND2_X2 \add_98_4/U338  ( .A1(\add_98_4/n278 ), .A2(\add_98_4/n279 ), .ZN(
        \add_98_4/n274 ) );
  NAND2_X2 \add_98_4/U337  ( .A1(rnd_q[50]), .A2(cv_q[50]), .ZN(
        \add_98_4/n269 ) );
  INV_X4 \add_98_4/U336  ( .A(rnd_q[50]), .ZN(\add_98_4/n276 ) );
  INV_X4 \add_98_4/U335  ( .A(cv_q[50]), .ZN(\add_98_4/n277 ) );
  NAND2_X2 \add_98_4/U334  ( .A1(\add_98_4/n276 ), .A2(\add_98_4/n277 ), .ZN(
        \add_98_4/n271 ) );
  NAND2_X2 \add_98_4/U333  ( .A1(\add_98_4/n269 ), .A2(\add_98_4/n271 ), .ZN(
        \add_98_4/n275 ) );
  XNOR2_X2 \add_98_4/U332  ( .A(\add_98_4/n274 ), .B(\add_98_4/n275 ), .ZN(
        N143) );
  INV_X4 \add_98_4/U331  ( .A(\add_98_4/n88 ), .ZN(\add_98_4/n272 ) );
  NAND2_X2 \add_98_4/U330  ( .A1(\add_98_4/n273 ), .A2(\add_98_4/n271 ), .ZN(
        \add_98_4/n258 ) );
  NAND2_X2 \add_98_4/U329  ( .A1(\add_98_4/n270 ), .A2(\add_98_4/n271 ), .ZN(
        \add_98_4/n268 ) );
  NAND2_X2 \add_98_4/U328  ( .A1(\add_98_4/n268 ), .A2(\add_98_4/n269 ), .ZN(
        \add_98_4/n197 ) );
  NAND2_X2 \add_98_4/U327  ( .A1(rnd_q[51]), .A2(cv_q[51]), .ZN(
        \add_98_4/n127 ) );
  INV_X4 \add_98_4/U326  ( .A(rnd_q[51]), .ZN(\add_98_4/n265 ) );
  INV_X4 \add_98_4/U325  ( .A(cv_q[51]), .ZN(\add_98_4/n266 ) );
  NAND2_X2 \add_98_4/U324  ( .A1(\add_98_4/n265 ), .A2(\add_98_4/n266 ), .ZN(
        \add_98_4/n196 ) );
  XNOR2_X2 \add_98_4/U323  ( .A(\add_98_4/n264 ), .B(\add_98_4/n23 ), .ZN(N144) );
  INV_X4 \add_98_4/U322  ( .A(\add_98_4/n221 ), .ZN(\add_98_4/n263 ) );
  XNOR2_X2 \add_98_4/U321  ( .A(\add_98_4/n221 ), .B(\add_98_4/n261 ), .ZN(
        N126) );
  INV_X4 \add_98_4/U320  ( .A(\add_98_4/n258 ), .ZN(\add_98_4/n257 ) );
  NAND2_X2 \add_98_4/U319  ( .A1(\add_98_4/n257 ), .A2(\add_98_4/n196 ), .ZN(
        \add_98_4/n129 ) );
  NAND2_X2 \add_98_4/U318  ( .A1(\add_98_4/n197 ), .A2(\add_98_4/n196 ), .ZN(
        \add_98_4/n126 ) );
  NAND2_X2 \add_98_4/U317  ( .A1(\add_98_4/n126 ), .A2(\add_98_4/n127 ), .ZN(
        \add_98_4/n255 ) );
  XNOR2_X2 \add_98_4/U316  ( .A(\add_98_4/n235 ), .B(\add_98_4/n253 ), .ZN(
        N145) );
  NAND2_X2 \add_98_4/U315  ( .A1(rnd_q[53]), .A2(cv_q[53]), .ZN(
        \add_98_4/n202 ) );
  INV_X4 \add_98_4/U314  ( .A(\add_98_4/n202 ), .ZN(\add_98_4/n250 ) );
  XNOR2_X2 \add_98_4/U313  ( .A(\add_98_4/n248 ), .B(\add_98_4/n249 ), .ZN(
        N146) );
  INV_X4 \add_98_4/U312  ( .A(\add_98_4/n236 ), .ZN(\add_98_4/n245 ) );
  INV_X4 \add_98_4/U311  ( .A(\add_98_4/n244 ), .ZN(\add_98_4/n243 ) );
  NAND2_X2 \add_98_4/U310  ( .A1(\add_98_4/n203 ), .A2(\add_98_4/n202 ), .ZN(
        \add_98_4/n242 ) );
  INV_X4 \add_98_4/U309  ( .A(rnd_q[54]), .ZN(\add_98_4/n239 ) );
  INV_X4 \add_98_4/U308  ( .A(cv_q[54]), .ZN(\add_98_4/n240 ) );
  NAND2_X2 \add_98_4/U307  ( .A1(\add_98_4/n239 ), .A2(\add_98_4/n240 ), .ZN(
        \add_98_4/n199 ) );
  NAND2_X2 \add_98_4/U306  ( .A1(rnd_q[54]), .A2(cv_q[54]), .ZN(
        \add_98_4/n204 ) );
  XNOR2_X2 \add_98_4/U305  ( .A(\add_98_4/n238 ), .B(\add_98_4/n26 ), .ZN(N147) );
  NAND2_X2 \add_98_4/U304  ( .A1(\add_98_4/n203 ), .A2(\add_98_4/n202 ), .ZN(
        \add_98_4/n237 ) );
  NAND2_X2 \add_98_4/U303  ( .A1(\add_98_4/n237 ), .A2(\add_98_4/n199 ), .ZN(
        \add_98_4/n234 ) );
  NAND2_X2 \add_98_4/U302  ( .A1(\add_98_4/n236 ), .A2(\add_98_4/n199 ), .ZN(
        \add_98_4/n229 ) );
  INV_X4 \add_98_4/U301  ( .A(rnd_q[55]), .ZN(\add_98_4/n232 ) );
  INV_X4 \add_98_4/U300  ( .A(cv_q[55]), .ZN(\add_98_4/n233 ) );
  NAND2_X2 \add_98_4/U299  ( .A1(\add_98_4/n232 ), .A2(\add_98_4/n233 ), .ZN(
        \add_98_4/n200 ) );
  NAND2_X2 \add_98_4/U298  ( .A1(rnd_q[55]), .A2(cv_q[55]), .ZN(
        \add_98_4/n152 ) );
  NAND2_X2 \add_98_4/U297  ( .A1(\add_98_4/n200 ), .A2(\add_98_4/n152 ), .ZN(
        \add_98_4/n231 ) );
  XNOR2_X2 \add_98_4/U296  ( .A(\add_98_4/n230 ), .B(\add_98_4/n231 ), .ZN(
        N148) );
  INV_X4 \add_98_4/U295  ( .A(\add_98_4/n229 ), .ZN(\add_98_4/n228 ) );
  NAND2_X2 \add_98_4/U294  ( .A1(\add_98_4/n228 ), .A2(\add_98_4/n200 ), .ZN(
        \add_98_4/n147 ) );
  NAND2_X2 \add_98_4/U293  ( .A1(rnd_q[37]), .A2(cv_q[37]), .ZN(
        \add_98_4/n227 ) );
  NAND2_X2 \add_98_4/U292  ( .A1(\add_98_4/n66 ), .A2(\add_98_4/n227 ), .ZN(
        \add_98_4/n226 ) );
  NAND2_X2 \add_98_4/U291  ( .A1(\add_98_4/n225 ), .A2(\add_98_4/n226 ), .ZN(
        \add_98_4/n224 ) );
  NAND2_X2 \add_98_4/U290  ( .A1(\add_98_4/n35 ), .A2(\add_98_4/n224 ), .ZN(
        \add_98_4/n222 ) );
  INV_X4 \add_98_4/U289  ( .A(\add_98_4/n215 ), .ZN(\add_98_4/n223 ) );
  NAND4_X2 \add_98_4/U288  ( .A1(\add_98_4/n222 ), .A2(\add_98_4/n3 ), .A3(
        \add_98_4/n314 ), .A4(\add_98_4/n223 ), .ZN(\add_98_4/n207 ) );
  NAND2_X2 \add_98_4/U287  ( .A1(rnd_q[33]), .A2(cv_q[33]), .ZN(
        \add_98_4/n220 ) );
  NAND2_X2 \add_98_4/U286  ( .A1(\add_98_4/n220 ), .A2(\add_98_4/n221 ), .ZN(
        \add_98_4/n219 ) );
  NAND2_X2 \add_98_4/U285  ( .A1(\add_98_4/n1 ), .A2(\add_98_4/n219 ), .ZN(
        \add_98_4/n217 ) );
  NAND2_X2 \add_98_4/U284  ( .A1(\add_98_4/n205 ), .A2(\add_98_4/n206 ), .ZN(
        \add_98_4/n189 ) );
  INV_X4 \add_98_4/U283  ( .A(\add_98_4/n146 ), .ZN(\add_98_4/n198 ) );
  NAND2_X2 \add_98_4/U282  ( .A1(\add_98_4/n198 ), .A2(\add_98_4/n152 ), .ZN(
        \add_98_4/n191 ) );
  INV_X4 \add_98_4/U281  ( .A(\add_98_4/n197 ), .ZN(\add_98_4/n194 ) );
  INV_X4 \add_98_4/U280  ( .A(\add_98_4/n196 ), .ZN(\add_98_4/n195 ) );
  NAND2_X2 \add_98_4/U279  ( .A1(\add_98_4/n189 ), .A2(\add_98_4/n190 ), .ZN(
        \add_98_4/n163 ) );
  NAND2_X2 \add_98_4/U278  ( .A1(rnd_q[56]), .A2(cv_q[56]), .ZN(
        \add_98_4/n187 ) );
  NAND2_X2 \add_98_4/U277  ( .A1(\add_98_4/n187 ), .A2(\add_98_4/n172 ), .ZN(
        \add_98_4/n188 ) );
  XNOR2_X2 \add_98_4/U276  ( .A(\add_98_4/n163 ), .B(\add_98_4/n188 ), .ZN(
        N149) );
  INV_X4 \add_98_4/U275  ( .A(\add_98_4/n181 ), .ZN(\add_98_4/n172 ) );
  NAND2_X2 \add_98_4/U274  ( .A1(\add_98_4/n172 ), .A2(\add_98_4/n163 ), .ZN(
        \add_98_4/n186 ) );
  NAND2_X2 \add_98_4/U273  ( .A1(\add_98_4/n186 ), .A2(\add_98_4/n187 ), .ZN(
        \add_98_4/n182 ) );
  NAND2_X2 \add_98_4/U272  ( .A1(rnd_q[57]), .A2(cv_q[57]), .ZN(
        \add_98_4/n161 ) );
  INV_X4 \add_98_4/U271  ( .A(rnd_q[57]), .ZN(\add_98_4/n184 ) );
  INV_X4 \add_98_4/U270  ( .A(cv_q[57]), .ZN(\add_98_4/n185 ) );
  NAND2_X2 \add_98_4/U269  ( .A1(\add_98_4/n184 ), .A2(\add_98_4/n185 ), .ZN(
        \add_98_4/n171 ) );
  NAND2_X2 \add_98_4/U268  ( .A1(\add_98_4/n161 ), .A2(\add_98_4/n171 ), .ZN(
        \add_98_4/n183 ) );
  XNOR2_X2 \add_98_4/U267  ( .A(\add_98_4/n182 ), .B(\add_98_4/n183 ), .ZN(
        N150) );
  INV_X4 \add_98_4/U266  ( .A(\add_98_4/n163 ), .ZN(\add_98_4/n180 ) );
  INV_X4 \add_98_4/U265  ( .A(\add_98_4/n171 ), .ZN(\add_98_4/n178 ) );
  NAND2_X2 \add_98_4/U264  ( .A1(cv_q[56]), .A2(rnd_q[56]), .ZN(
        \add_98_4/n179 ) );
  NAND2_X2 \add_98_4/U263  ( .A1(\add_98_4/n9 ), .A2(\add_98_4/n161 ), .ZN(
        \add_98_4/n177 ) );
  INV_X4 \add_98_4/U262  ( .A(rnd_q[58]), .ZN(\add_98_4/n174 ) );
  INV_X4 \add_98_4/U261  ( .A(cv_q[58]), .ZN(\add_98_4/n175 ) );
  NAND2_X2 \add_98_4/U260  ( .A1(\add_98_4/n174 ), .A2(\add_98_4/n175 ), .ZN(
        \add_98_4/n159 ) );
  NAND2_X2 \add_98_4/U259  ( .A1(rnd_q[58]), .A2(cv_q[58]), .ZN(
        \add_98_4/n162 ) );
  XNOR2_X2 \add_98_4/U258  ( .A(\add_98_4/n173 ), .B(\add_98_4/n25 ), .ZN(N151) );
  NAND2_X2 \add_98_4/U257  ( .A1(\add_98_4/n31 ), .A2(\add_98_4/n163 ), .ZN(
        \add_98_4/n168 ) );
  NAND2_X2 \add_98_4/U256  ( .A1(\add_98_4/n170 ), .A2(\add_98_4/n159 ), .ZN(
        \add_98_4/n169 ) );
  NAND2_X2 \add_98_4/U255  ( .A1(\add_98_4/n168 ), .A2(\add_98_4/n169 ), .ZN(
        \add_98_4/n164 ) );
  INV_X4 \add_98_4/U254  ( .A(rnd_q[59]), .ZN(\add_98_4/n166 ) );
  INV_X4 \add_98_4/U253  ( .A(cv_q[59]), .ZN(\add_98_4/n167 ) );
  NAND2_X2 \add_98_4/U252  ( .A1(\add_98_4/n166 ), .A2(\add_98_4/n167 ), .ZN(
        \add_98_4/n150 ) );
  NAND2_X2 \add_98_4/U251  ( .A1(rnd_q[59]), .A2(cv_q[59]), .ZN(
        \add_98_4/n158 ) );
  NAND2_X2 \add_98_4/U250  ( .A1(\add_98_4/n150 ), .A2(\add_98_4/n158 ), .ZN(
        \add_98_4/n165 ) );
  XNOR2_X2 \add_98_4/U249  ( .A(\add_98_4/n164 ), .B(\add_98_4/n165 ), .ZN(
        N152) );
  NAND2_X2 \add_98_4/U248  ( .A1(\add_98_4/n157 ), .A2(\add_98_4/n158 ), .ZN(
        \add_98_4/n153 ) );
  INV_X4 \add_98_4/U247  ( .A(rnd_q[60]), .ZN(\add_98_4/n155 ) );
  INV_X4 \add_98_4/U246  ( .A(cv_q[60]), .ZN(\add_98_4/n156 ) );
  NAND2_X2 \add_98_4/U245  ( .A1(\add_98_4/n155 ), .A2(\add_98_4/n156 ), .ZN(
        \add_98_4/n151 ) );
  NAND2_X2 \add_98_4/U244  ( .A1(rnd_q[60]), .A2(cv_q[60]), .ZN(
        \add_98_4/n101 ) );
  XNOR2_X2 \add_98_4/U243  ( .A(\add_98_4/n154 ), .B(\add_98_4/n27 ), .ZN(N153) );
  INV_X4 \add_98_4/U242  ( .A(\add_98_4/n152 ), .ZN(\add_98_4/n149 ) );
  INV_X4 \add_98_4/U241  ( .A(\add_98_4/n122 ), .ZN(\add_98_4/n104 ) );
  INV_X4 \add_98_4/U240  ( .A(\add_98_4/n101 ), .ZN(\add_98_4/n148 ) );
  INV_X4 \add_98_4/U239  ( .A(\add_98_4/n147 ), .ZN(\add_98_4/n103 ) );
  INV_X4 \add_98_4/U238  ( .A(\add_98_4/n129 ), .ZN(\add_98_4/n87 ) );
  NAND2_X2 \add_98_4/U237  ( .A1(\add_98_4/n126 ), .A2(\add_98_4/n127 ), .ZN(
        \add_98_4/n102 ) );
  NAND2_X2 \add_98_4/U236  ( .A1(\add_98_4/n102 ), .A2(\add_98_4/n13 ), .ZN(
        \add_98_4/n145 ) );
  NAND2_X2 \add_98_4/U235  ( .A1(\add_98_4/n146 ), .A2(\add_98_4/n104 ), .ZN(
        \add_98_4/n93 ) );
  NAND4_X2 \add_98_4/U234  ( .A1(\add_98_4/n143 ), .A2(\add_98_4/n144 ), .A3(
        \add_98_4/n145 ), .A4(\add_98_4/n93 ), .ZN(\add_98_4/n139 ) );
  NAND2_X2 \add_98_4/U233  ( .A1(rnd_q[61]), .A2(cv_q[61]), .ZN(\add_98_4/n91 ) );
  INV_X4 \add_98_4/U232  ( .A(rnd_q[61]), .ZN(\add_98_4/n141 ) );
  INV_X4 \add_98_4/U231  ( .A(cv_q[61]), .ZN(\add_98_4/n142 ) );
  NAND2_X2 \add_98_4/U230  ( .A1(\add_98_4/n141 ), .A2(\add_98_4/n142 ), .ZN(
        \add_98_4/n117 ) );
  NAND2_X2 \add_98_4/U229  ( .A1(\add_98_4/n91 ), .A2(\add_98_4/n117 ), .ZN(
        \add_98_4/n140 ) );
  XNOR2_X2 \add_98_4/U228  ( .A(\add_98_4/n139 ), .B(\add_98_4/n140 ), .ZN(
        N154) );
  XNOR2_X2 \add_98_4/U227  ( .A(\add_98_4/n80 ), .B(\add_98_4/n136 ), .ZN(N127) );
  INV_X4 \add_98_4/U226  ( .A(\add_98_4/n134 ), .ZN(\add_98_4/n130 ) );
  NAND2_X2 \add_98_4/U225  ( .A1(\add_98_4/n132 ), .A2(\add_98_4/n133 ), .ZN(
        \add_98_4/n131 ) );
  NAND2_X2 \add_98_4/U224  ( .A1(\add_98_4/n126 ), .A2(\add_98_4/n127 ), .ZN(
        \add_98_4/n125 ) );
  NAND2_X2 \add_98_4/U223  ( .A1(\add_98_4/n103 ), .A2(\add_98_4/n117 ), .ZN(
        \add_98_4/n123 ) );
  NAND2_X2 \add_98_4/U222  ( .A1(\add_98_4/n21 ), .A2(\add_98_4/n117 ), .ZN(
        \add_98_4/n113 ) );
  INV_X4 \add_98_4/U221  ( .A(\add_98_4/n93 ), .ZN(\add_98_4/n120 ) );
  NAND2_X2 \add_98_4/U220  ( .A1(\add_98_4/n120 ), .A2(\add_98_4/n117 ), .ZN(
        \add_98_4/n114 ) );
  INV_X4 \add_98_4/U219  ( .A(\add_98_4/n91 ), .ZN(\add_98_4/n118 ) );
  INV_X4 \add_98_4/U218  ( .A(\add_98_4/n117 ), .ZN(\add_98_4/n105 ) );
  NAND2_X2 \add_98_4/U217  ( .A1(\add_98_4/n11 ), .A2(\add_98_4/n117 ), .ZN(
        \add_98_4/n116 ) );
  NAND4_X2 \add_98_4/U216  ( .A1(\add_98_4/n113 ), .A2(\add_98_4/n114 ), .A3(
        \add_98_4/n115 ), .A4(\add_98_4/n116 ), .ZN(\add_98_4/n112 ) );
  INV_X4 \add_98_4/U215  ( .A(rnd_q[62]), .ZN(\add_98_4/n109 ) );
  INV_X4 \add_98_4/U214  ( .A(cv_q[62]), .ZN(\add_98_4/n110 ) );
  NAND2_X2 \add_98_4/U213  ( .A1(rnd_q[62]), .A2(cv_q[62]), .ZN(
        \add_98_4/n100 ) );
  INV_X4 \add_98_4/U212  ( .A(\add_98_4/n100 ), .ZN(\add_98_4/n108 ) );
  XNOR2_X2 \add_98_4/U211  ( .A(\add_98_4/n106 ), .B(\add_98_4/n107 ), .ZN(
        N155) );
  NAND2_X2 \add_98_4/U210  ( .A1(\add_98_4/n12 ), .A2(\add_98_4/n102 ), .ZN(
        \add_98_4/n83 ) );
  NAND2_X2 \add_98_4/U209  ( .A1(\add_98_4/n94 ), .A2(\add_98_4/n148 ), .ZN(
        \add_98_4/n99 ) );
  NAND2_X2 \add_98_4/U208  ( .A1(\add_98_4/n99 ), .A2(\add_98_4/n100 ), .ZN(
        \add_98_4/n95 ) );
  NAND2_X2 \add_98_4/U207  ( .A1(\add_98_4/n21 ), .A2(\add_98_4/n94 ), .ZN(
        \add_98_4/n97 ) );
  NAND2_X2 \add_98_4/U206  ( .A1(\add_98_4/n11 ), .A2(\add_98_4/n94 ), .ZN(
        \add_98_4/n98 ) );
  NAND2_X2 \add_98_4/U205  ( .A1(\add_98_4/n97 ), .A2(\add_98_4/n98 ), .ZN(
        \add_98_4/n96 ) );
  INV_X4 \add_98_4/U204  ( .A(\add_98_4/n94 ), .ZN(\add_98_4/n92 ) );
  NAND4_X2 \add_98_4/U203  ( .A1(\add_98_4/n83 ), .A2(\add_98_4/n84 ), .A3(
        \add_98_4/n85 ), .A4(\add_98_4/n86 ), .ZN(\add_98_4/n81 ) );
  XNOR2_X2 \add_98_4/U202  ( .A(rnd_q[63]), .B(cv_q[63]), .ZN(\add_98_4/n82 )
         );
  XNOR2_X2 \add_98_4/U201  ( .A(\add_98_4/n81 ), .B(\add_98_4/n82 ), .ZN(N156)
         );
  XNOR2_X2 \add_98_4/U200  ( .A(\add_98_4/n74 ), .B(\add_98_4/n75 ), .ZN(N128)
         );
  INV_X4 \add_98_4/U199  ( .A(\add_98_4/n66 ), .ZN(\add_98_4/n72 ) );
  XNOR2_X2 \add_98_4/U198  ( .A(\add_98_4/n30 ), .B(\add_98_4/n73 ), .ZN(N129)
         );
  INV_X4 \add_98_4/U197  ( .A(\add_98_4/n63 ), .ZN(\add_98_4/n70 ) );
  XNOR2_X2 \add_98_4/U196  ( .A(\add_98_4/n68 ), .B(\add_98_4/n69 ), .ZN(N130)
         );
  NAND2_X2 \add_98_4/U195  ( .A1(rnd_q[38]), .A2(cv_q[38]), .ZN(\add_98_4/n58 ) );
  NAND2_X2 \add_98_4/U194  ( .A1(\add_98_4/n58 ), .A2(\add_98_4/n6 ), .ZN(
        \add_98_4/n61 ) );
  NAND2_X2 \add_98_4/U193  ( .A1(\add_98_4/n30 ), .A2(\add_98_4/n66 ), .ZN(
        \add_98_4/n65 ) );
  NAND2_X2 \add_98_4/U192  ( .A1(\add_98_4/n64 ), .A2(\add_98_4/n65 ), .ZN(
        \add_98_4/n62 ) );
  NAND2_X2 \add_98_4/U191  ( .A1(\add_98_4/n62 ), .A2(\add_98_4/n63 ), .ZN(
        \add_98_4/n59 ) );
  XNOR2_X2 \add_98_4/U190  ( .A(\add_98_4/n61 ), .B(\add_98_4/n59 ), .ZN(N131)
         );
  NAND2_X2 \add_98_4/U189  ( .A1(\add_98_4/n59 ), .A2(\add_98_4/n6 ), .ZN(
        \add_98_4/n57 ) );
  NAND2_X2 \add_98_4/U188  ( .A1(\add_98_4/n57 ), .A2(\add_98_4/n58 ), .ZN(
        \add_98_4/n54 ) );
  NAND2_X2 \add_98_4/U187  ( .A1(\add_98_4/n56 ), .A2(\add_98_4/n3 ), .ZN(
        \add_98_4/n55 ) );
  XNOR2_X2 \add_98_4/U186  ( .A(\add_98_4/n54 ), .B(\add_98_4/n55 ), .ZN(N132)
         );
  INV_X4 \add_98_4/U185  ( .A(\add_98_4/n52 ), .ZN(\add_98_4/n45 ) );
  XNOR2_X2 \add_98_4/U184  ( .A(\add_98_4/n50 ), .B(\add_98_4/n51 ), .ZN(N133)
         );
  XNOR2_X2 \add_98_4/U183  ( .A(\add_98_4/n41 ), .B(\add_98_4/n42 ), .ZN(N134)
         );
  NAND2_X2 \add_98_4/U182  ( .A1(\add_98_4/n260 ), .A2(\add_98_4/n134 ), .ZN(
        \add_98_4/n259 ) );
  NOR2_X2 \add_98_4/U181  ( .A1(\add_98_4/n20 ), .A2(\add_98_4/n108 ), .ZN(
        \add_98_4/n107 ) );
  NOR2_X2 \add_98_4/U180  ( .A1(\add_98_4/n244 ), .A2(\add_98_4/n250 ), .ZN(
        \add_98_4/n249 ) );
  AND2_X2 \add_98_4/U179  ( .A1(cv_q[40]), .A2(rnd_q[40]), .ZN(\add_98_4/n354 ) );
  NOR2_X2 \add_98_4/U178  ( .A1(\add_98_4/n39 ), .A2(\add_98_4/n252 ), .ZN(
        \add_98_4/n253 ) );
  NOR2_X2 \add_98_4/U177  ( .A1(\add_98_4/n40 ), .A2(\add_98_4/n43 ), .ZN(
        \add_98_4/n42 ) );
  NOR2_X2 \add_98_4/U176  ( .A1(\add_98_4/n76 ), .A2(\add_98_4/n77 ), .ZN(
        \add_98_4/n75 ) );
  NOR2_X2 \add_98_4/U175  ( .A1(\add_98_4/n262 ), .A2(\add_98_4/n137 ), .ZN(
        \add_98_4/n261 ) );
  AND2_X2 \add_98_4/U174  ( .A1(rnd_q[41]), .A2(cv_q[41]), .ZN(\add_98_4/n40 )
         );
  AND2_X2 \add_98_4/U173  ( .A1(rnd_q[52]), .A2(cv_q[52]), .ZN(\add_98_4/n39 )
         );
  AND2_X2 \add_98_4/U172  ( .A1(rnd_q[34]), .A2(cv_q[34]), .ZN(\add_98_4/n38 )
         );
  OR2_X2 \add_98_4/U171  ( .A1(cv_q[49]), .A2(rnd_q[49]), .ZN(\add_98_4/n37 )
         );
  NOR2_X2 \add_98_4/U170  ( .A1(cv_q[49]), .A2(rnd_q[49]), .ZN(\add_98_4/n280 ) );
  NOR2_X2 \add_98_4/U169  ( .A1(\add_98_4/n280 ), .A2(\add_98_4/n281 ), .ZN(
        \add_98_4/n273 ) );
  NOR2_X2 \add_98_4/U168  ( .A1(cv_q[37]), .A2(rnd_q[37]), .ZN(\add_98_4/n297 ) );
  NOR2_X2 \add_98_4/U167  ( .A1(cv_q[38]), .A2(rnd_q[38]), .ZN(\add_98_4/n298 ) );
  NOR2_X2 \add_98_4/U166  ( .A1(\add_98_4/n297 ), .A2(\add_98_4/n298 ), .ZN(
        \add_98_4/n225 ) );
  NOR2_X2 \add_98_4/U165  ( .A1(rnd_q[36]), .A2(cv_q[36]), .ZN(\add_98_4/n36 )
         );
  NOR2_X2 \add_98_4/U164  ( .A1(cv_q[41]), .A2(rnd_q[41]), .ZN(\add_98_4/n356 ) );
  NOR2_X2 \add_98_4/U163  ( .A1(\add_98_4/n356 ), .A2(\add_98_4/n357 ), .ZN(
        \add_98_4/n355 ) );
  AND2_X2 \add_98_4/U162  ( .A1(\add_98_4/n56 ), .A2(\add_98_4/n377 ), .ZN(
        \add_98_4/n35 ) );
  NOR2_X2 \add_98_4/U161  ( .A1(cv_q[49]), .A2(rnd_q[49]), .ZN(\add_98_4/n283 ) );
  NOR2_X2 \add_98_4/U160  ( .A1(\add_98_4/n309 ), .A2(\add_98_4/n313 ), .ZN(
        \add_98_4/n311 ) );
  NOR2_X2 \add_98_4/U159  ( .A1(cv_q[52]), .A2(rnd_q[52]), .ZN(\add_98_4/n247 ) );
  NOR2_X2 \add_98_4/U158  ( .A1(cv_q[53]), .A2(rnd_q[53]), .ZN(\add_98_4/n246 ) );
  NOR2_X2 \add_98_4/U157  ( .A1(\add_98_4/n246 ), .A2(\add_98_4/n247 ), .ZN(
        \add_98_4/n236 ) );
  NOR2_X2 \add_98_4/U156  ( .A1(cv_q[37]), .A2(rnd_q[37]), .ZN(\add_98_4/n387 ) );
  NOR2_X2 \add_98_4/U155  ( .A1(\add_98_4/n46 ), .A2(\add_98_4/n45 ), .ZN(
        \add_98_4/n51 ) );
  NOR2_X2 \add_98_4/U154  ( .A1(\add_98_4/n38 ), .A2(\add_98_4/n79 ), .ZN(
        \add_98_4/n136 ) );
  NOR2_X2 \add_98_4/U153  ( .A1(\add_98_4/n344 ), .A2(\add_98_4/n319 ), .ZN(
        \add_98_4/n343 ) );
  NOR2_X2 \add_98_4/U152  ( .A1(\add_98_4/n70 ), .A2(\add_98_4/n67 ), .ZN(
        \add_98_4/n69 ) );
  NOR2_X2 \add_98_4/U151  ( .A1(\add_98_4/n318 ), .A2(\add_98_4/n16 ), .ZN(
        \add_98_4/n320 ) );
  NOR2_X2 \add_98_4/U150  ( .A1(\add_98_4/n36 ), .A2(\add_98_4/n72 ), .ZN(
        \add_98_4/n73 ) );
  NOR2_X2 \add_98_4/U149  ( .A1(cv_q[53]), .A2(rnd_q[53]), .ZN(\add_98_4/n244 ) );
  OR2_X2 \add_98_4/U148  ( .A1(\add_98_4/n283 ), .A2(\add_98_4/n284 ), .ZN(
        \add_98_4/n34 ) );
  NAND3_X2 \add_98_4/U147  ( .A1(cv_q[52]), .A2(rnd_q[52]), .A3(
        \add_98_4/n243 ), .ZN(\add_98_4/n203 ) );
  NOR2_X2 \add_98_4/U146  ( .A1(cv_q[52]), .A2(rnd_q[52]), .ZN(\add_98_4/n252 ) );
  NOR2_X2 \add_98_4/U145  ( .A1(cv_q[33]), .A2(rnd_q[33]), .ZN(\add_98_4/n137 ) );
  NOR2_X2 \add_98_4/U144  ( .A1(cv_q[48]), .A2(rnd_q[48]), .ZN(\add_98_4/n281 ) );
  NOR2_X2 \add_98_4/U143  ( .A1(cv_q[38]), .A2(rnd_q[38]), .ZN(\add_98_4/n60 )
         );
  NOR2_X2 \add_98_4/U142  ( .A1(cv_q[56]), .A2(rnd_q[56]), .ZN(\add_98_4/n181 ) );
  NOR2_X2 \add_98_4/U141  ( .A1(cv_q[37]), .A2(rnd_q[37]), .ZN(\add_98_4/n67 )
         );
  NOR2_X2 \add_98_4/U140  ( .A1(\add_98_4/n76 ), .A2(\add_98_4/n383 ), .ZN(
        \add_98_4/n218 ) );
  NOR2_X2 \add_98_4/U139  ( .A1(cv_q[40]), .A2(rnd_q[40]), .ZN(\add_98_4/n46 )
         );
  NOR2_X2 \add_98_4/U138  ( .A1(cv_q[41]), .A2(rnd_q[41]), .ZN(\add_98_4/n43 )
         );
  NOR2_X2 \add_98_4/U137  ( .A1(cv_q[46]), .A2(rnd_q[46]), .ZN(\add_98_4/n309 ) );
  NOR2_X2 \add_98_4/U136  ( .A1(cv_q[44]), .A2(rnd_q[44]), .ZN(\add_98_4/n319 ) );
  NOR3_X2 \add_98_4/U135  ( .A1(\add_98_4/n308 ), .A2(\add_98_4/n309 ), .A3(
        \add_98_4/n310 ), .ZN(\add_98_4/n307 ) );
  NOR2_X2 \add_98_4/U134  ( .A1(cv_q[45]), .A2(rnd_q[45]), .ZN(\add_98_4/n310 ) );
  NAND3_X2 \add_98_4/U133  ( .A1(\add_98_4/n202 ), .A2(\add_98_4/n203 ), .A3(
        \add_98_4/n204 ), .ZN(\add_98_4/n201 ) );
  AND2_X4 \add_98_4/U132  ( .A1(\add_98_4/n199 ), .A2(\add_98_4/n200 ), .ZN(
        \add_98_4/n33 ) );
  AND2_X2 \add_98_4/U131  ( .A1(\add_98_4/n201 ), .A2(\add_98_4/n33 ), .ZN(
        \add_98_4/n146 ) );
  NOR2_X2 \add_98_4/U130  ( .A1(\add_98_4/n348 ), .A2(\add_98_4/n349 ), .ZN(
        \add_98_4/n347 ) );
  NAND3_X2 \add_98_4/U129  ( .A1(\add_98_4/n346 ), .A2(\add_98_4/n15 ), .A3(
        \add_98_4/n347 ), .ZN(\add_98_4/n316 ) );
  NOR2_X2 \add_98_4/U128  ( .A1(\add_98_4/n263 ), .A2(\add_98_4/n218 ), .ZN(
        \add_98_4/n303 ) );
  NAND3_X2 \add_98_4/U127  ( .A1(\add_98_4/n378 ), .A2(\add_98_4/n372 ), .A3(
        \add_98_4/n379 ), .ZN(\add_98_4/n370 ) );
  NOR2_X2 \add_98_4/U126  ( .A1(\add_98_4/n40 ), .A2(\add_98_4/n388 ), .ZN(
        \add_98_4/n369 ) );
  NAND3_X2 \add_98_4/U125  ( .A1(\add_98_4/n369 ), .A2(\add_98_4/n370 ), .A3(
        \add_98_4/n371 ), .ZN(\add_98_4/n367 ) );
  NAND3_X2 \add_98_4/U124  ( .A1(\add_98_4/n337 ), .A2(\add_98_4/n4 ), .A3(
        \add_98_4/n7 ), .ZN(\add_98_4/n336 ) );
  NAND3_X2 \add_98_4/U123  ( .A1(\add_98_4/n24 ), .A2(\add_98_4/n330 ), .A3(
        \add_98_4/n336 ), .ZN(\add_98_4/n334 ) );
  NOR2_X2 \add_98_4/U122  ( .A1(\add_98_4/n79 ), .A2(\add_98_4/n80 ), .ZN(
        \add_98_4/n78 ) );
  NOR2_X2 \add_98_4/U121  ( .A1(\add_98_4/n78 ), .A2(\add_98_4/n38 ), .ZN(
        \add_98_4/n74 ) );
  NOR2_X2 \add_98_4/U120  ( .A1(\add_98_4/n18 ), .A2(\add_98_4/n153 ), .ZN(
        \add_98_4/n154 ) );
  NOR2_X2 \add_98_4/U119  ( .A1(\add_98_4/n60 ), .A2(\add_98_4/n67 ), .ZN(
        \add_98_4/n375 ) );
  NOR2_X2 \add_98_4/U118  ( .A1(\add_98_4/n235 ), .A2(\add_98_4/n245 ), .ZN(
        \add_98_4/n241 ) );
  NOR2_X2 \add_98_4/U117  ( .A1(\add_98_4/n241 ), .A2(\add_98_4/n242 ), .ZN(
        \add_98_4/n238 ) );
  NOR2_X2 \add_98_4/U116  ( .A1(\add_98_4/n30 ), .A2(\add_98_4/n49 ), .ZN(
        \add_98_4/n48 ) );
  NOR2_X2 \add_98_4/U115  ( .A1(\add_98_4/n48 ), .A2(\add_98_4/n19 ), .ZN(
        \add_98_4/n47 ) );
  NOR2_X2 \add_98_4/U114  ( .A1(\add_98_4/n46 ), .A2(\add_98_4/n47 ), .ZN(
        \add_98_4/n44 ) );
  NOR2_X2 \add_98_4/U113  ( .A1(\add_98_4/n44 ), .A2(\add_98_4/n45 ), .ZN(
        \add_98_4/n41 ) );
  NOR2_X2 \add_98_4/U112  ( .A1(\add_98_4/n252 ), .A2(\add_98_4/n235 ), .ZN(
        \add_98_4/n251 ) );
  NOR2_X2 \add_98_4/U111  ( .A1(\add_98_4/n251 ), .A2(\add_98_4/n39 ), .ZN(
        \add_98_4/n248 ) );
  NOR2_X2 \add_98_4/U110  ( .A1(\add_98_4/n30 ), .A2(\add_98_4/n36 ), .ZN(
        \add_98_4/n71 ) );
  NOR2_X2 \add_98_4/U109  ( .A1(\add_98_4/n71 ), .A2(\add_98_4/n72 ), .ZN(
        \add_98_4/n68 ) );
  NOR3_X2 \add_98_4/U108  ( .A1(\add_98_4/n180 ), .A2(\add_98_4/n178 ), .A3(
        \add_98_4/n181 ), .ZN(\add_98_4/n176 ) );
  NOR2_X2 \add_98_4/U107  ( .A1(\add_98_4/n176 ), .A2(\add_98_4/n177 ), .ZN(
        \add_98_4/n173 ) );
  NOR2_X2 \add_98_4/U106  ( .A1(\add_98_4/n36 ), .A2(\add_98_4/n67 ), .ZN(
        \add_98_4/n64 ) );
  NAND3_X2 \add_98_4/U105  ( .A1(\add_98_4/n314 ), .A2(\add_98_4/n315 ), .A3(
        \add_98_4/n316 ), .ZN(\add_98_4/n133 ) );
  NOR2_X2 \add_98_4/U104  ( .A1(\add_98_4/n20 ), .A2(\add_98_4/n91 ), .ZN(
        \add_98_4/n90 ) );
  NOR2_X2 \add_98_4/U103  ( .A1(\add_98_4/n105 ), .A2(\add_98_4/n101 ), .ZN(
        \add_98_4/n119 ) );
  NOR2_X2 \add_98_4/U102  ( .A1(\add_98_4/n319 ), .A2(\add_98_4/n14 ), .ZN(
        \add_98_4/n325 ) );
  OR2_X4 \add_98_4/U101  ( .A1(\add_98_4/n137 ), .A2(\add_98_4/n221 ), .ZN(
        \add_98_4/n32 ) );
  AND2_X2 \add_98_4/U100  ( .A1(\add_98_4/n138 ), .A2(\add_98_4/n32 ), .ZN(
        \add_98_4/n80 ) );
  NOR2_X2 \add_98_4/U99  ( .A1(\add_98_4/n43 ), .A2(\add_98_4/n52 ), .ZN(
        \add_98_4/n388 ) );
  NAND3_X2 \add_98_4/U98  ( .A1(\add_98_4/n161 ), .A2(\add_98_4/n9 ), .A3(
        \add_98_4/n162 ), .ZN(\add_98_4/n160 ) );
  NAND3_X2 \add_98_4/U97  ( .A1(\add_98_4/n159 ), .A2(\add_98_4/n150 ), .A3(
        \add_98_4/n160 ), .ZN(\add_98_4/n157 ) );
  NOR2_X2 \add_98_4/U96  ( .A1(\add_98_4/n147 ), .A2(\add_98_4/n127 ), .ZN(
        \add_98_4/n193 ) );
  NOR3_X2 \add_98_4/U95  ( .A1(\add_98_4/n135 ), .A2(\add_98_4/n130 ), .A3(
        \add_98_4/n131 ), .ZN(\add_98_4/n128 ) );
  NOR2_X2 \add_98_4/U94  ( .A1(\add_98_4/n128 ), .A2(\add_98_4/n129 ), .ZN(
        \add_98_4/n124 ) );
  NOR2_X2 \add_98_4/U93  ( .A1(\add_98_4/n124 ), .A2(\add_98_4/n125 ), .ZN(
        \add_98_4/n121 ) );
  NOR2_X2 \add_98_4/U92  ( .A1(\add_98_4/n318 ), .A2(\add_98_4/n319 ), .ZN(
        \add_98_4/n317 ) );
  NAND3_X2 \add_98_4/U91  ( .A1(\add_98_4/n4 ), .A2(\add_98_4/n10 ), .A3(
        \add_98_4/n317 ), .ZN(\add_98_4/n214 ) );
  AND3_X2 \add_98_4/U90  ( .A1(\add_98_4/n171 ), .A2(\add_98_4/n159 ), .A3(
        \add_98_4/n172 ), .ZN(\add_98_4/n31 ) );
  NAND3_X2 \add_98_4/U89  ( .A1(\add_98_4/n150 ), .A2(\add_98_4/n151 ), .A3(
        \add_98_4/n31 ), .ZN(\add_98_4/n122 ) );
  NOR3_X2 \add_98_4/U88  ( .A1(\add_98_4/n194 ), .A2(\add_98_4/n147 ), .A3(
        \add_98_4/n195 ), .ZN(\add_98_4/n192 ) );
  NOR2_X2 \add_98_4/U87  ( .A1(\add_98_4/n319 ), .A2(\add_98_4/n14 ), .ZN(
        \add_98_4/n337 ) );
  NOR2_X2 \add_98_4/U86  ( .A1(\add_98_4/n46 ), .A2(\add_98_4/n43 ), .ZN(
        \add_98_4/n372 ) );
  NAND3_X2 \add_98_4/U85  ( .A1(\add_98_4/n216 ), .A2(\add_98_4/n217 ), .A3(
        \add_98_4/n381 ), .ZN(\add_98_4/n212 ) );
  NOR2_X2 \add_98_4/U84  ( .A1(\add_98_4/n36 ), .A2(\add_98_4/n387 ), .ZN(
        \add_98_4/n386 ) );
  NAND3_X2 \add_98_4/U83  ( .A1(\add_98_4/n3 ), .A2(\add_98_4/n6 ), .A3(
        \add_98_4/n386 ), .ZN(\add_98_4/n49 ) );
  NOR2_X2 \add_98_4/U82  ( .A1(\add_98_4/n20 ), .A2(\add_98_4/n105 ), .ZN(
        \add_98_4/n94 ) );
  AND3_X2 \add_98_4/U81  ( .A1(\add_98_4/n381 ), .A2(\add_98_4/n216 ), .A3(
        \add_98_4/n380 ), .ZN(\add_98_4/n30 ) );
  OR3_X4 \add_98_4/U80  ( .A1(\add_98_4/n311 ), .A2(\add_98_4/n312 ), .A3(
        \add_98_4/n16 ), .ZN(\add_98_4/n29 ) );
  OR2_X2 \add_98_4/U79  ( .A1(\add_98_4/n29 ), .A2(\add_98_4/n307 ), .ZN(
        \add_98_4/n305 ) );
  NOR2_X2 \add_98_4/U78  ( .A1(\add_98_4/n210 ), .A2(\add_98_4/n211 ), .ZN(
        \add_98_4/n209 ) );
  NAND3_X2 \add_98_4/U77  ( .A1(\add_98_4/n212 ), .A2(\add_98_4/n213 ), .A3(
        \add_98_4/n378 ), .ZN(\add_98_4/n208 ) );
  NAND3_X2 \add_98_4/U76  ( .A1(\add_98_4/n208 ), .A2(\add_98_4/n209 ), .A3(
        \add_98_4/n207 ), .ZN(\add_98_4/n206 ) );
  NAND3_X2 \add_98_4/U75  ( .A1(\add_98_4/n234 ), .A2(\add_98_4/n204 ), .A3(
        \add_98_4/n17 ), .ZN(\add_98_4/n230 ) );
  NAND3_X2 \add_98_4/U74  ( .A1(\add_98_4/n162 ), .A2(\add_98_4/n9 ), .A3(
        \add_98_4/n161 ), .ZN(\add_98_4/n170 ) );
  NOR3_X2 \add_98_4/U73  ( .A1(\add_98_4/n259 ), .A2(\add_98_4/n211 ), .A3(
        \add_98_4/n210 ), .ZN(\add_98_4/n256 ) );
  NOR2_X2 \add_98_4/U72  ( .A1(\add_98_4/n256 ), .A2(\add_98_4/n129 ), .ZN(
        \add_98_4/n254 ) );
  NOR2_X2 \add_98_4/U71  ( .A1(\add_98_4/n254 ), .A2(\add_98_4/n255 ), .ZN(
        \add_98_4/n235 ) );
  NOR3_X2 \add_98_4/U70  ( .A1(\add_98_4/n218 ), .A2(\add_98_4/n77 ), .A3(
        \add_98_4/n1 ), .ZN(\add_98_4/n302 ) );
  NOR2_X2 \add_98_4/U69  ( .A1(\add_98_4/n352 ), .A2(\add_98_4/n362 ), .ZN(
        \add_98_4/n361 ) );
  NAND3_X2 \add_98_4/U68  ( .A1(\add_98_4/n359 ), .A2(\add_98_4/n360 ), .A3(
        \add_98_4/n361 ), .ZN(\add_98_4/n215 ) );
  NOR2_X2 \add_98_4/U67  ( .A1(\add_98_4/n214 ), .A2(\add_98_4/n215 ), .ZN(
        \add_98_4/n293 ) );
  NOR3_X2 \add_98_4/U66  ( .A1(\add_98_4/n191 ), .A2(\add_98_4/n192 ), .A3(
        \add_98_4/n193 ), .ZN(\add_98_4/n190 ) );
  NOR2_X2 \add_98_4/U65  ( .A1(\add_98_4/n30 ), .A2(\add_98_4/n49 ), .ZN(
        \add_98_4/n363 ) );
  NOR2_X2 \add_98_4/U64  ( .A1(\add_98_4/n363 ), .A2(\add_98_4/n19 ), .ZN(
        \add_98_4/n358 ) );
  NOR2_X2 \add_98_4/U63  ( .A1(\add_98_4/n358 ), .A2(\add_98_4/n215 ), .ZN(
        \add_98_4/n345 ) );
  NOR2_X2 \add_98_4/U62  ( .A1(\add_98_4/n345 ), .A2(\add_98_4/n328 ), .ZN(
        \add_98_4/n342 ) );
  NOR2_X2 \add_98_4/U61  ( .A1(\add_98_4/n118 ), .A2(\add_98_4/n119 ), .ZN(
        \add_98_4/n115 ) );
  NOR3_X2 \add_98_4/U60  ( .A1(\add_98_4/n121 ), .A2(\add_98_4/n122 ), .A3(
        \add_98_4/n123 ), .ZN(\add_98_4/n111 ) );
  NOR2_X2 \add_98_4/U59  ( .A1(\add_98_4/n111 ), .A2(\add_98_4/n112 ), .ZN(
        \add_98_4/n106 ) );
  NOR2_X2 \add_98_4/U58  ( .A1(\add_98_4/n30 ), .A2(\add_98_4/n49 ), .ZN(
        \add_98_4/n53 ) );
  NOR2_X2 \add_98_4/U57  ( .A1(\add_98_4/n53 ), .A2(\add_98_4/n19 ), .ZN(
        \add_98_4/n50 ) );
  NOR2_X2 \add_98_4/U56  ( .A1(\add_98_4/n272 ), .A2(\add_98_4/n258 ), .ZN(
        \add_98_4/n267 ) );
  NOR2_X2 \add_98_4/U55  ( .A1(\add_98_4/n267 ), .A2(\add_98_4/n197 ), .ZN(
        \add_98_4/n264 ) );
  NOR2_X2 \add_98_4/U54  ( .A1(\add_98_4/n129 ), .A2(\add_98_4/n147 ), .ZN(
        \add_98_4/n205 ) );
  NOR2_X2 \add_98_4/U53  ( .A1(\add_98_4/n92 ), .A2(\add_98_4/n93 ), .ZN(
        \add_98_4/n89 ) );
  NOR2_X2 \add_98_4/U52  ( .A1(\add_98_4/n214 ), .A2(\add_98_4/n215 ), .ZN(
        \add_98_4/n213 ) );
  NOR2_X2 \add_98_4/U51  ( .A1(\add_98_4/n325 ), .A2(\add_98_4/n326 ), .ZN(
        \add_98_4/n324 ) );
  NOR3_X2 \add_98_4/U50  ( .A1(\add_98_4/n323 ), .A2(\add_98_4/n324 ), .A3(
        \add_98_4/n22 ), .ZN(\add_98_4/n322 ) );
  NOR2_X2 \add_98_4/U49  ( .A1(\add_98_4/n312 ), .A2(\add_98_4/n322 ), .ZN(
        \add_98_4/n321 ) );
  NOR2_X2 \add_98_4/U48  ( .A1(\add_98_4/n30 ), .A2(\add_98_4/n49 ), .ZN(
        \add_98_4/n327 ) );
  NAND3_X2 \add_98_4/U47  ( .A1(\add_98_4/n88 ), .A2(\add_98_4/n13 ), .A3(
        \add_98_4/n87 ), .ZN(\add_98_4/n144 ) );
  NOR3_X2 \add_98_4/U46  ( .A1(\add_98_4/n11 ), .A2(\add_98_4/n21 ), .A3(
        \add_98_4/n148 ), .ZN(\add_98_4/n143 ) );
  NOR2_X2 \add_98_4/U45  ( .A1(\add_98_4/n95 ), .A2(\add_98_4/n96 ), .ZN(
        \add_98_4/n84 ) );
  NOR2_X2 \add_98_4/U44  ( .A1(\add_98_4/n89 ), .A2(\add_98_4/n90 ), .ZN(
        \add_98_4/n85 ) );
  NOR4_X2 \add_98_4/U43  ( .A1(\add_98_4/n327 ), .A2(\add_98_4/n328 ), .A3(
        \add_98_4/n19 ), .A4(\add_98_4/n326 ), .ZN(\add_98_4/n323 ) );
  NOR2_X2 \add_98_4/U42  ( .A1(\add_98_4/n262 ), .A2(\add_98_4/n77 ), .ZN(
        \add_98_4/n304 ) );
  NOR2_X2 \add_98_4/U41  ( .A1(\add_98_4/n49 ), .A2(\add_98_4/n302 ), .ZN(
        \add_98_4/n301 ) );
  NOR2_X2 \add_98_4/U40  ( .A1(\add_98_4/n214 ), .A2(\add_98_4/n215 ), .ZN(
        \add_98_4/n299 ) );
  NAND3_X2 \add_98_4/U39  ( .A1(\add_98_4/n299 ), .A2(\add_98_4/n300 ), .A3(
        \add_98_4/n301 ), .ZN(\add_98_4/n134 ) );
  NAND3_X2 \add_98_4/U38  ( .A1(\add_98_4/n87 ), .A2(\add_98_4/n88 ), .A3(
        \add_98_4/n12 ), .ZN(\add_98_4/n86 ) );
  NOR2_X2 \add_98_4/U37  ( .A1(\add_98_4/n211 ), .A2(\add_98_4/n210 ), .ZN(
        \add_98_4/n291 ) );
  NAND3_X2 \add_98_4/U36  ( .A1(\add_98_4/n291 ), .A2(\add_98_4/n134 ), .A3(
        \add_98_4/n260 ), .ZN(\add_98_4/n88 ) );
  OR2_X4 \add_98_4/U35  ( .A1(rnd_q[32]), .A2(cv_q[32]), .ZN(\add_98_4/n382 )
         );
  NOR2_X1 \add_98_4/U34  ( .A1(cv_q[42]), .A2(rnd_q[42]), .ZN(\add_98_4/n357 )
         );
  NOR2_X1 \add_98_4/U33  ( .A1(cv_q[34]), .A2(rnd_q[34]), .ZN(\add_98_4/n79 )
         );
  NOR2_X1 \add_98_4/U32  ( .A1(cv_q[35]), .A2(rnd_q[35]), .ZN(\add_98_4/n76 )
         );
  OR2_X4 \add_98_4/U31  ( .A1(rnd_q[43]), .A2(cv_q[43]), .ZN(\add_98_4/n315 )
         );
  NOR2_X1 \add_98_4/U30  ( .A1(cv_q[42]), .A2(rnd_q[42]), .ZN(\add_98_4/n352 )
         );
  AND2_X4 \add_98_4/U29  ( .A1(\add_98_4/n382 ), .A2(\add_98_4/n221 ), .ZN(
        N125) );
  AND2_X4 \add_98_4/U28  ( .A1(\add_98_4/n151 ), .A2(\add_98_4/n101 ), .ZN(
        \add_98_4/n27 ) );
  AND2_X4 \add_98_4/U27  ( .A1(\add_98_4/n199 ), .A2(\add_98_4/n204 ), .ZN(
        \add_98_4/n26 ) );
  AND2_X4 \add_98_4/U26  ( .A1(\add_98_4/n159 ), .A2(\add_98_4/n162 ), .ZN(
        \add_98_4/n25 ) );
  OR2_X4 \add_98_4/U25  ( .A1(\add_98_4/n310 ), .A2(\add_98_4/n329 ), .ZN(
        \add_98_4/n24 ) );
  AND2_X4 \add_98_4/U24  ( .A1(\add_98_4/n127 ), .A2(\add_98_4/n196 ), .ZN(
        \add_98_4/n23 ) );
  OR2_X4 \add_98_4/U23  ( .A1(\add_98_4/n309 ), .A2(\add_98_4/n310 ), .ZN(
        \add_98_4/n22 ) );
  AND2_X4 \add_98_4/U22  ( .A1(\add_98_4/n149 ), .A2(\add_98_4/n104 ), .ZN(
        \add_98_4/n21 ) );
  AND2_X4 \add_98_4/U21  ( .A1(\add_98_4/n109 ), .A2(\add_98_4/n110 ), .ZN(
        \add_98_4/n20 ) );
  AND2_X4 \add_98_4/U20  ( .A1(\add_98_4/n373 ), .A2(\add_98_4/n3 ), .ZN(
        \add_98_4/n19 ) );
  AND3_X4 \add_98_4/U19  ( .A1(\add_98_4/n31 ), .A2(\add_98_4/n150 ), .A3(
        \add_98_4/n163 ), .ZN(\add_98_4/n18 ) );
  OR2_X4 \add_98_4/U18  ( .A1(\add_98_4/n235 ), .A2(\add_98_4/n229 ), .ZN(
        \add_98_4/n17 ) );
  AND2_X4 \add_98_4/U17  ( .A1(rnd_q[47]), .A2(cv_q[47]), .ZN(\add_98_4/n16 )
         );
  OR2_X4 \add_98_4/U16  ( .A1(\add_98_4/n352 ), .A2(\add_98_4/n353 ), .ZN(
        \add_98_4/n15 ) );
  AND2_X4 \add_98_4/U15  ( .A1(\add_98_4/n215 ), .A2(\add_98_4/n341 ), .ZN(
        \add_98_4/n14 ) );
  AND2_X4 \add_98_4/U14  ( .A1(\add_98_4/n103 ), .A2(\add_98_4/n104 ), .ZN(
        \add_98_4/n13 ) );
  AND3_X4 \add_98_4/U13  ( .A1(\add_98_4/n103 ), .A2(\add_98_4/n94 ), .A3(
        \add_98_4/n104 ), .ZN(\add_98_4/n12 ) );
  AND2_X4 \add_98_4/U12  ( .A1(\add_98_4/n153 ), .A2(\add_98_4/n151 ), .ZN(
        \add_98_4/n11 ) );
  OR2_X4 \add_98_4/U11  ( .A1(cv_q[46]), .A2(rnd_q[46]), .ZN(\add_98_4/n10 )
         );
  OR2_X4 \add_98_4/U10  ( .A1(\add_98_4/n178 ), .A2(\add_98_4/n179 ), .ZN(
        \add_98_4/n9 ) );
  OR2_X4 \add_98_4/U9  ( .A1(cv_q[33]), .A2(rnd_q[33]), .ZN(\add_98_4/n8 ) );
  OR3_X4 \add_98_4/U8  ( .A1(\add_98_4/n327 ), .A2(\add_98_4/n19 ), .A3(
        \add_98_4/n328 ), .ZN(\add_98_4/n7 ) );
  OR2_X4 \add_98_4/U7  ( .A1(cv_q[38]), .A2(rnd_q[38]), .ZN(\add_98_4/n6 ) );
  OR2_X4 \add_98_4/U6  ( .A1(cv_q[35]), .A2(rnd_q[35]), .ZN(\add_98_4/n5 ) );
  OR2_X4 \add_98_4/U5  ( .A1(cv_q[45]), .A2(rnd_q[45]), .ZN(\add_98_4/n4 ) );
  OR2_X4 \add_98_4/U4  ( .A1(cv_q[39]), .A2(rnd_q[39]), .ZN(\add_98_4/n3 ) );
  OR2_X4 \add_98_4/U3  ( .A1(cv_q[34]), .A2(rnd_q[34]), .ZN(\add_98_4/n2 ) );
  AND3_X4 \add_98_4/U2  ( .A1(\add_98_4/n2 ), .A2(\add_98_4/n5 ), .A3(
        \add_98_4/n8 ), .ZN(\add_98_4/n1 ) );
endmodule

