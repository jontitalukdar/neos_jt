module s5378(blif_clk_net, blif_reset_net, n3065gat, n3066gat,n3067gat, n3068gat, n3069gat, n3070gat, n3071gat, n3072gat,n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat,n3079gat, n3080gat, n3081gat, n3082gat, n3083gat, n3084gat,n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat,n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat,n3098gat, n3099gat, n3100gat, n3104gat, n3105gat, n3106gat,n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat,n3113gat, n3114gat, n3115gat, n3116gat, n3117gat, n3118gat,n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat,n3131gat, n3132gat, n3133gat, n3134gat, n3135gat, n3136gat,n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat,n3143gat, n3144gat, n3145gat, n3146gat, n3147gat, n3148gat,n3149gat, n3150gat, n3151gat, n3152gat);
input blif_clk_net, blif_reset_net, n3065gat, n3066gat, n3067gat,n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat,n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat,n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat,n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat,n3099gat, n3100gat;
output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat,n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat,n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat,n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat,n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat,n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat,n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat,n3152gat;
wire blif_clk_net, blif_reset_net, n3065gat, n3066gat, n3067gat,n3068gat, n3069gat, n3070gat, n3071gat, n3072gat, n3073gat,n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat,n3080gat, n3081gat, n3082gat, n3083gat, n3084gat, n3085gat,n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, n3091gat,n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat,n3099gat, n3100gat;
wire n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat,n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, n3115gat,n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat,n3122gat, n3123gat, n3124gat, n3125gat, n3126gat, n3127gat,n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat,n3134gat, n3135gat, n3136gat, n3137gat, n3138gat, n3139gat,n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat,n3152gat;
wire n148gat, n152gat, n156gat, n160gat, n256gat, n271gat, n314gat,n322gat;
wire n327gat, n331gat, n337gat, n341gat, n366gat, n384gat, n388gat,n398gat;
wire n402gat, n463gat, n470gat, n553gat, n561gat, n580gat, n584gat,n614gat;
wire n659gat, n667gat, n673gat, n680gat, n684gat, n699gat, n707gat,n777gat;
wire n816gat, n820gat, n824gat, n830gat, n834gat, n838gat, n842gat,n861gat;
wire n865gat, n883gat, n919gat, n931gat, n957gat, n1035gat, n1045gat,n1068gat;
wire n1072gat, n1080gat, n1121gat, n1135gat, n1148gat, n1197gat,n1226gat, n1241gat;
wire n1282gat, n1294gat, n1312gat, n1316gat, n1332gat, n1336gat,n1340gat, n1363gat;
wire n1389gat, n1394gat, n1433gat, n1456gat, n1462gat, n1496gat,n1508gat, n1525gat;
wire n1588gat, n1596gat, n1675gat, n1678gat, n1740gat, n1748gat,n1763gat, n1767gat;
wire n1771gat, n1775gat, n1807gat, n1821gat, n1829gat, n1834gat,n1850gat, n1871gat;
wire n1880gat, n1899gat, n1975gat, n2021gat, n2025gat, n2029gat,n2033gat, n2037gat;
wire n2040gat, n2044gat, n2084gat, n2091gat, n2095gat, n2099gat,n2102gat, n2110gat;
wire n2117gat, n2121gat, n2125gat, n2135gat, n2155gat, n2169gat,n2176gat, n2179gat;
wire n2182gat, n2190gat, n2203gat, n2207gat, n2262gat, n2266gat,n2319gat, n2343gat;
wire n2347gat, n2394gat, n2399gat, n2403gat, n2407gat, n2440gat,n2446gat, n2450gat;
wire n2454gat, n2458gat, n2464gat, n2468gat, n2472gat, n2476gat,n2490gat, n2495gat;
wire n2502gat, n2506gat, n2510gat, n2514gat, n2518gat, n2522gat,n2526gat, n2543gat;
wire n2562gat, n2588gat, n2592gat, n2599gat, n2622gat, n2626gat,n2630gat, n2634gat;
wire n2640gat, n2644gat, n2658gat, n_0, n_1, n_2, n_3, n_4;
wire n_5, n_8, n_9, n_10, n_12, n_13, n_15, n_18;
wire n_20, n_21, n_23, n_26, n_27, n_31, n_36, n_38;
wire n_42, n_44, n_46, n_50, n_51, n_54, n_55, n_63;
wire n_65, n_66, n_72, n_73, n_74, n_75, n_80, n_83;
wire n_85, n_90, n_95, n_96, n_100, n_106, n_111, n_116;
wire n_117, n_121, n_122, n_129, n_130, n_131, n_132, n_135;
wire n_136, n_140, n_141, n_142, n_143, n_145, n_153, n_154;
wire n_156, n_157, n_158, n_159, n_162, n_164, n_165, n_167;
wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_177;
wire n_185, n_194, n_195, n_196, n_197, n_198, n_199, n_202;
wire n_203, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
wire n_213, n_215, n_217, n_218, n_219, n_220, n_221, n_226;
wire n_227, n_228, n_229, n_231, n_235, n_237, n_238, n_239;
wire n_240, n_241, n_242, n_243, n_244, n_248, n_249, n_251;
wire n_252, n_253, n_254, n_256, n_257, n_258, n_259, n_260;
wire n_261, n_262, n_266, n_268, n_269, n_270, n_271, n_273;
wire n_274, n_277, n_278, n_279, n_281, n_282, n_287, n_289;
wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_302;
wire n_303, n_306, n_310, n_311, n_312, n_313, n_314, n_315;
wire n_316, n_318, n_319, n_320, n_322, n_324, n_325, n_326;
wire n_328, n_329, n_330, n_333, n_335, n_336, n_338, n_339;
wire n_342, n_343, n_344, n_347, n_350, n_351, n_355, n_356;
wire n_357, n_364, n_365, n_366, n_367, n_369, n_374, n_375;
wire n_376, n_377, n_378, n_380, n_381, n_382, n_384, n_385;
wire n_386, n_387, n_388, n_389, n_390, n_391, n_395, n_396;
wire n_397, n_398, n_400, n_401, n_402, n_403, n_404, n_405;
wire n_406, n_407, n_409, n_410, n_411, n_412, n_413, n_414;
wire n_415, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
wire n_426, n_427, n_428, n_431, n_432, n_435, n_436, n_437;
wire n_442, n_444, n_447, n_448, n_451, n_452, n_454, n_455;
wire n_457, n_458, n_461, n_462, n_463, n_464, n_466, n_467;
wire n_468, n_475, n_476, n_479, n_481, n_482, n_483, n_484;
wire n_487, n_489, n_490, n_491, n_493, n_494, n_495, n_496;
wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
wire n_506, n_511, n_515, n_518, n_519, n_521, n_522, n_523;
wire n_524, n_527, n_529, n_530, n_531, n_532, n_533, n_535;
wire n_536, n_537, n_547, n_549, n_553, n_554, n_555, n_556;
wire n_557, n_558, n_560, n_561, n_562, n_563, n_565, n_566;
wire n_567, n_568, n_569, n_570, n_573, n_574, n_575, n_578;
wire n_579, n_580, n_581, n_584, n_585, n_586, n_587, n_588;
wire n_590, n_591, n_592, n_593, n_595, n_597, n_598, n_600;
wire n_602, n_603, n_604, n_610, n_611, n_612, n_613, n_614;
wire n_615, n_616, n_617, n_619, n_620, n_621, n_622, n_623;
wire n_627, n_630, n_631, n_632, n_633, n_634, n_637, n_638;
wire n_639, n_642, n_643, n_644, n_645, n_646, n_648, n_649;
wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
wire n_659, n_660, n_661, n_667, n_671, n_676, n_679, n_680;
wire n_681, n_683, n_684, n_685, n_687, n_689, n_690, n_691;
wire n_694, n_696, n_697, n_699, n_700, n_701, n_703, n_704;
wire n_705, n_706, n_708, n_714, n_716, n_719, n_720, n_722;
wire n_723, n_724, n_725, n_726, n_728, n_730, n_731, n_732;
wire n_733, n_736, n_738, n_739, n_743, n_744, n_747, n_748;
wire n_749, n_750, n_751, n_755, n_756, n_757, n_758, n_760;
wire n_761, n_763, n_764, n_766, n_767, n_769, n_770, n_771;
wire n_772, n_774, n_775, n_776, n_777, n_778, n_779, n_781;
wire n_782, n_786, n_787, n_788, n_789, n_791, n_795, n_796;
wire n_798, n_800, n_802, n_805, n_806, n_807, n_808, n_809;
wire n_812, n_813, n_815, n_816, n_817, n_819, n_820, n_821;
wire n_822, n_823, n_824, n_829, n_830, n_831, n_832, n_833;
wire n_834, n_835, n_836, n_840, n_841, n_842, n_852, n_854;
wire n_855, n_856, n_857, n_859, n_860, n_861, n_862, n_863;
wire n_864, n_866, n_867, n_868, n_870, n_872, n_876, n_877;
wire n_878, n_879, n_880, n_882, n_883, n_884, n_885, n_887;
wire n_888, n_889, n_892, n_894, n_901, n_902, n_903, n_904;
wire n_905, n_906, n_908, n_909, n_911, n_913, n_914, n_915;
wire n_917, n_918, n_919, n_920, n_921, n_922, n_924, n_925;
wire n_926, n_928, n_929, n_930, n_931, n_936, n_937, n_938;
wire n_939, n_940, n_941, n_943, n_944, n_948, n_950, n_951;
wire n_952, n_953, n_954, n_955, n_956, n_957, n_959, n_961;
wire n_963, n_965, n_966, n_967, n_968, n_970, n_971, n_972;
wire n_973, n_976, n_979, n_980, n_981, n_982, n_984, n_985;
wire n_987, n_988, n_989, n_990, n_993, n_994, n_997, n_998;
wire n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1006, n_1009;
wire n_1010, n_1011, n_1014, n_1017, n_1019, n_1020, n_1021, n_1023;
wire n_1024, n_1026, n_1027, n_1030, n_1033, n_1034, n_1036, n_1037;
wire n_1038, n_1039, n_1040, n_1041, n_1044, n_1045, n_1046, n_1047;
wire n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056;
wire n_1057, n_1058, n_1060, n_1061, n_1062, n_1063, n_1064, n_1066;
wire n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075;
wire n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1084;
wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
wire n_1094, n_1095, n_1096, n_1097, n_1099, n_1100, n_1101, n_1103;
wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
wire n_1132, n_1133, n_1140, n_1147, n_1148, n_1149, n_1150, n_1151;
wire n_1153, n_1154, n_1155, n_1158, n_1159, n_1160, n_1161, n_1164;
wire n_1165, n_1167, n_1168, n_1169, n_1170, n_1171, n_1191, n_1196;
wire n_1197, n_1198, n_1201, n_1208, n_1211, n_1216, n_1241, n_1245;
wire n_1253, n_1259, n_1262, n_1267, n_1268, n_1269, n_1272, n_1275;
wire n_1276, n_1277, n_1282, n_1283, n_1289, n_1294, n_1295, n_1310;
wire n_1326, n_1337, n_1338, n_1339, n_1342, n_1343, n_1344, n_1345;
wire n_1354, n_1362, n_1363, n_1366, n_1371, n_1373, n_1376, n_1377;
wire n_1378, n_1380, n_1381, n_1382, n_1396, n_1397, n_1398, n_1399;
wire n_1402, n_1419, n_1420, n_1421, n_1430, n_1431, n_1442, n_1443;
wire n_1453, n_1464, n_1483, n_1485, n_1486, n_1493, n_1494, n_1497;
wire n_1498, n_1504, n_1505, n_1506, n_1508, n_1510, n_1513, n_1514;
wire n_1515, n_1525, n_1526, n_1527, n_1528, n_1531, n_1544, n_1546;
wire n_1547, n_1548, n_1550, n_1551, n_1552, n_1559, n_1562, n_1566;
wire n_1571, n_1573, n_1577, n_1580, n_1581, n_1588, n_1589, n_1590;
wire n_1591, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599;
wire n_1600, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613;
wire n_1621, n_1637, n_1646, n_1647, n_1648, n_1650, n_1651, n_1652;
wire n_1653, n_1658, n_1659, n_1660, n_1661, n_1664, n_1668, n_1669;
wire n_1670, n_1680, n_1683, n_1684, n_1685, n_1686, n_1687, n_1697;
wire n_1698, n_1699, n_1702, n_1707, n_1708, n_1715, n_1718, n_1719;
wire n_1720, n_1721, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729;
wire n_1730, n_1731, n_1732, n_1733, n_1734, n_1748, n_1749, n_1751;
wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
wire n_1761, n_1766, n_1770, n_1771, n_1774, n_1775, n_1776, n_1777;
wire n_1779, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790;
wire n_1792, n_1793, n_1794, n_1796, n_1797, n_1798, n_1799, n_1800;
wire n_1801, n_1802, n_1803, n_1807, n_1808, n_1809, n_1810, n_1811;
wire n_1812, n_1814, n_1816, n_1818, n_1819, n_1821, n_1823, n_1824;
wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1834, n_1837;
wire n_1842, n_1843, n_1851, n_1852, n_1857, n_1859, n_1860, n_1862;
wire n_1864, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1877;
wire n_1878, n_1881, n_1882, n_1884, n_1885, n_1886, n_1887, n_1888;
wire n_1889, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1898;
wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
wire n_1909, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918;
wire n_1919, n_1920, n_1922, n_1923, n_1924, n_1926, n_1927, n_1928;
wire n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936;
wire n_1937, n_1938, n_1939, n_1947, n_1948, n_1949, n_1950, n_1951;
wire n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964;
wire n_1965, n_1966, n_1967, n_1981, n_1984, n_1990, n_1992, n_1994;
wire n_1995, n_2002, n_2003, n_2004, n_2007, n_2008, n_2014, n_2015;
wire n_2019, n_2021, n_2022, n_2024, n_2027, n_2029, n_2030, n_2031;
wire n_2032, n_2033, n_2035, n_2041, n_2042, n_2043, n_2044, n_2046;
wire n_2048, n_2049, n_2050, n_2051, n_2055, n_2056, n_2059, n_2063;
wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
wire n_2072, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080;
wire n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089;
wire n_2090, n_2091, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098;
wire n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2106, n_2107;
wire n_2108, n_2109, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
wire n_2120, n_2121;
assign n3152gat = 1'b1;
assign n3142gat = n3141gat;
assign n3140gat = n3139gat;
assign n3115gat = 1'b1;
assign n3112gat = 1'b1;
OR2X1 g6944(.A (n_2109), .B (n_592), .Y (n3143gat));
OR2X1 g6945(.A (n_2109), .B (n_621), .Y (n3144gat));
DFFSRX1 n2588gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1170), .Q (n2588gat), .QN ());
NAND2X1 g6950(.A (n_1169), .B (n_1019), .Y (n3125gat));
INVX1 g6951(.A (n_1171), .Y (n3129gat));
AOI21X1 g6952(.A0 (n_1168), .A1 (n_1125), .B0 (n_1155), .Y (n_1171));
OR4X1 g6953(.A (n_1160), .B (n2464gat), .C (n3090gat), .D (n2599gat),.Y (n_1170));
NAND2X1 g6954(.A (n_1168), .B (n_1120), .Y (n_1169));
NAND3X1 g6955(.A (n_2114), .B (n_2115), .C (n_1080), .Y (n_1167));
NAND3X1 g6956(.A (n_556), .B (n_570), .C (n_1161), .Y (n_1168));
NAND2X1 g6958(.A (n_1109), .B (n_1164), .Y (n3123gat));
DFFSRX1 n2599gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1164), .Q (), .QN (n2599gat));
XOR2X1 g6961(.A (n667gat), .B (n_1938), .Y (n_1164));
XOR2X1 g6962(.A (n_574), .B (n_1938), .Y (n_2114));
AOI22X1 g6960(.A0 (n_1939), .A1 (n_1075), .B0 (n842gat), .B1(n_1071), .Y (n_1161));
NAND4X1 g6959(.A (n_1159), .B (n2476gat), .C (n2468gat), .D(n2526gat), .Y (n_1160));
NOR2X1 g6963(.A (n2518gat), .B (n2522gat), .Y (n_1159));
NAND2X1 g6971(.A (n_1153), .B (n_1132), .Y (n_1158));
NAND2X1 g6966(.A (n_1107), .B (n_2082), .Y (n3124gat));
DFFSRX1 n2518gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_2082), .Q (), .QN (n2518gat));
AOI21X1 g6965(.A0 (n_1148), .A1 (n_557), .B0 (n_1140), .Y (n_1155));
NAND2X1 g6968(.A (n_1151), .B (n_1133), .Y (n_1154));
OAI21X1 g6974(.A0 (n_1149), .A1 (n_1150), .B0 (n_1147), .Y (n_1153));
XOR2X1 g6972(.A (n_1150), .B (n_1149), .Y (n_1151));
NAND2X1 g6970(.A (n3116gat), .B (n_1075), .Y (n_1148));
NAND2X1 g6975(.A (n_1149), .B (n_1150), .Y (n_1147));
NAND2X2 g6977(.A (n_1127), .B (n_1097), .Y (n_1149));
NAND2X1 g6983(.A (n_1115), .B (n_1039), .Y (n3121gat));
NAND2X1 g6984(.A (n_1113), .B (n_973), .Y (n3122gat));
NAND2X1 g6981(.A (n_1122), .B (n_691), .Y (n3117gat));
NAND2X1 g6985(.A (n_1111), .B (n_1613), .Y (n3118gat));
NAND2X1 g6986(.A (n_1105), .B (n_821), .Y (n3119gat));
OAI21X1 g6991(.A0 (n_642), .A1 (n_1140), .B0 (n_1126), .Y (n3130gat));
OAI21X1 g6987(.A0 (n_1040), .A1 (n_1140), .B0 (n_1124), .Y(n3131gat));
OAI21X1 g6988(.A0 (n_1038), .A1 (n_1140), .B0 (n_1123), .Y(n3132gat));
OAI21X1 g6992(.A0 (n_1000), .A1 (n_1140), .B0 (n_1119), .Y(n3134gat));
OAI21X1 g6993(.A0 (n_999), .A1 (n_1140), .B0 (n_1118), .Y (n3135gat));
OAI21X1 g6994(.A0 (n_997), .A1 (n_1140), .B0 (n_1117), .Y (n3136gat));
OAI21X1 g6990(.A0 (n_994), .A1 (n_1140), .B0 (n_1116), .Y (n3137gat));
INVX1 g6978(.A (n_1132), .Y (n_1133));
NAND2X1 g6982(.A (n_1100), .B (n_1613), .Y (n3120gat));
OAI21X1 g6989(.A0 (n_1036), .A1 (n_1140), .B0 (n_1101), .Y(n3133gat));
NAND4X1 g7072(.A (n_1047), .B (n_761), .C (n_733), .D (n_1086), .Y(n3141gat));
AND2X1 g7239(.A (n_1103), .B (n_771), .Y (n3146gat));
AOI21X1 g6979(.A0 (n_1060), .A1 (n314gat), .B0 (n_1095), .Y (n_1132));
NAND4X1 g7225(.A (n_889), .B (n_1090), .C (n_758), .D (n_747), .Y(n3139gat));
NAND2X1 g6980(.A (n_1094), .B (n659gat), .Y (n_1127));
NAND2X1 g6996(.A (n_1121), .B (n_1125), .Y (n_1126));
NAND2X1 g6997(.A (n_1110), .B (n_1125), .Y (n_1124));
NAND2X1 g6998(.A (n_1104), .B (n_1125), .Y (n_1123));
NAND2X1 g6999(.A (n_1121), .B (n_1120), .Y (n_1122));
NAND2X1 g7001(.A (n_1114), .B (n_1125), .Y (n_1119));
NAND2X1 g7002(.A (n_1112), .B (n_1125), .Y (n_1118));
NAND2X1 g7003(.A (n_1108), .B (n_1125), .Y (n_1117));
NAND2X1 g7004(.A (n_1125), .B (n_1106), .Y (n_1116));
NAND2X1 g7006(.A (n_1114), .B (n_1120), .Y (n_1115));
NAND2X1 g7007(.A (n_1112), .B (n_1120), .Y (n_1113));
NAND2X1 g7008(.A (n_1110), .B (n_1120), .Y (n_1111));
NAND2X1 g7009(.A (n_1108), .B (n_1120), .Y (n_1109));
NAND2X1 g7010(.A (n_1106), .B (n_1120), .Y (n_1107));
NAND2X1 g7011(.A (n_1104), .B (n_1120), .Y (n_1105));
NOR2X1 g7251(.A (n_1087), .B (n2033gat), .Y (n_1103));
NAND2X1 g7000(.A (n_1099), .B (n_1125), .Y (n_1101));
NAND2X1 g7005(.A (n_1099), .B (n_1120), .Y (n_1100));
NAND2X1 g7014(.A (n_1085), .B (n_1079), .Y (n_1097));
NAND2X1 g7024(.A (n_530), .B (n_1066), .Y (n_1110));
OR2X1 g7025(.A (n_1077), .B (n_1088), .Y (n_1096));
NAND2X1 g7026(.A (n_862), .B (n_1064), .Y (n_1108));
DFFSRX1 n1316gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n1433gat), .Q (n1316gat), .QN ());
AOI21X1 g7015(.A0 (n_1045), .A1 (n_1049), .B0 (n314gat), .Y (n_1095));
NAND2X1 g7016(.A (n_1061), .B (n_1052), .Y (n_1094));
NAND3X1 g7018(.A (n_602), .B (n_1053), .C (n_817), .Y (n_1106));
NAND2X1 g7019(.A (n_553), .B (n_1076), .Y (n_1114));
NAND2X1 g7020(.A (n_555), .B (n_1074), .Y (n_1104));
NAND2X1 g7021(.A (n_802), .B (n_1072), .Y (n_1121));
NAND2X1 g7023(.A (n_532), .B (n_1070), .Y (n_1112));
AND2X1 g7263(.A (n_1058), .B (n_774), .Y (n_1090));
OR2X1 g7029(.A (n_1054), .B (n_1088), .Y (n_1089));
NAND4X1 g7274(.A (n_1057), .B (n2110gat), .C (n2176gat), .D(n2037gat), .Y (n_1087));
OAI21X1 g7135(.A0 (n_763), .A1 (n_867), .B0 (n1456gat), .Y (n_1086));
NAND2X1 g7042(.A (n_1051), .B (n_1050), .Y (n_1085));
NAND2X1 g7012(.A (n_1091), .B (n_1092), .Y (n_1084));
NAND2X1 g7022(.A (n_770), .B (n_1055), .Y (n_1099));
DFFSRX1 n1871gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1046), .Q (n1871gat), .QN ());
AOI21X1 g7303(.A0 (n2514gat), .A1 (n_1017), .B0 (n_724), .Y(n3145gat));
NAND3X1 g7030(.A (n_287), .B (n_854), .C (n_1062), .Y (n_1082));
AOI22X1 g7032(.A0 (n_1080), .A1 (n_1079), .B0 (n_833), .B1 (n322gat),.Y (n_1081));
AOI22X1 g7033(.A0 (n_377), .A1 (n_1073), .B0 (n_856), .B1 (n_1990),.Y (n_1078));
AOI22X1 g7034(.A0 (n_829), .A1 (n_1063), .B0 (n_835), .B1 (n_1068),.Y (n_1077));
AOI21X1 g7035(.A0 (n_1030), .A1 (n_1075), .B0 (n_494), .Y (n_1076));
AOI22X1 g7036(.A0 (n_1069), .A1 (n816gat), .B0 (n_1073), .B1(n_1075), .Y (n_1074));
AOI22X1 g7037(.A0 (n_1075), .A1 (n_1079), .B0 (n_1071), .B1(n271gat), .Y (n_1072));
AOI22X1 g7039(.A0 (n_1069), .A1 (n684gat), .B0 (n_1068), .B1(n_1075), .Y (n_1070));
AOI22X1 g7040(.A0 (n_1069), .A1 (n580gat), .B0 (n_1990), .B1(n_1075), .Y (n_1066));
AOI22X1 g7041(.A0 (n_1063), .A1 (n_1075), .B0 (n_2007), .B1 (n_1071),.Y (n_1064));
XOR2X1 g7043(.A (n_1062), .B (n_1063), .Y (n_1150));
NAND2X1 g7047(.A (n_1041), .B (n_1990), .Y (n_1061));
DFFSRX1 n1433gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1044), .Q (), .QN (n1433gat));
XOR2X1 g7017(.A (n_1068), .B (n322gat), .Y (n_1060));
MX2X1 g7027(.A (n_1004), .B (n_1020), .S0 (n1072gat), .Y (n_1091));
DFFSRX1 n2454gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1196), .Q (n2454gat), .QN ());
DFFSRX1 n2339gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1027), .Q (), .QN (n3126gat));
DFFSRX1 n2495gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1026), .Q (n2495gat), .QN ());
NAND4X1 g7293(.A (n1775gat), .B (n_1056), .C (n_15), .D (n_1006), .Y(n_1058));
NAND4X1 g7308(.A (n2514gat), .B (n1771gat), .C (n_1056), .D (n_931),.Y (n_1057));
DFFSRX1 n1456gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1197), .Q (), .QN (n1456gat));
AOI22X1 g7038(.A0 (n322gat), .A1 (n_1075), .B0 (n341gat), .B1(n_1071), .Y (n_1055));
NAND2X1 g7044(.A (n_1686), .B (n_1030), .Y (n_1054));
NAND2X1 g7045(.A (n_1062), .B (n_1075), .Y (n_1053));
NAND2X1 g7046(.A (n_1073), .B (n777gat), .Y (n_1052));
OR2X1 g7048(.A (n_1073), .B (n_1990), .Y (n_1051));
NAND2X1 g7049(.A (n_1073), .B (n_1990), .Y (n_1050));
NAND2X1 g7051(.A (n_1068), .B (n322gat), .Y (n_1049));
DFFSRX1 n2099gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2025gat), .Q (n2099gat), .QN ());
DFFSRX1 n2037gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2044gat), .Q (n2037gat), .QN ());
OR2X1 g7103(.A (n_1011), .B (n1135gat), .Y (n3113gat));
NAND2X1 g7102(.A (n_842), .B (n1748gat), .Y (n_1047));
INVX2 g7155(.A (n_1033), .Y (n_1046));
OR2X1 g7050(.A (n_1068), .B (n322gat), .Y (n_1045));
OAI33X1 g7180(.A0 (n_1003), .A1 (n_1779), .A2 (n_1295), .B0 (n_1779),.B1 (n_1295), .B2 (n2182gat), .Y (n_1044));
INVX1 g7053(.A (n_1073), .Y (n_1041));
AOI21X1 g7073(.A0 (n337gat), .A1 (n_1037), .B0 (n_1024), .Y (n_1040));
DFFSRX1 n2464gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1039), .Q (), .QN (n2464gat));
AOI21X1 g7074(.A0 (n_554), .A1 (n_1037), .B0 (n_1023), .Y (n_1038));
AOI21X1 g7075(.A0 (n341gat), .A1 (n_1037), .B0 (n_1021), .Y (n_1036));
AOI21X1 g7031(.A0 (n_988), .A1 (n_987), .B0 (n1045gat), .Y (n_1034));
DFFSRX1 n2514gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2458gat), .Q (n2514gat), .QN ());
NAND3X1 g7156(.A (n_1262), .B (n_1245), .C (n_1963), .Y (n_1033));
INVX2 g7054(.A (n553gat), .Y (n_1073));
INVX1 g7057(.A (n659gat), .Y (n_1079));
INVX1 g7059(.A (n314gat), .Y (n_1030));
INVX1 g7067(.A (n561gat), .Y (n_1063));
INVX1 g7069(.A (n366gat), .Y (n_1062));
NOR2X1 g7191(.A (n_1771), .B (n_1010), .Y (n_1027));
OR2X1 g7204(.A (n_1002), .B (n_1771), .Y (n_1026));
OAI21X1 g7089(.A0 (n_493), .A1 (n838gat), .B0 (n_993), .Y (n_1024));
OAI21X1 g7090(.A0 (n_493), .A1 (n707gat), .B0 (n_982), .Y (n_1023));
OAI21X1 g7091(.A0 (n_493), .A1 (n614gat), .B0 (n_990), .Y (n_1021));
OAI21X1 g7093(.A0 (n1121gat), .A1 (n1035gat), .B0 (n_989), .Y(n_1020));
DFFSRX1 n2502gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1019), .Q (n2502gat), .QN ());
DFFSRX1 n2270gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_968), .Q (), .QN (n3127gat));
NOR2X1 g7358(.A (n_1017), .B (n3106gat), .Y (n3107gat));
DFFSRX1 n2044gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_985), .Q (), .QN (n2044gat));
DFFSRX1 n2025gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1191), .Q (), .QN (n2025gat));
DFFSRX1 n1748gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_984), .Q (), .QN (n1748gat));
NAND3X1 g7161(.A (n_1607), .B (n_1531), .C (n_401), .Y (n_1014));
DFFSRX1 n553gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1653), .Q (n553gat), .QN ());
DFFSRX1 n322gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1720), .Q (), .QN (n322gat));
DFFSRX1 n659gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_971), .Q (n659gat), .QN ());
DFFSRX1 n314gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_980), .Q (n314gat), .QN ());
DFFSRX1 n318gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_979), .Q (), .QN (n_1068));
DFFSRX1 n777gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1829), .Q (n777gat), .QN ());
DFFSRX1 n561gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_972), .Q (n561gat), .QN ());
DFFSRX1 n366gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_976), .Q (n366gat), .QN ());
DFFSRX1 n667gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_970), .Q (), .QN (n667gat));
MX2X1 g7209(.A (n_957), .B (n_965), .S0 (n_879), .Y (n_1039));
INVX1 g7210(.A (n_1010), .Y (n_1011));
XOR2X1 g7092(.A (n931gat), .B (n1135gat), .Y (n_1009));
XOR2X1 g7094(.A (n1226gat), .B (n1282gat), .Y (n_1092));
OR2X1 g7104(.A (n_967), .B (n1282gat), .Y (n3114gat));
AOI21X1 g7313(.A0 (n_961), .A1 (n1821gat), .B0 (n_831), .Y (n_1006));
DFFSRX1 n2458gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2592gat), .Q (), .QN (n2458gat));
XOR2X1 g7052(.A (n1035gat), .B (n1121gat), .Y (n_1004));
NAND3X1 g7195(.A (n2179gat), .B (n_1001), .C (n_162), .Y (n_1003));
XOR2X1 g7227(.A (n2266gat), .B (n_963), .Y (n_1002));
XOR2X1 g7228(.A (n2135gat), .B (n_1001), .Y (n_1010));
AOI22X1 g7085(.A0 (n_998), .A1 (n_2035), .B0 (n_1075), .B1(n1045gat), .Y (n_1000));
AOI22X1 g7086(.A0 (n_998), .A1 (n_531), .B0 (n_1075), .B1 (n1135gat),.Y (n_999));
AOI22X1 g7087(.A0 (n_998), .A1 (n_2007), .B0 (n_1075), .B1(n1282gat), .Y (n_997));
AOI22X1 g7088(.A0 (n_998), .A1 (n_600), .B0 (n_1075), .B1 (n1226gat),.Y (n_994));
NAND2X1 g7096(.A (n_1075), .B (n1072gat), .Y (n_993));
OR2X1 g7099(.A (n_914), .B (n1072gat), .Y (n3109gat));
NAND2X1 g7101(.A (n_929), .B (n1121gat), .Y (n3110gat));
OR2X1 g7098(.A (n_981), .B (n931gat), .Y (n_990));
NAND2X1 g7100(.A (n1121gat), .B (n1035gat), .Y (n_989));
OR2X1 g7105(.A (n1135gat), .B (n931gat), .Y (n_988));
NAND2X1 g7106(.A (n1135gat), .B (n931gat), .Y (n_987));
NAND2X1 g7095(.A (n_1646), .B (n931gat), .Y (n3111gat));
AND2X1 g7356(.A (n_959), .B (n2040gat), .Y (n_985));
AND2X1 g7383(.A (n1771gat), .B (n_931), .Y (n_1017));
NOR2X1 g7174(.A (n_1967), .B (n_1373), .Y (n_984));
OR2X1 g7097(.A (n_981), .B (n1121gat), .Y (n_982));
NAND3X1 g7076(.A (n_1830), .B (n_952), .C (n_951), .Y (n_980));
NAND3X1 g7077(.A (n_1830), .B (n_950), .C (n_948), .Y (n_979));
NAND3X1 g7079(.A (n_1830), .B (n_944), .C (n_943), .Y (n_976));
DFFSRX1 n2526gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_973), .Q (n2526gat), .QN ());
NAND3X1 g7081(.A (n_1830), .B (n_941), .C (n_940), .Y (n_972));
NAND3X1 g7082(.A (n_1830), .B (n_939), .C (n_938), .Y (n_971));
XOR2X1 g7229(.A (n_954), .B (n_140), .Y (n_1019));
NAND3X1 g7083(.A (n_1830), .B (n_937), .C (n_936), .Y (n_970));
NOR2X1 g7233(.A (n_1771), .B (n_966), .Y (n_968));
INVX1 g7255(.A (n_966), .Y (n_967));
OAI21X1 g7276(.A0 (n_955), .A1 (n_956), .B0 (n_953), .Y (n_965));
DFFSRX1 n2592gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n1775gat), .Q (), .QN (n2592gat));
NOR2X1 g7254(.A (n2262gat), .B (n2190gat), .Y (n_1001));
AND2X1 g7256(.A (n2262gat), .B (n2190gat), .Y (n_966));
NOR2X1 g7257(.A (n2262gat), .B (n_27), .Y (n_963));
DFFSRX1 n1035gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_925), .Q (n1035gat), .QN ());
DFFSRX1 n2343gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_928), .Q (n2343gat), .QN ());
DFFSRX1 n2399gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_930), .Q (n2399gat), .QN ());
DFFSRX1 n1121gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_921), .Q (n1121gat), .QN ());
DFFSRX1 n931gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_926), .Q (n931gat), .QN ());
DFFSRX1 n1072gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_922), .Q (), .QN (n1072gat));
DFFSRX1 n1282gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_917), .Q (), .QN (n1282gat));
DFFSRX1 n1135gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_920), .Q (), .QN (n1135gat));
DFFSRX1 n1226gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_918), .Q (), .QN (n1226gat));
DFFSRX1 n1197gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_919), .Q (), .QN (n1197gat));
DFFSRX1 n1045gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_924), .Q (), .QN (n1045gat));
NAND3X1 g7357(.A (n3097gat), .B (n_1259), .C (n1775gat), .Y (n_961));
NOR2X1 g7379(.A (n1316gat), .B (n_931), .Y (n_959));
MX2X1 g7241(.A (n_911), .B (n_902), .S0 (n_622), .Y (n_973));
XOR2X1 g7242(.A (n_956), .B (n_955), .Y (n_957));
XOR2X1 g7260(.A (n2495gat), .B (n3128gat), .Y (n_954));
DFFSRX1 n2630gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_904), .Q (n2630gat), .QN ());
DFFSRX1 n2622gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_905), .Q (n2622gat), .QN ());
DFFSRX1 n2490gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_908), .Q (n2490gat), .QN ());
DFFSRX1 n2207gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_913), .Q (n2207gat), .QN ());
DFFSRX1 n2203gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_915), .Q (n2203gat), .QN ());
DFFSRX1 n2640gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_909), .Q (n2640gat), .QN ());
DFFSRX1 n2543gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_906), .Q (n2543gat), .QN ());
NAND2X1 g7288(.A (n_955), .B (n_956), .Y (n_953));
NAND2X1 g7117(.A (n3069gat), .B (n_1651), .Y (n_952));
NAND2X1 g7118(.A (n3078gat), .B (n_1824), .Y (n_951));
NAND2X1 g7119(.A (n3070gat), .B (n_1651), .Y (n_950));
NAND2X1 g7120(.A (n3079gat), .B (n_1824), .Y (n_948));
NAND2X1 g7123(.A (n_1651), .B (n3072gat), .Y (n_944));
NAND2X1 g7124(.A (n_1824), .B (n3081gat), .Y (n_943));
NAND2X1 g7126(.A (n_1651), .B (n3071gat), .Y (n_941));
NAND2X1 g7127(.A (n_1824), .B (n3080gat), .Y (n_940));
NAND2X1 g7128(.A (n_1651), .B (n3065gat), .Y (n_939));
NAND2X1 g7129(.A (n3074gat), .B (n_1824), .Y (n_938));
NAND2X1 g7130(.A (n_1651), .B (n3073gat), .Y (n_937));
NAND2X1 g7131(.A (n_1824), .B (n3082gat), .Y (n_936));
OR2X1 g7382(.A (n1312gat), .B (n1775gat), .Y (n_1245));
DFFSRX1 n2634gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_903), .Q (n2634gat), .QN ());
DFFSRX1 n2262gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3128gat), .Q (n2262gat), .QN ());
NOR2X1 g7267(.A (n_929), .B (n_1992), .Y (n_930));
NOR2X1 g7268(.A (n_1646), .B (n_1992), .Y (n_928));
NAND2X1 g7146(.A (n_661), .B (n_1830), .Y (n_926));
NAND2X1 g7147(.A (n_660), .B (n_1830), .Y (n_925));
NAND2X1 g7148(.A (n_658), .B (n_1830), .Y (n_924));
NAND2X1 g7149(.A (n_657), .B (n_1830), .Y (n_922));
NAND2X1 g7150(.A (n_656), .B (n_1830), .Y (n_921));
NAND2X1 g7151(.A (n_655), .B (n_1830), .Y (n_920));
NAND2X1 g7152(.A (n_654), .B (n_1830), .Y (n_919));
NAND2X1 g7153(.A (n_653), .B (n_1830), .Y (n_918));
NAND2X1 g7154(.A (n_652), .B (n_1830), .Y (n_917));
INVX1 g7401(.A (n1775gat), .Y (n_931));
AND2X1 g7264(.A (n_914), .B (n_1995), .Y (n_915));
AND2X1 g7265(.A (n_380), .B (n_1995), .Y (n_913));
DFFSRX1 n1763gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_884), .Q (n1763gat), .QN ());
AOI21X1 g7309(.A0 (n_859), .A1 (n883gat), .B0 (n_887), .Y (n_955));
OAI21X1 g7310(.A0 (n_1790), .A1 (n_901), .B0 (n_888), .Y (n_911));
DFFSRX1 n1771gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_882), .Q (n1771gat), .QN ());
DFFSRX1 n1775gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_885), .Q (), .QN (n1775gat));
NAND2X1 g7266(.A (n_535), .B (n_1995), .Y (n_909));
DFFSRX1 n2626gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1802), .Q (n2626gat), .QN ());
AND2X1 g7234(.A (n_1802), .B (n_302), .Y (n_908));
AND2X1 g7235(.A (n_490), .B (n_1802), .Y (n_906));
AND2X1 g7236(.A (n_428), .B (n_1802), .Y (n_905));
AND2X1 g7237(.A (n_667), .B (n_1802), .Y (n_904));
NAND2X1 g7238(.A (n_529), .B (n_1802), .Y (n_903));
DFFSRX1 n2562gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1994), .Q (n2562gat), .QN ());
XOR2X1 g7277(.A (n_901), .B (n_1790), .Y (n_902));
DFFSRX1 n2390gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_880), .Q (), .QN (n3128gat));
AOI21X1 g7337(.A0 (n_270), .A1 (n_861), .B0 (n_877), .Y (n_894));
NOR2X1 g7404(.A (n_876), .B (n_870), .Y (n_892));
AOI22X1 g7259(.A0 (n_866), .A1 (n1508gat), .B0 (n_760), .B1(n1525gat), .Y (n_889));
NAND2X1 g7317(.A (n_1790), .B (n_901), .Y (n_888));
NOR2X1 g7322(.A (n_872), .B (n883gat), .Y (n_887));
NOR2X1 g7417(.A (n_632), .B (n_883), .Y (n_885));
NOR2X1 g7418(.A (n_883), .B (n_257), .Y (n_884));
NOR2X1 g7419(.A (n_883), .B (n_631), .Y (n_882));
INVX1 g7297(.A (n_1771), .Y (n_880));
AOI21X1 g7351(.A0 (n_820), .A1 (n699gat), .B0 (n_863), .Y (n_879));
AOI22X1 g7384(.A0 (n_364), .A1 (n_840), .B0 (n_375), .B1 (n_805), .Y(n_878));
NAND2X1 g7386(.A (n_855), .B (n_830), .Y (n_877));
NAND2X1 g7466(.A (n_852), .B (n_680), .Y (n_876));
MX2X1 g7352(.A (n_812), .B (n_808), .S0 (n838gat), .Y (n_901));
AOI21X1 g7353(.A0 (n824gat), .A1 (n820gat), .B0 (n_841), .Y (n_872));
OAI21X1 g7428(.A0 (n_366), .A1 (n_800), .B0 (n_1687), .Y (n_870));
OR2X1 g7437(.A (n_832), .B (n_603), .Y (n_883));
AOI21X1 g7275(.A0 (n1508gat), .A1 (n_867), .B0 (n_824), .Y (n_868));
NAND2X1 g7292(.A (n_764), .B (n_822), .Y (n_866));
AOI22X1 g7376(.A0 (n_378), .A1 (n_777), .B0 (n_365), .B1 (n_807), .Y(n_864));
NOR2X1 g7381(.A (n_813), .B (n699gat), .Y (n_863));
AOI22X1 g7385(.A0 (n_1069), .A1 (n824gat), .B0 (n_860), .B1 (n_1037),.Y (n_862));
AOI21X1 g7387(.A0 (n_778), .A1 (n580gat), .B0 (n_819), .Y (n_956));
MX2X1 g7388(.A (n824gat), .B (n_860), .S0 (n3149gat), .Y (n_861));
XOR2X1 g7390(.A (n820gat), .B (n824gat), .Y (n_859));
NAND3X1 g7406(.A (n_815), .B (n_376), .C (n_856), .Y (n_857));
NAND3X1 g7408(.A (n_816), .B (n_854), .C (n_1685), .Y (n_855));
NAND3X1 g7492(.A (n_809), .B (n_1080), .C (n_1685), .Y (n_852));
DFFSRX1 n152gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_779), .Q (n152gat), .QN ());
NAND3X1 g7136(.A (n_748), .B (n_823), .C (n_720), .Y (n_842));
NOR2X1 g7405(.A (n824gat), .B (n820gat), .Y (n_841));
AOI21X1 g7422(.A0 (n3149gat), .A1 (n160gat), .B0 (n_806), .Y (n_840));
NAND3X1 g7442(.A (n_798), .B (n_1685), .C (n_835), .Y (n_836));
NAND3X1 g7443(.A (n_796), .B (n_833), .C (n_1685), .Y (n_834));
DFFSRX1 n331gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n824gat), .Q (n331gat), .QN ());
OR2X1 g7460(.A (n2472gat), .B (n_831), .Y (n_832));
NAND3X1 g7484(.A (n_795), .B (n_829), .C (n_1685), .Y (n_830));
DFFSRX1 n699gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1733), .Q (n699gat), .QN ());
NOR2X1 g7316(.A (n_823), .B (n1678gat), .Y (n_824));
NAND2X1 g7321(.A (n_615), .B (n_867), .Y (n_822));
DFFSRX1 n2468gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_821), .Q (n2468gat), .QN ());
XOR2X1 g7391(.A (n584gat), .B (n684gat), .Y (n_820));
AOI21X1 g7407(.A0 (n_767), .A1 (n_766), .B0 (n580gat), .Y (n_819));
AOI22X1 g7421(.A0 (n_1069), .A1 (n883gat), .B0 (n673gat), .B1(n_1037), .Y (n_817));
MX2X1 g7423(.A (n684gat), .B (n1080gat), .S0 (n3149gat), .Y (n_816));
MX2X1 g7424(.A (n883gat), .B (n673gat), .S0 (n3149gat), .Y (n_815));
XOR2X1 g7426(.A (n584gat), .B (n684gat), .Y (n_813));
OAI21X1 g7427(.A0 (n834gat), .A1 (n707gat), .B0 (n_781), .Y (n_812));
NAND2X1 g7513(.A (n_519), .B (n2084gat), .Y (n_809));
DFFSRX1 n256gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_782), .Q (n256gat), .QN ());
DFFSRX1 n327gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n684gat), .Q (n327gat), .QN ());
XOR2X1 g7392(.A (n834gat), .B (n707gat), .Y (n_808));
DFFSRX1 n2476gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1613), .Q (n2476gat), .QN ());
DFFSRX1 n2522gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1613), .Q (), .QN (n2522gat));
OAI21X1 g7409(.A0 (n3149gat), .A1 (n838gat), .B0 (n_775), .Y (n_807));
DFFSRX1 n824gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_772), .Q (), .QN (n824gat));
NOR2X1 g7439(.A (n3149gat), .B (n_779), .Y (n_806));
OAI21X1 g7446(.A0 (n3149gat), .A1 (n614gat), .B0 (n_776), .Y (n_805));
AOI22X1 g7464(.A0 (n_1069), .A1 (n680gat), .B0 (n_1037), .B1(n1068gat), .Y (n_802));
DFFSRX1 n388gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n883gat), .Q (n388gat), .QN ());
AOI21X1 g7468(.A0 (n3149gat), .A1 (n1068gat), .B0 (n_769), .Y(n_800));
MX2X1 g7470(.A (n584gat), .B (n865gat), .S0 (n3149gat), .Y (n_798));
MX2X1 g7471(.A (n580gat), .B (n861gat), .S0 (n3149gat), .Y (n_796));
AND2X1 g7487(.A (n1829gat), .B (n1821gat), .Y (n_831));
AOI22X1 g7523(.A0 (n_1680), .A1 (n699gat), .B0 (n3149gat), .B1(n1148gat), .Y (n_795));
DFFSRX1 n2446gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_786), .Q (n2446gat), .QN ());
NOR2X1 g7290(.A (n_442), .B (n_1345), .Y (n_791));
NAND4X1 g7306(.A (n_2014), .B (n_788), .C (n_787), .D (n_597), .Y(n_789));
NAND2X1 g7335(.A (n_2021), .B (n3149gat), .Y (n_823));
AND2X1 g7343(.A (n_2024), .B (n3149gat), .Y (n_867));
MX2X1 g7389(.A (n_732), .B (n_744), .S0 (n_619), .Y (n_821));
DFFSRX1 n830gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_756), .Q (n830gat), .QN ());
DFFSRX1 n834gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_757), .Q (n834gat), .QN ());
NAND2X1 g7440(.A (n834gat), .B (n707gat), .Y (n_781));
OAI21X1 g7474(.A0 (n816gat), .A1 (n680gat), .B0 (n_755), .Y (n_778));
MX2X1 g7522(.A (n_23), .B (n271gat), .S0 (n3149gat), .Y (n_777));
DFFSRX1 n2084gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3149gat), .Q (n2084gat), .QN ());
NAND2X1 g7542(.A (n3149gat), .B (n341gat), .Y (n_776));
NAND2X1 g7543(.A (n3149gat), .B (n337gat), .Y (n_775));
OR2X1 g7287(.A (n_751), .B (n1678gat), .Y (n_774));
DFFSRX1 n1508gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_750), .Q (), .QN (n1508gat));
DFFSRX1 n820gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1812), .Q (n820gat), .QN ());
INVX1 g7431(.A (n838gat), .Y (n_782));
NAND3X1 g7444(.A (n_644), .B (n_725), .C (n_704), .Y (n_772));
INVX1 g7454(.A (n707gat), .Y (n_779));
DFFSRX1 n883gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1874), .Q (), .QN (n883gat));
DFFSRX1 n684gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_743), .Q (), .QN (n684gat));
NOR2X1 g7463(.A (n2169gat), .B (n_685), .Y (n_771));
AOI22X1 g7465(.A0 (n_1069), .A1 (n584gat), .B0 (n865gat), .B1(n_1037), .Y (n_770));
NOR2X1 g7482(.A (n3149gat), .B (n_739), .Y (n_769));
OR2X1 g7486(.A (n816gat), .B (n_739), .Y (n_767));
NAND2X1 g7488(.A (n816gat), .B (n_739), .Y (n_766));
DFFSRX1 n1829gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2029gat), .Q (), .QN (n1829gat));
DFFSRX1 n2021gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_723), .Q (n2021gat), .QN ());
NAND2X1 g7296(.A (n_763), .B (n_1382), .Y (n_764));
NAND2X1 g7315(.A (n_760), .B (n1675gat), .Y (n_761));
NAND2X1 g7318(.A (n2155gat), .B (n_141), .Y (n_2120));
NAND4X1 g7319(.A (n_736), .B (n_568), .C (n1596gat), .D (n_612), .Y(n_758));
NAND4X1 g7359(.A (n_55), .B (n2502gat), .C (n2658gat), .D (n2510gat),.Y (n_786));
DFFSRX1 n838gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_728), .Q (n838gat), .QN ());
NAND4X1 g7445(.A (n_651), .B (n_706), .C (n_687), .D (n_648), .Y(n_757));
MX2X1 g7449(.A (n3073gat), .B (n_1916), .S0 (n_2117), .Y (n_756));
DFFSRX1 n707gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_726), .Q (n707gat), .QN ());
NAND2X1 g7489(.A (n816gat), .B (n680gat), .Y (n_755));
DFFSRX1 n614gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_708), .Q (n614gat), .QN ());
AOI22X1 g7307(.A0 (n_2019), .A1 (n1462gat), .B0 (n_719), .B1(n1596gat), .Y (n_751));
INVX1 g7325(.A (n_738), .Y (n_750));
INVX1 g7329(.A (n2155gat), .Y (n_749));
NAND3X1 g7145(.A (n_2021), .B (n1336gat), .C (n_1748), .Y (n_748));
NAND3X1 g7347(.A (n_2029), .B (n2091gat), .C (n1496gat), .Y (n_788));
NAND2X1 g7349(.A (n_585), .B (n_2022), .Y (n_747));
OAI21X1 g7472(.A0 (n_730), .A1 (n_731), .B0 (n_716), .Y (n_744));
DFFSRX1 n2169gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_714), .Q (), .QN (n2169gat));
OAI21X1 g7480(.A0 (n_697), .A1 (n_1877), .B0 (n_676), .Y (n_743));
INVX1 g7503(.A (n680gat), .Y (n_739));
DFFSRX1 n2029gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_722), .Q (), .QN (n2029gat));
DFFSRX1 n1389gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_696), .Q (n1389gat), .QN ());
NOR2X1 g7320(.A (n_694), .B (n1340gat), .Y (n_763));
NAND4X1 g7326(.A (n_2024), .B (n_1198), .C (n_420), .D (n_461), .Y(n_738));
DFFSRX1 n2155gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_2019), .Q (n2155gat), .QN ());
NOR2X1 g7344(.A (n_2024), .B (n_2104), .Y (n_736));
NAND3X1 g7345(.A (n_2024), .B (n1807gat), .C (n1340gat), .Y (n_733));
NOR2X1 g7348(.A (n_671), .B (n_2024), .Y (n_760));
XOR2X1 g7429(.A (n_731), .B (n_730), .Y (n_732));
MX2X1 g7467(.A (n3066gat), .B (n_1950), .S0 (n_2117), .Y (n_728));
NAND3X1 g7494(.A (n_679), .B (n_684), .C (n_649), .Y (n_726));
AOI22X1 g7495(.A0 (n_683), .A1 (n_2056), .B0 (n_1871), .B1(n3071gat), .Y (n_725));
DFFSRX1 n816gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_703), .Q (), .QN (n816gat));
DFFSRX1 n584gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_701), .Q (), .QN (n584gat));
DFFSRX1 n680gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_700), .Q (), .QN (n680gat));
DFFSRX1 n580gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_699), .Q (), .QN (n580gat));
DFFSRX1 n2040gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_724), .Q (), .QN (n2040gat));
OR2X1 g7514(.A (n_633), .B (n_724), .Y (n_723));
INVX1 g7572(.A (n1821gat), .Y (n_722));
INVX1 g7338(.A (n_719), .Y (n_720));
NAND2X1 g7481(.A (n_730), .B (n_731), .Y (n_716));
INVX1 g7509(.A (n2176gat), .Y (n_714));
MX2X1 g7517(.A (n3068gat), .B (n_637), .S0 (n_2117), .Y (n_708));
NAND2X1 g7541(.A (n_643), .B (n_2117), .Y (n_706));
AND2X1 g7544(.A (n384gat), .B (n_2101), .Y (n_705));
NAND2X1 g7546(.A (n_613), .B (n_1878), .Y (n_704));
NAND4X1 g7556(.A (n_519), .B (n_527), .C (n_1550), .D (n_575), .Y(n_724));
OAI21X1 g7558(.A0 (n_1875), .A1 (n_36), .B0 (n_645), .Y (n_703));
OAI21X1 g7560(.A0 (n_1875), .A1 (n_38), .B0 (n_634), .Y (n_701));
OAI21X1 g7561(.A0 (n_1875), .A1 (n_46), .B0 (n_646), .Y (n_700));
OAI21X1 g7563(.A0 (n_1875), .A1 (n_44), .B0 (n_623), .Y (n_699));
DFFSRX1 n2091gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1748), .Q (), .QN (n2091gat));
XOR2X1 g7565(.A (n327gat), .B (n_611), .Y (n_697));
NOR2X1 g7301(.A (n_630), .B (n_523), .Y (n_696));
AND2X1 g7339(.A (n_2021), .B (n_2103), .Y (n_719));
AND2X1 g7342(.A (n_627), .B (n_2024), .Y (n_1531));
OAI21X1 g7350(.A0 (n_1748), .A1 (n_2104), .B0 (n_2019), .Y (n_694));
DFFSRX1 n2510gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_691), .Q (n2510gat), .QN ());
DFFSRX1 n1821gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_639), .Q (n1821gat), .QN ());
XOR2X1 g7473(.A (n_689), .B (n_1924), .Y (n_690));
NAND4X1 g7485(.A (n_2117), .B (n148gat), .C (n_1947), .D (n_1949), .Y(n_687));
DFFSRX1 n2176gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_685), .Q (n2176gat), .QN ());
NAND2X1 g7539(.A (n_616), .B (n3067gat), .Y (n_684));
NOR2X1 g7545(.A (n331gat), .B (n_1734), .Y (n_683));
NAND2X1 g7548(.A (n_1924), .B (n_689), .Y (n_681));
NAND3X1 g7549(.A (n_1685), .B (n_578), .C (n_856), .Y (n_680));
NAND2X1 g7550(.A (n_614), .B (n_2117), .Y (n_679));
AOI22X1 g7562(.A0 (n_1871), .A1 (n3070gat), .B0 (n3079gat), .B1(n_1872), .Y (n_676));
DFFSRX1 n2506gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_593), .Q (n2506gat), .QN ());
DFFSRX1 n1880gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_604), .Q (n1880gat), .QN ());
DFFSRX1 n1496gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n1394gat), .Q (), .QN (n1496gat));
NAND2X1 g7592(.A (n_1748), .B (n1394gat), .Y (n_671));
OR2X1 g7511(.A (n_617), .B (n_667), .Y (n3104gat));
DFFSRX1 n1767gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_595), .Q (), .QN (n1767gat));
DFFSRX1 n2658gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_620), .Q (n2658gat), .QN ());
AND2X1 g7185(.A (n_610), .B (n_390), .Y (n3138gat));
AOI21X1 g7518(.A0 (n_566), .A1 (n673gat), .B0 (n_591), .Y (n_730));
NAND2X1 g7529(.A (n_659), .B (n3068gat), .Y (n_661));
NAND2X1 g7530(.A (n_659), .B (n3065gat), .Y (n_660));
NAND2X1 g7531(.A (n_659), .B (n3069gat), .Y (n_658));
NAND2X1 g7532(.A (n_659), .B (n3066gat), .Y (n_657));
NAND2X1 g7533(.A (n_659), .B (n3067gat), .Y (n_656));
NAND2X1 g7534(.A (n_659), .B (n3070gat), .Y (n_655));
NAND2X1 g7535(.A (n_659), .B (n3073gat), .Y (n_654));
NAND2X1 g7536(.A (n_659), .B (n3072gat), .Y (n_653));
NAND2X1 g7537(.A (n_659), .B (n3071gat), .Y (n_652));
NAND2X1 g7538(.A (n_616), .B (n3065gat), .Y (n_651));
NAND3X1 g7551(.A (n_2117), .B (n_0), .C (n156gat), .Y (n_649));
NAND3X1 g7552(.A (n_2118), .B (n_198), .C (n256gat), .Y (n_648));
DFFSRX1 n2182gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_579), .Q (n2182gat), .QN ());
NAND2X1 g7585(.A (n3074gat), .B (n_1872), .Y (n_646));
NAND2X1 g7586(.A (n_1872), .B (n3076gat), .Y (n_645));
NAND2X1 g7587(.A (n3080gat), .B (n_1872), .Y (n_644));
NOR2X1 g7589(.A (n148gat), .B (n_1949), .Y (n_643));
AOI21X1 g7590(.A0 (n271gat), .A1 (n_1037), .B0 (n_573), .Y (n_642));
NOR2X1 g7602(.A (n_581), .B (n_1120), .Y (n_1140));
NOR2X1 g7625(.A (n2319gat), .B (n3099gat), .Y (n_639));
NOR2X1 g7629(.A (n_567), .B (n_1754), .Y (n_638));
OAI21X1 g7639(.A0 (n156gat), .A1 (n_549), .B0 (n_1917), .Y (n_637));
NAND2X1 g7540(.A (n_584), .B (n_489), .Y (n3105gat));
NAND2X1 g7581(.A (n3077gat), .B (n_1872), .Y (n_634));
NAND2X1 g7679(.A (n_632), .B (n_631), .Y (n_633));
INVX1 g7323(.A (n_1702), .Y (n_630));
NAND2X1 g7580(.A (n3075gat), .B (n_1872), .Y (n_623));
NAND2X1 g7420(.A (n_432), .B (n_563), .Y (n_622));
MX2X1 g7451(.A (n_499), .B (n_537), .S0 (n_167), .Y (n_691));
INVX1 g7566(.A (n_620), .Y (n_621));
AOI21X1 g7519(.A0 (n_522), .A1 (n861gat), .B0 (n_590), .Y (n_731));
AOI21X1 g7520(.A0 (n_536), .A1 (n1148gat), .B0 (n_586), .Y (n_619));
INVX1 g7524(.A (n2095gat), .Y (n_685));
OAI22X1 g7557(.A0 (n_588), .A1 (n_421), .B0 (n_587), .B1 (n_320), .Y(n_617));
INVX1 g7582(.A (n_2118), .Y (n_616));
NOR2X1 g7600(.A (n1462gat), .B (n1394gat), .Y (n_615));
OAI21X1 g7601(.A0 (n_580), .A1 (n_196), .B0 (n_329), .Y (n_1125));
OAI21X1 g7604(.A0 (n_410), .A1 (n_202), .B0 (n_561), .Y (n_659));
MX2X1 g7607(.A (n_1396), .B (n_1951), .S0 (n152gat), .Y (n_614));
MX2X1 g7610(.A (n388gat), .B (n_1497), .S0 (n331gat), .Y (n_613));
DFFSRX1 n2179gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1216), .Q (), .QN (n2179gat));
INVX1 g7620(.A (n_1721), .Y (n_611));
AND2X1 g7626(.A (n_1486), .B (n_1216), .Y (n_610));
NOR2X1 g7579(.A (n_558), .B (n_603), .Y (n_604));
AOI22X1 g7656(.A0 (n_569), .A1 (n673gat), .B0 (n_600), .B1 (n_1071),.Y (n_602));
OR2X1 g7312(.A (n_2033), .B (n_597), .Y (n_598));
INVX1 g7742(.A (n_632), .Y (n_595));
INVX1 g7164(.A (n_592), .Y (n_593));
XOR2X1 g7567(.A (n_424), .B (n_533), .Y (n_620));
DFFSRX1 n2095gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_562), .Q (n2095gat), .QN ());
AOI21X1 g7553(.A0 (n_481), .A1 (n_475), .B0 (n673gat), .Y (n_591));
AOI21X1 g7554(.A0 (n_479), .A1 (n_476), .B0 (n861gat), .Y (n_590));
NAND3X1 g7588(.A (n_588), .B (n_587), .C (n_303), .Y (n3151gat));
NOR2X1 g7591(.A (n_521), .B (n1148gat), .Y (n_586));
NOR2X1 g7599(.A (n1588gat), .B (n1596gat), .Y (n_585));
AOI22X1 g7603(.A0 (n_560), .A1 (n_466), .B0 (n_409), .B1 (n_220), .Y(n_584));
INVX1 g7613(.A (n1394gat), .Y (n_612));
DFFSRX1 n1340gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_524), .Q (n1340gat), .QN ());
NOR2X1 g7624(.A (n_580), .B (n_195), .Y (n_581));
OR2X1 g7627(.A (n_2074), .B (n_2104), .Y (n_579));
OR2X1 g7632(.A (n_518), .B (n_2103), .Y (n_578));
NOR2X1 g7637(.A (n_574), .B (n_1216), .Y (n_575));
OAI22X1 g7640(.A0 (n_493), .A1 (n834gat), .B0 (n_981), .B1(n1035gat), .Y (n_573));
AOI22X1 g7648(.A0 (n_396), .A1 (n_402), .B0 (n_569), .B1 (n_506), .Y(n_570));
INVX1 g7660(.A (n1678gat), .Y (n_568));
INVX1 g7662(.A (n1834gat), .Y (n_567));
DFFSRX1 n2319gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2472gat), .Q (), .QN (n2319gat));
OAI21X1 g7708(.A0 (n_860), .A1 (n1241gat), .B0 (n_511), .Y (n_566));
NAND2X1 g7743(.A (n_505), .B (n_458), .Y (n_632));
AOI21X1 g7802(.A0 (n_389), .A1 (n341gat), .B0 (n_501), .Y (n_565));
AOI21X1 g7165(.A0 (n_503), .A1 (n_502), .B0 (n_504), .Y (n_592));
AOI21X1 g7448(.A0 (n614gat), .A1 (n_1898), .B0 (n_431), .Y (n_563));
DFFSRX1 n1740gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n1332gat), .Q (n1740gat), .QN ());
OAI21X1 g7605(.A0 (n_1595), .A1 (n_463), .B0 (n_411), .Y (n_562));
DFFSRX1 n1394gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_496), .Q (), .QN (n1394gat));
NAND2X1 g7631(.A (n_462), .B (n_560), .Y (n_561));
NAND2X1 g7641(.A (n2117gat), .B (n2125gat), .Y (n_558));
AOI21X1 g7650(.A0 (n842gat), .A1 (n_1037), .B0 (n_495), .Y (n_557));
AOI21X1 g7651(.A0 (n1241gat), .A1 (n_1037), .B0 (n_491), .Y (n_556));
AOI22X1 g7652(.A0 (n_448), .A1 (n_1037), .B0 (n_554), .B1 (n_1071),.Y (n_555));
AOI22X1 g7653(.A0 (n_447), .A1 (n_1037), .B0 (n_2035), .B1 (n_1071),.Y (n_553));
DFFSRX1 n1678gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_483), .Q (n1678gat), .QN ());
DFFSRX1 n1834gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_484), .Q (n1834gat), .QN ());
NAND2X1 g7687(.A (n_2055), .B (n388gat), .Y (n_1571));
NAND3X1 g7695(.A (n_2050), .B (n327gat), .C (n_1498), .Y (n_547));
NAND2X1 g7333(.A (n_2015), .B (n_2), .Y (n_787));
NAND2X1 g7340(.A (n_2015), .B (n1740gat), .Y (n_597));
XOR2X1 g7493(.A (n_498), .B (n_468), .Y (n_537));
XOR2X1 g7608(.A (n865gat), .B (n1080gat), .Y (n_536));
XOR2X1 g7609(.A (n2644gat), .B (n_423), .Y (n_535));
DFFSRX1 n1596gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_464), .Q (), .QN (n1596gat));
NAND3X1 g7645(.A (n_418), .B (n_419), .C (n_374), .Y (n_588));
AOI21X1 g7649(.A0 (n_336), .A1 (n_145), .B0 (n_455), .Y (n_533));
AOI22X1 g7654(.A0 (n1080gat), .A1 (n_1037), .B0 (n_531), .B1(n_1071), .Y (n_532));
AOI22X1 g7655(.A0 (n861gat), .A1 (n_1037), .B0 (n337gat), .B1(n_1071), .Y (n_530));
XOR2X1 g7657(.A (n1975gat), .B (n_415), .Y (n_529));
OR2X1 g7670(.A (n_1069), .B (n_1037), .Y (n_998));
NOR2X1 g7697(.A (n_523), .B (n_482), .Y (n_524));
OAI21X1 g7704(.A0 (n_311), .A1 (n_226), .B0 (n_451), .Y (n_580));
XOR2X1 g7709(.A (n957gat), .B (n1068gat), .Y (n_522));
XOR2X1 g7710(.A (n865gat), .B (n1080gat), .Y (n_521));
DFFSRX1 n2472gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_437), .Q (), .QN (n2472gat));
INVX1 g7734(.A (n_518), .Y (n_519));
NOR2X1 g7740(.A (n_1698), .B (n_1697), .Y (n_515));
NAND2X1 g7787(.A (n_860), .B (n1241gat), .Y (n_511));
DFFSRX1 n1336gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_435), .Q (n1336gat), .QN ());
NOR2X1 g7871(.A (n_600), .B (n_500), .Y (n_505));
NOR2X1 g7175(.A (n_503), .B (n_502), .Y (n_504));
NOR2X1 g7881(.A (n_500), .B (n341gat), .Y (n_501));
XOR2X1 g7568(.A (n_498), .B (n_467), .Y (n_499));
NAND2X1 g7623(.A (n_381), .B (n1035gat), .Y (n3108gat));
DFFSRX1 n1462gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_427), .Q (n1462gat), .QN ());
DFFSRX1 n1332gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_405), .Q (), .QN (n1332gat));
DFFSRX1 n2117gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2121gat), .Q (n2117gat), .QN ());
DFFSRX1 n1588gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_404), .Q (n1588gat), .QN ());
AND2X1 g7675(.A (n_413), .B (n_310), .Y (n_496));
NOR2X1 g7676(.A (n_493), .B (n830gat), .Y (n_495));
NOR2X1 g7690(.A (n_493), .B (n699gat), .Y (n_494));
NOR2X1 g7696(.A (n_493), .B (n820gat), .Y (n_491));
INVX1 g7698(.A (n_489), .Y (n_490));
NOR2X1 g7702(.A (n_418), .B (n_1600), .Y (n_560));
DFFSRX1 n1525gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_397), .Q (), .QN (n1525gat));
INVX1 g7732(.A (n_1396), .Y (n_549));
INVX1 g7736(.A (n_1834), .Y (n_518));
INVX1 g7749(.A (n_487), .Y (n_574));
INVX1 g7756(.A (n_981), .Y (n_1075));
INVX1 g7763(.A (n_631), .Y (n_484));
INVX1 g7770(.A (n_482), .Y (n_483));
NAND2X1 g7775(.A (n1294gat), .B (n1241gat), .Y (n_481));
NAND2X1 g7778(.A (n957gat), .B (n1068gat), .Y (n_479));
OR2X1 g7788(.A (n957gat), .B (n1068gat), .Y (n_476));
OR2X1 g7789(.A (n1294gat), .B (n1241gat), .Y (n_475));
INVX1 g7807(.A (n673gat), .Y (n_506));
MX2X1 g7606(.A (n_326), .B (n_259), .S0 (n337gat), .Y (n_689));
INVX1 g7646(.A (n_467), .Y (n_468));
DFFSRX1 n1807gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_2031), .Q (), .QN (n1807gat));
INVX1 g7685(.A (n_1596), .Y (n_466));
NOR2X1 g7689(.A (n_426), .B (n_1373), .Y (n_464));
INVX1 g7691(.A (n_462), .Y (n_463));
NOR2X1 g7699(.A (n_369), .B (n_461), .Y (n_489));
NAND2X1 g7750(.A (n_1551), .B (n_458), .Y (n_487));
NAND2X1 g7758(.A (n_454), .B (n_406), .Y (n_981));
NAND2X1 g7764(.A (n_458), .B (n_1552), .Y (n_631));
NOR2X1 g7765(.A (n_339), .B (n_145), .Y (n_455));
AND2X1 g7767(.A (n_454), .B (n_249), .Y (n_569));
NAND2X1 g7768(.A (n_357), .B (n_458), .Y (n_527));
NAND3X1 g7771(.A (n_111), .B (n_303), .C (n_1559), .Y (n_482));
INVX1 g7781(.A (n_493), .Y (n_1069));
AOI21X1 g7803(.A0 (n_1211), .A1 (n_350), .B0 (n_351), .Y (n_452));
AOI22X1 g7791(.A0 (n_312), .A1 (n_221), .B0 (n_1670), .B1 (n_277), .Y(n_451));
INVX1 g7812(.A (n1294gat), .Y (n_860));
INVX1 g7816(.A (n957gat), .Y (n_448));
INVX1 g7819(.A (n1148gat), .Y (n_447));
NOR2X1 g7847(.A (n830gat), .B (n_384), .Y (n_444));
INVX1 g7859(.A (n_1453), .Y (n_442));
OR2X1 g7868(.A (n_1514), .B (n_342), .Y (n_1697));
NOR2X1 g7873(.A (n_344), .B (n_355), .Y (n_437));
NOR2X1 g7879(.A (n_386), .B (n842gat), .Y (n_436));
INVX1 g7181(.A (n_391), .Y (n_435));
AOI21X1 g7183(.A0 (n_237), .A1 (n_157), .B0 (n_347), .Y (n_503));
AOI21X1 g7447(.A0 (n614gat), .A1 (n_1211), .B0 (n_338), .Y (n_432));
NOR2X1 g7462(.A (n614gat), .B (n_388), .Y (n_431));
INVX1 g7967(.A (n_1898), .Y (n_500));
OR2X1 g7703(.A (n_210), .B (n_428), .Y (n3150gat));
AOI21X1 g7647(.A0 (n_164), .A1 (n3084gat), .B0 (n_328), .Y (n_467));
NOR2X1 g7671(.A (n_426), .B (n_2032), .Y (n_427));
AOI22X1 g7658(.A0 (n_235), .A1 (n_100), .B0 (n_274), .B1 (n_85), .Y(n_424));
NOR2X1 g7681(.A (n_325), .B (n_143), .Y (n_423));
NOR2X1 g7692(.A (n_422), .B (n_421), .Y (n_462));
XOR2X1 g7711(.A (n_420), .B (n_414), .Y (n_667));
DFFSRX1 n1675gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_315), .Q (), .QN (n1675gat));
DFFSRX1 n2121gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2125gat), .Q (), .QN (n2121gat));
INVX1 g7720(.A (n_1600), .Y (n_419));
INVX1 g7722(.A (n_1598), .Y (n_418));
AND2X1 g7728(.A (n_316), .B (n_414), .Y (n_415));
NOR2X1 g7729(.A (n_403), .B (n_412), .Y (n_413));
AND2X1 g7741(.A (n_407), .B (n_249), .Y (n_1037));
NAND2X1 g7744(.A (n_203), .B (n_2098), .Y (n_411));
NAND2X1 g7751(.A (n_409), .B (n_83), .Y (n_410));
AND2X1 g7766(.A (n_407), .B (n_406), .Y (n_1071));
NOR2X1 g7769(.A (n_319), .B (n_523), .Y (n_405));
NOR2X1 g7779(.A (n_403), .B (n_1), .Y (n_404));
NAND3X1 g7786(.A (n_402), .B (n_395), .C (n_406), .Y (n_493));
INVX1 g7795(.A (n_400), .Y (n_401));
DFFSRX1 n673gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_289), .Q (), .QN (n673gat));
DFFSRX1 n1068gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_330), .Q (), .QN (n1068gat));
DFFSRX1 n1294gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_294), .Q (n1294gat), .QN ());
DFFSRX1 n1080gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_295), .Q (), .QN (n1080gat));
DFFSRX1 n957gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_292), .Q (n957gat), .QN ());
DFFSRX1 n1148gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_313), .Q (n1148gat), .QN ());
DFFSRX1 n865gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_293), .Q (), .QN (n865gat));
AND2X1 g7852(.A (n_306), .B (n_256), .Y (n_397));
NOR2X1 g7855(.A (n_395), .B (n_249), .Y (n_396));
NAND4X1 g7182(.A (n_390), .B (n_271), .C (n_145), .D (n_174), .Y(n_391));
INVX1 g7958(.A (n_388), .Y (n_389));
INVX1 g7960(.A (n_386), .Y (n_387));
INVX1 g7976(.A (n_384), .Y (n_385));
INVX1 g7979(.A (n_1902), .Y (n_382));
INVX1 g7712(.A (n_380), .Y (n_381));
DFFSRX1 n1241gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_291), .Q (), .QN (n1241gat));
DFFSRX1 n861gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_296), .Q (), .QN (n861gat));
AND2X1 g7846(.A (n_377), .B (n_376), .Y (n_378));
AND2X1 g7843(.A (n_376), .B (n_835), .Y (n_375));
DFFSRX1 n2347gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_95), .Q (n2347gat), .QN ());
NAND2X1 g7961(.A (n_356), .B (n_2003), .Y (n_386));
XOR2X1 g7713(.A (n2407gat), .B (n_324), .Y (n_380));
INVX1 g7718(.A (n_422), .Y (n_374));
NAND3X1 g7725(.A (n_262), .B (n_207), .C (n_172), .Y (n_502));
OR4X1 g7738(.A (n_1669), .B (n_1505), .C (n_333), .D (n3085gat), .Y(n_587));
OAI21X1 g7792(.A0 (n_1984), .A1 (n_1547), .B0 (n_273), .Y (n_369));
INVX1 g7796(.A (n_1888), .Y (n_400));
NOR2X1 g7836(.A (n_402), .B (n_395), .Y (n_454));
INVX1 g8058(.A (n_367), .Y (n_600));
NAND2X1 g7842(.A (n_377), .B (n_1685), .Y (n_366));
AND2X1 g7845(.A (n_833), .B (n_376), .Y (n_365));
AND2X1 g7854(.A (n_1686), .B (n_376), .Y (n_364));
NOR2X1 g7872(.A (n_356), .B (n_355), .Y (n_357));
NOR2X1 g7880(.A (n_355), .B (n_350), .Y (n_351));
OAI21X1 g7188(.A0 (n2634gat), .A1 (n_290), .B0 (n_244), .Y (n_347));
NAND2X1 g7959(.A (n_531), .B (n_2035), .Y (n_388));
INVX1 g7963(.A (n_1922), .Y (n_344));
INVX1 g7970(.A (n_1892), .Y (n_343));
INVX1 g7971(.A (n_1892), .Y (n_342));
NAND2X1 g7977(.A (n_356), .B (n_2007), .Y (n_384));
AOI21X1 g7989(.A0 (n_1494), .A1 (n_335), .B0 (n_269), .Y (n_339));
NOR2X1 g7461(.A (n614gat), .B (n_355), .Y (n_338));
DFFSRX1 n2102gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_258), .Q (n2102gat), .QN ());
XOR2X1 g7805(.A (n_335), .B (n_1494), .Y (n_336));
NOR2X1 g7844(.A (n_1669), .B (n_333), .Y (n_409));
XOR2X1 g7804(.A (n_1559), .B (n_1984), .Y (n_428));
OR2X1 g7638(.A (n_229), .B (n_1354), .Y (n_914));
OR2X1 g7727(.A (n_75), .B (n_1708), .Y (n_2033));
INVX1 g8005(.A (n_239), .Y (n_330));
NAND4X1 g7705(.A (n_322), .B (n_218), .C (n_227), .D (n_209), .Y(n_329));
OAI21X1 g7706(.A0 (n_136), .A1 (n3084gat), .B0 (n_205), .Y (n_328));
XOR2X1 g7707(.A (n_554), .B (n271gat), .Y (n_326));
INVX1 g8059(.A (n_356), .Y (n_367));
NAND3X1 g7719(.A (n3087gat), .B (n_1506), .C (n_1528), .Y (n_422));
NAND2X1 g7753(.A (n_74), .B (n_324), .Y (n_325));
AND2X1 g7793(.A (n_213), .B (n_322), .Y (n_1120));
NAND2X1 g7826(.A (n_318), .B (n_1198), .Y (n_403));
AND2X1 g7830(.A (n_252), .B (n_395), .Y (n_407));
NAND4X1 g7850(.A (n_268), .B (n_63), .C (n_266), .D (n_26), .Y(n_426));
NAND2X1 g7856(.A (n_318), .B (n_1984), .Y (n_319));
NAND2X1 g7882(.A (n_231), .B (n_1201), .Y (n_316));
INVX1 g7883(.A (n_314), .Y (n_315));
INVX1 g8001(.A (n_240), .Y (n_313));
AND2X1 g7896(.A (n_196), .B (n_311), .Y (n_312));
NOR2X1 g7898(.A (n_194), .B (n2407gat), .Y (n_310));
DFFSRX1 n2407gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_1493), .Q (n2407gat), .QN ());
NOR2X1 g7937(.A (n_217), .B (n_1241), .Y (n_306));
INVX1 g7947(.A (n_302), .Y (n_303));
INVX1 g7991(.A (n_279), .Y (n_296));
INVX1 g7993(.A (n_243), .Y (n_295));
INVX1 g7995(.A (n_242), .Y (n_294));
INVX1 g7997(.A (n_241), .Y (n_293));
INVX1 g7999(.A (n_260), .Y (n_292));
INVX1 g8003(.A (n_282), .Y (n_291));
NOR2X1 g7196(.A (n_215), .B (n_290), .Y (n_390));
INVX1 g8007(.A (n_238), .Y (n_289));
NOR2X1 g8138(.A (n_1494), .B (n_145), .Y (n_2115));
DFFSRX1 n2125gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_211), .Q (), .QN (n2125gat));
AOI22X1 g8004(.A0 (n3082gat), .A1 (n_278), .B0 (n3073gat), .B1(n_277), .Y (n_282));
DFFSRX1 n2139gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_129), .Q (n_1581), .QN ());
AND2X1 g7862(.A (n_281), .B (n3147gat), .Y (n_603));
DFFSRX1 n2403gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_156), .Q (), .QN (n2403gat));
AOI22X1 g7992(.A0 (n3075gat), .A1 (n_278), .B0 (n3066gat), .B1(n_277), .Y (n_279));
OAI21X1 g7794(.A0 (n2640gat), .A1 (n2562gat), .B0 (n_185), .Y(n_274));
NAND3X1 g7831(.A (n_1984), .B (n_1559), .C (n_1547), .Y (n_273));
DFFSRX1 n2440gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_177), .Q (n2440gat), .QN ());
NAND2X1 g7832(.A (n_169), .B (n_1984), .Y (n_414));
AND2X1 g7839(.A (n_1080), .B (n_376), .Y (n_270));
NOR2X1 g8110(.A (n_1494), .B (n_335), .Y (n_269));
NAND4X1 g7857(.A (n_268), .B (n_143), .C (n_266), .D (n_142), .Y(n_523));
DFFSRX1 n2394gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_100), .Q (n2394gat), .QN ());
NAND4X1 g7884(.A (n_111), .B (n_1241), .C (n_1559), .D (n_1580), .Y(n_314));
AOI22X1 g7886(.A0 (n_141), .A1 (n_170), .B0 (n_261), .B1 (n_171), .Y(n_262));
XOR2X1 g7887(.A (n_266), .B (n_130), .Y (n_929));
AOI22X1 g8000(.A0 (n3076gat), .A1 (n_278), .B0 (n3067gat), .B1(n_277), .Y (n_260));
XOR2X1 g7888(.A (n160gat), .B (n271gat), .Y (n_259));
NOR2X1 g7895(.A (n_248), .B (n_174), .Y (n_854));
XOR2X1 g8011(.A (n3089gat), .B (n3088gat), .Y (n_498));
INVX1 g7901(.A (n_257), .Y (n_258));
NOR2X1 g7905(.A (n_254), .B (n_174), .Y (n_835));
NOR2X1 g7906(.A (n_1566), .B (n_174), .Y (n_833));
NOR2X1 g7907(.A (n_1577), .B (n_1559), .Y (n_256));
NOR2X1 g7912(.A (n_1566), .B (n_253), .Y (n_377));
INVX1 g7914(.A (n_252), .Y (n_402));
AND2X1 g7929(.A (n_1852), .B (n_2008), .Y (n_458));
INVX1 g7932(.A (n_249), .Y (n_406));
NOR2X1 g7938(.A (n_248), .B (n_177), .Y (n_829));
INVX1 g7984(.A (n_1882), .Y (n_355));
NAND2X1 g7192(.A (n_158), .B (n2634gat), .Y (n_244));
AOI22X1 g7994(.A0 (n3079gat), .A1 (n_278), .B0 (n3070gat), .B1(n_277), .Y (n_243));
AOI22X1 g7996(.A0 (n3080gat), .A1 (n_278), .B0 (n3071gat), .B1(n_277), .Y (n_242));
AOI22X1 g7998(.A0 (n3077gat), .A1 (n_278), .B0 (n3068gat), .B1(n_277), .Y (n_241));
NAND2X1 g7949(.A (n_1759), .B (n_1580), .Y (n_302));
AOI22X1 g8002(.A0 (n3078gat), .A1 (n_278), .B0 (n3069gat), .B1(n_277), .Y (n_240));
AOI22X1 g8006(.A0 (n3074gat), .A1 (n_278), .B0 (n3065gat), .B1(n_277), .Y (n_239));
AOI22X1 g8008(.A0 (n3081gat), .A1 (n_278), .B0 (n3072gat), .B1(n_277), .Y (n_238));
XOR2X1 g7199(.A (n2634gat), .B (n_2063), .Y (n_237));
INVX1 g8093(.A (n_1088), .Y (n_287));
XOR2X1 g8009(.A (n2640gat), .B (n_174), .Y (n_235));
INVX1 g8060(.A (n919gat), .Y (n_356));
NAND2X1 g7957(.A (n_1241), .B (n_1559), .Y (n_231));
INVX1 g7197(.A (n_154), .Y (n_2121));
DFFSRX1 n1850gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_2063), .Q (n1850gat), .QN ());
AOI21X1 g7701(.A0 (n_228), .A1 (n_266), .B0 (n2347gat), .Y (n_229));
NOR2X1 g7933(.A (n_227), .B (n_226), .Y (n_249));
OAI21X1 g7824(.A0 (n_1670), .A1 (n3085gat), .B0 (n3095gat), .Y(n_322));
NAND2X1 g7835(.A (n_121), .B (n_228), .Y (n_324));
NAND2X1 g8094(.A (n_1493), .B (n_145), .Y (n_1088));
AND2X1 g7897(.A (n_208), .B (n_226), .Y (n_221));
NAND2X1 g7902(.A (n_1852), .B (n271gat), .Y (n_257));
INVX1 g7903(.A (n_219), .Y (n_220));
OR2X1 g7915(.A (n_218), .B (n_311), .Y (n_252));
NOR2X1 g7916(.A (n_217), .B (n_1559), .Y (n_318));
NAND2X1 g7918(.A (n_206), .B (n_170), .Y (n_215));
NOR2X1 g7919(.A (n2454gat), .B (n_2004), .Y (n_457));
OR2X1 g7921(.A (n_218), .B (n_227), .Y (n_213));
INVX1 g7889(.A (n2110gat), .Y (n_211));
AND2X1 g7925(.A (n_1852), .B (n337gat), .Y (n_210));
OR2X1 g7934(.A (n_209), .B (n_208), .Y (n_395));
NAND2X1 g7943(.A (n_206), .B (n_129), .Y (n_207));
NAND2X1 g7944(.A (n_1668), .B (n3085gat), .Y (n_205));
NOR2X1 g7946(.A (n_1559), .B (n_1547), .Y (n_461));
NOR2X1 g7952(.A (n_117), .B (n_202), .Y (n_203));
NAND2X1 g7926(.A (n2099gat), .B (n_106), .Y (n_199));
INVX1 g8026(.A (n148gat), .Y (n_198));
INVX1 g8075(.A (n_197), .Y (n_531));
INVX1 g8141(.A (n_195), .Y (n_196));
NAND2X1 g8144(.A (n_143), .B (n2347gat), .Y (n_194));
AND2X1 g7917(.A (n_1483), .B (n_2067), .Y (n_271));
DFFSRX1 n1899gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_90), .Q (n1899gat), .QN ());
NAND2X1 g8139(.A (n2640gat), .B (n2562gat), .Y (n_185));
NAND2X1 g8090(.A (n_85), .B (n_156), .Y (n_254));
DFFSRX1 n2061gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_2048), .Q (n_1562), .QN ());
DFFSRX1 n2110gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n2033gat), .Q (n2110gat), .QN ());
DFFSRX1 n148gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_23), .Q (n148gat), .QN ());
NAND3X1 g7840(.A (n_73), .B (n_175), .C (n_143), .Y (n_627));
AND2X1 g7927(.A (n_2066), .B (n_177), .Y (n_856));
NOR2X1 g7945(.A (n_1759), .B (n_1577), .Y (n_1984));
AND2X1 g7894(.A (n_2066), .B (n_174), .Y (n_1080));
NAND2X1 g7904(.A (n_173), .B (n_83), .Y (n_219));
NAND3X1 g7922(.A (n_171), .B (n_2046), .C (n_170), .Y (n_172));
AND2X1 g7928(.A (n_1559), .B (n_1544), .Y (n_169));
XOR2X1 g8012(.A (n3087gat), .B (n3086gat), .Y (n_167));
XOR2X1 g7990(.A (n_135), .B (n3085gat), .Y (n_164));
DFFSRX1 n384gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_21), .Q (), .QN (n384gat));
INVX1 g8044(.A (n2135gat), .Y (n_162));
INVX1 g8056(.A (n341gat), .Y (n_350));
INVX1 g8072(.A (n160gat), .Y (n_554));
INVX1 g8076(.A (n_1881), .Y (n_197));
OR2X1 g8084(.A (n3087gat), .B (n_1267), .Y (n_333));
NAND2X1 g8098(.A (n_63), .B (n2394gat), .Y (n_159));
NOR2X1 g7208(.A (n_157), .B (n_2059), .Y (n_158));
NAND2X1 g8104(.A (n_100), .B (n_156), .Y (n_248));
NOR2X1 g7198(.A (n_66), .B (n_153), .Y (n_154));
DFFSRX1 n1312gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n1363gat), .Q (n1312gat), .QN ());
NAND2X1 g8143(.A (n_277), .B (n3088gat), .Y (n_195));
NAND2X1 g7920(.A (n2446gat), .B (n2450gat), .Y (n3147gat));
DFFSRX1 n919gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3072gat), .Q (n919gat), .QN ());
INVX1 g8122(.A (n_132), .Y (n_141));
DFFSRX1 n337gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3066gat), .Q (), .QN (n337gat));
XOR2X1 g8010(.A (n_31), .B (n_54), .Y (n_140));
DFFSRX1 n2143gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_157), .Q (n_1548), .QN ());
OR2X1 g8101(.A (n_135), .B (n3085gat), .Y (n_136));
NOR2X1 g8091(.A (n_1647), .B (n2347gat), .Y (n_268));
AND2X1 g7953(.A (n_175), .B (n_50), .Y (n_131));
INVX2 g8119(.A (n_228), .Y (n_130));
INVX1 g8153(.A (n_156), .Y (n_335));
NOR2X1 g8099(.A (n_1493), .B (n_145), .Y (n_376));
NAND2X1 g7853(.A (n_398), .B (n_1647), .Y (n_1698));
NOR2X1 g7205(.A (n_2064), .B (n_90), .Y (n_122));
AND2X1 g7941(.A (n_266), .B (n_72), .Y (n_121));
AND2X1 g8097(.A (n_1525), .B (n_80), .Y (n_165));
DFFSRX1 n2190gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3127gat), .Q (n2190gat), .QN ());
INVX1 g8051(.A (n2450gat), .Y (n3148gat));
DFFSRX1 n2135gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3126gat), .Q (n2135gat), .QN ());
INVX1 g8088(.A (n_116), .Y (n_117));
OR2X1 g7207(.A (n_157), .B (n_2063), .Y (n_290));
NOR2X1 g8100(.A (n_171), .B (n_2048), .Y (n_206));
AND2X1 g8105(.A (n3093gat), .B (n3087gat), .Y (n_208));
INVX1 g8113(.A (n_111), .Y (n_217));
AND2X1 g8117(.A (n3093gat), .B (n3085gat), .Y (n_226));
INVX1 g8133(.A (n_1259), .Y (n_106));
DFFSRX1 n160gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3067gat), .Q (n160gat), .QN ());
NAND2X1 g8111(.A (n3086gat), .B (n3085gat), .Y (n_202));
AND2X1 g8116(.A (n3093gat), .B (n3086gat), .Y (n_311));
DFFSRX1 n271gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3065gat), .Q (), .QN (n271gat));
AND2X1 g8106(.A (n3095gat), .B (n3086gat), .Y (n_227));
DFFSRX1 n341gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3068gat), .Q (), .QN (n341gat));
DFFSRX1 n463gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_10), .Q (n463gat), .QN ());
BUFX3 g8279(.A (n3093gat), .Y (n_277));
AND2X1 g8120(.A (n_63), .B (n_4), .Y (n_228));
AND2X1 g8125(.A (n_5), .B (n_95), .Y (n_96));
DFFSRX1 n2450gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(1'b0), .Q (n2450gat), .QN ());
DFFSRX1 n156gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_42), .Q (n156gat), .QN ());
NAND2X1 g8124(.A (n_90), .B (n_2049), .Y (n_132));
INVX1 g8244(.A (n_85), .Y (n_100));
NOR2X1 g8114(.A (n_1544), .B (n_1504), .Y (n_111));
OR2X1 g7913(.A (n_142), .B (n2403gat), .Y (n_412));
INVX1 g8128(.A (n_320), .Y (n_83));
DFFSRX1 n398gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3069gat), .Q (n398gat), .QN ());
AND2X1 g8089(.A (n3087gat), .B (n_1267), .Y (n_116));
DFFSRX1 n1975gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_3), .Q (), .QN (n1975gat));
INVX1 g8154(.A (n_80), .Y (n_156));
AND2X1 g8130(.A (n_2049), .B (n_65), .Y (n_261));
AND2X1 g8118(.A (n3095gat), .B (n3088gat), .Y (n_209));
DFFSRX1 n402gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3070gat), .Q (n402gat), .QN ());
NAND2X1 g8115(.A (n_1573), .B (n_1546), .Y (n_75));
INVX1 g7899(.A (n_73), .Y (n_74));
AND2X1 g8102(.A (n_1505), .B (n3085gat), .Y (n_173));
DFFSRX1 n2644gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_18), .Q (), .QN (n2644gat));
DFFSRX1 n1363gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_12), .Q (), .QN (n1363gat));
DFFSRX1 n470gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_9), .Q (), .QN (n470gat));
DFFSRX1 n2033gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_8), .Q (), .QN (n2033gat));
OR2X1 g7206(.A (n_2065), .B (n_65), .Y (n_66));
AND2X1 g8109(.A (n3095gat), .B (n3087gat), .Y (n_218));
CLKBUFX1 g8158(.A (n3095gat), .Y (n_278));
INVX1 g8170(.A (n_170), .Y (n_129));
DFFSRX1 n842gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3073gat), .Q (), .QN (n842gat));
DFFSRX1 n2266gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n_20), .Q (n2266gat), .QN ());
INVX1 g8209(.A (n_174), .Y (n_177));
DFFSRX1 n846gat_reg(.RN (1'b1), .SN (n_1165), .CK (blif_clk_net), .D(n3071gat), .Q (n_2002), .QN ());
AND2X1 g8107(.A (n2506gat), .B (n2588gat), .Y (n_55));
INVX1 g8149(.A (n_90), .Y (n_171));
INVX1 g8219(.A (n_1504), .Y (n_420));
INVX2 g8210(.A (n_253), .Y (n_174));
INVX1 g8023(.A (n_50), .Y (n_266));
INVX1 g8171(.A (n_65), .Y (n_170));
INVX1 g8245(.A (n_1525), .Y (n_85));
AND2X1 g7935(.A (n2403gat), .B (n2347gat), .Y (n_398));
INVX1 g8155(.A (n_1526), .Y (n_80));
INVX1 g8217(.A (n_63), .Y (n_143));
INVX1 g8166(.A (n3106gat), .Y (n_1056));
INVX1 g8247(.A (n_1647), .Y (n_251));
NOR2X1 g8129(.A (n3092gat), .B (n3091gat), .Y (n_320));
CLKBUFX1 g7219(.A (n_153), .Y (n_157));
INVX1 g8255(.A (n_142), .Y (n_26));
INVX1 g8236(.A (n_95), .Y (n_145));
NOR2X1 g8126(.A (n2407gat), .B (n2347gat), .Y (n_175));
NOR2X1 g7900(.A (n2394gat), .B (n2403gat), .Y (n_73));
INVX1 g8151(.A (n2495gat), .Y (n_20));
INVX1 g8263(.A (n3066gat), .Y (n_44));
INVX1 g7476(.A (n614gat), .Y (n_42));
INVX1 g8228(.A (n3127gat), .Y (n_31));
INVX1 g8172(.A (n2490gat), .Y (n_65));
INVX1 g8251(.A (n2640gat), .Y (n_18));
INVX1 g8269(.A (n3067gat), .Y (n_36));
INVX1 g8273(.A (n3098gat), .Y (n_15));
INVX1 g8282(.A (n2021gat), .Y (n_13));
INVX1 g8272(.A (n1316gat), .Y (n_12));
INVX1 g8174(.A (n3068gat), .Y (n_38));
INVX1 g8238(.A (n3083gat), .Y (n_135));
INVX1 g8211(.A (n2562gat), .Y (n_253));
INVX1 g8241(.A (n2347gat), .Y (n_72));
INVX1 g8261(.A (n820gat), .Y (n_10));
INVX1 g8163(.A (n830gat), .Y (n_9));
INVX1 g8157(.A (n2037gat), .Y (n_8));
INVX1 g8024(.A (n2403gat), .Y (n_50));
INVX1 g8038(.A (n2190gat), .Y (n_27));
INVX1 g8259(.A (n3084gat), .Y (n_51));
INVX2 g8237(.A (n2203gat), .Y (n_95));
INVX2 g8150(.A (n2626gat), .Y (n_90));
INVX1 g8212(.A (n2562gat), .Y (n_5));
INVX1 g8283(.A (n3094gat), .Y (n_421));
INVX1 g7220(.A (n2543gat), .Y (n_153));
INVX1 g8256(.A (n2394gat), .Y (n_142));
INVX1 g8257(.A (n2394gat), .Y (n_4));
INVX1 g8223(.A (n2634gat), .Y (n_3));
INVX1 g8287(.A (n699gat), .Y (n_21));
INVX1 g8271(.A (n3065gat), .Y (n_46));
INVX1 g8147(.A (n1740gat), .Y (n_2));
INVX1 g8199(.A (blif_reset_net), .Y (n_1165));
INVX1 g8218(.A (n2440gat), .Y (n_63));
INVX1 g8197(.A (n834gat), .Y (n_23));
INVX1 g7891(.A (n1312gat), .Y (n_1));
INVX1 g8161(.A (n152gat), .Y (n_0));
INVX1 g8201(.A (n3126gat), .Y (n_54));
INVX1 g8198(.A (n3100gat), .Y (n_281));
CLKBUFX1 g8455(.A (n_1262), .Y (n_1191));
INVX1 g8457(.A (n_1966), .Y (n_1196));
INVX2 g8458(.A (n_1014), .Y (n_1197));
INVX1 g8459(.A (n_1201), .Y (n_1198));
CLKBUFX1 g8462(.A (n_1885), .Y (n_1201));
INVX1 g8466(.A (n_1734), .Y (n_1208));
INVX1 g8470(.A (n_1837), .Y (n_1211));
INVX1 g52(.A (n_1936), .Y (n_1262));
INVX1 g62(.A (n_1792), .Y (n_1253));
NOR2X1 g65(.A (n_1754), .B (n_13), .Y (n_1259));
INVX1 g29(.A (n3088gat), .Y (n_1267));
NAND2X1 g24_dup(.A (n_1506), .B (n_1528), .Y (n_1272));
INVX1 g28(.A (n3095gat), .Y (n_1268));
NAND2X1 g26(.A (n_51), .B (n_135), .Y (n_1269));
NOR2X1 g8496(.A (n_1275), .B (n_1276), .Y (n_1277));
AOI21X1 g8497(.A0 (n_1078), .A1 (n_1081), .B0 (n_1088), .Y (n_1275));
NAND3X1 g8498(.A (n_1096), .B (n_1089), .C (n_1082), .Y (n_1276));
AND2X1 g8502(.A (n673gat), .B (n_1056), .Y (n_1282));
NOR2X1 g8503(.A (n_612), .B (n_868), .Y (n_1283));
NOR2X1 g44(.A (n_787), .B (n_400), .Y (n_1289));
NOR2X1 g40(.A (n_1294), .B (n_1796), .Y (n_1295));
OR2X1 g42(.A (n_1289), .B (n_1799), .Y (n_1294));
NAND2X1 g8517(.A (n_1310), .B (n_1510), .Y (n_1699));
INVX1 g8518(.A (n_2083), .Y (n_1310));
NAND2X1 g8525(.A (n_1819), .B (n_131), .Y (n_1326));
INVX1 g8533(.A (n_1338), .Y (n_1339));
NAND3X1 g8534(.A (n_1443), .B (n_1337), .C (n_398), .Y (n_1338));
NOR2X1 g8535(.A (n_251), .B (n_159), .Y (n_1337));
NAND3X1 g55(.A (n_1419), .B (n_1431), .C (n_1510), .Y (n_1342));
NAND2X1 g8536(.A (n_1343), .B (n_1419), .Y (n_1344));
INVX1 g8537(.A (n_1860), .Y (n_1343));
NAND2X1 g25_dup(.A (n_1905), .B (n_1702), .Y (n_1345));
NAND3X1 g8542(.A (n_1443), .B (n_1354), .C (n_1362), .Y (n_1363));
AND2X1 g47(.A (n_398), .B (n_228), .Y (n_1354));
NOR2X1 g8549(.A (n2407gat), .B (n_2083), .Y (n_1362));
NAND2X1 g8554(.A (n_1548), .B (n2102gat), .Y (n_1366));
NAND3X1 g8556(.A (n_1371), .B (n_1573), .C (n_1547), .Y (n_1373));
INVX1 g8557(.A (n_1708), .Y (n_1371));
NOR2X1 g8562(.A (n_2121), .B (n_2120), .Y (n_1376));
NAND3X1 g33(.A (n_122), .B (n_261), .C (n_1377), .Y (n_1378));
AND2X1 g8563(.A (n_749), .B (n_153), .Y (n_1377));
NAND2X1 g31(.A (n_165), .B (n_1381), .Y (n_1382));
INVX1 g34(.A (n_1380), .Y (n_1381));
NAND3X1 g35(.A (n_1483), .B (n_95), .C (n2562gat), .Y (n_1380));
CLKBUFX1 g8566(.A (n_2069), .Y (n_1396));
INVX1 g8568(.A (n_1669), .Y (n_1397));
NOR2X1 g8569(.A (n_1398), .B (n_219), .Y (n_1399));
NAND2X1 g8570(.A (n3088gat), .B (n3087gat), .Y (n_1398));
NOR2X1 g32_dup(.A (n_1596), .B (n_1595), .Y (n_1402));
NAND2X1 g8586(.A (n_1862), .B (n_1419), .Y (n_1420));
NOR2X1 g8588(.A (n_251), .B (n_2085), .Y (n_1419));
NAND2X1 g8589(.A (n_1339), .B (n_2086), .Y (n_1421));
AND2X1 g8596(.A (n_1430), .B (n_1453), .Y (n_1431));
NOR2X1 g8597(.A (n_1514), .B (n_1464), .Y (n_1430));
INVX2 g8598(.A (n_1442), .Y (n_1443));
NAND2X1 g8599(.A (n_1901), .B (n_1464), .Y (n_1442));
NAND2X2 g8615(.A (n_1551), .B (n_457), .Y (n_1550));
NAND2X1 g8616(.A (n_2069), .B (n_2051), .Y (n_1216));
NOR2X1 g8619(.A (n_2083), .B (n_1901), .Y (n_1453));
INVX1 g8625(.A (n_1891), .Y (n_1464));
NAND2X1 g8645(.A (n_1382), .B (n_1483), .Y (n_1485));
INVX1 g8647(.A (n2207gat), .Y (n_1483));
AND2X1 g8648(.A (n_271), .B (n_96), .Y (n_1486));
INVX1 g8650(.A (n_1493), .Y (n_1494));
CLKBUFX1 g8651(.A (n_1483), .Y (n_1493));
NOR2X1 g16(.A (n388gat), .B (n_2051), .Y (n_1497));
INVX1 g8654(.A (n331gat), .Y (n_1498));
CLKBUFX1 g8658(.A (n_1886), .Y (n_1504));
INVX1 g8660(.A (n3086gat), .Y (n_1505));
NAND2X1 g8661(.A (n_1506), .B (n_1528), .Y (n_1508));
NOR2X1 g8662(.A (n_1269), .B (n_1268), .Y (n_1506));
NOR2X1 g8664(.A (n_1513), .B (n_1514), .Y (n_1515));
NAND2X1 g24(.A (n_1510), .B (n_1891), .Y (n_1513));
NOR2X1 g8665(.A (n2403gat), .B (n_72), .Y (n_1510));
NAND2X1 g25(.A (n_142), .B (n_143), .Y (n_1514));
AND2X1 g8670(.A (n2343gat), .B (n2399gat), .Y (n_2067));
INVX1 g8671(.A (n2343gat), .Y (n_1525));
INVX1 g8672(.A (n2399gat), .Y (n_1526));
AND2X1 g8673(.A (n_1527), .B (n1871gat), .Y (n_1528));
INVX1 g8674(.A (n3085gat), .Y (n_1527));
INVX1 g8682(.A (n_1547), .Y (n_1544));
INVX1 g8683(.A (n_1547), .Y (n_1546));
CLKBUFX3 g8684(.A (n_1548), .Y (n_1547));
INVX2 g8686(.A (n_1884), .Y (n_1551));
INVX1 g8687(.A (n_1928), .Y (n_1552));
CLKBUFX1 g8695(.A (n_1751), .Y (n_1559));
INVX1 g8699(.A (n_165), .Y (n_1566));
INVX1 g8707(.A (n_1573), .Y (n_1577));
INVX1 g8709(.A (n_1580), .Y (n_1573));
CLKBUFX3 g8710(.A (n_1581), .Y (n_1580));
OR2X1 g8715(.A (n_1588), .B (n_1508), .Y (n_1589));
NAND3X1 g27(.A (n3086gat), .B (n3088gat), .C (n3094gat), .Y (n_1588));
NAND2X1 g8718(.A (n_422), .B (n_1590), .Y (n_1591));
INVX2 g8719(.A (n_1272), .Y (n_1590));
NAND3X1 g8720(.A (n_1593), .B (n_1590), .C (n_1594), .Y (n_1595));
INVX1 g8721(.A (n_1508), .Y (n_1593));
NOR2X1 g8722(.A (n_1267), .B (n_1505), .Y (n_1594));
NAND2X1 g8723(.A (n_422), .B (n3094gat), .Y (n_1596));
NOR2X1 g30(.A (n_1505), .B (n_1597), .Y (n_1598));
INVX1 g8724(.A (n_1593), .Y (n_1597));
NOR2X1 g8725(.A (n_1267), .B (n_1599), .Y (n_1600));
INVX1 g8726(.A (n_1590), .Y (n_1599));
INVX1 g8733(.A (n_1967), .Y (n_1607));
NAND2X2 g8735(.A (n_1610), .B (n_1612), .Y (n_1613));
NAND3X1 g23(.A (n_1609), .B (n_565), .C (n_452), .Y (n_1610));
NAND2X1 g8736(.A (n_1608), .B (n_681), .Y (n_1609));
OR2X1 g8737(.A (n_1924), .B (n_689), .Y (n_1608));
NAND2X1 g8738(.A (n_690), .B (n_1611), .Y (n_1612));
NAND2X1 g8739(.A (n_565), .B (n_452), .Y (n_1611));
NAND2X1 g8745(.A (n_1793), .B (n_106), .Y (n_1621));
INVX1 g8757(.A (n_1926), .Y (n_1637));
INVX1 g8764(.A (n_1814), .Y (n_1646));
INVX1 g8765(.A (n2407gat), .Y (n_1647));
NAND3X1 g8766(.A (n_1648), .B (n_1652), .C (n_2096), .Y (n_1653));
NAND2X1 g8767(.A (n_1824), .B (n3076gat), .Y (n_1648));
NAND2X1 g8768(.A (n_1651), .B (n3067gat), .Y (n_1652));
INVX4 g8769(.A (n_1650), .Y (n_1651));
NAND2X2 g8770(.A (n_2096), .B (n_277), .Y (n_1650));
NAND2X1 g8775(.A (n_1749), .B (n_1715), .Y (n_1658));
NAND4X1 g8778(.A (n_1659), .B (n_836), .C (n_857), .D (n_834), .Y(n_1660));
AND2X1 g8779(.A (n_878), .B (n_864), .Y (n_1659));
NAND2X1 g54(.A (n_894), .B (n_892), .Y (n_1661));
AND2X1 g51(.A (n_1282), .B (n2592gat), .Y (n_1664));
NAND3X1 g8781(.A (n1871gat), .B (n_1668), .C (n3093gat), .Y (n_1669));
AND2X1 g8783(.A (n_51), .B (n_135), .Y (n_1668));
INVX1 g8784(.A (n_1668), .Y (n_1670));
INVX1 g8785(.A (n1871gat), .Y (n3106gat));
NAND4X1 g8791(.A (n_1683), .B (n_1684), .C (n_1685), .D (n_1686), .Y(n_1687));
OR2X1 g8792(.A (n816gat), .B (n3149gat), .Y (n_1683));
INVX2 g8795(.A (n_1905), .Y (n_1680));
NAND2X1 g8798(.A (n3149gat), .B (n957gat), .Y (n_1684));
NOR2X1 g8799(.A (n_95), .B (n_1493), .Y (n_1685));
NOR2X1 g8800(.A (n_253), .B (n_254), .Y (n_1686));
INVX4 g8801(.A (n_1680), .Y (n3149gat));
NAND2X1 g8807(.A (n_1761), .B (n_1784), .Y (n_1702));
OR2X1 g13(.A (n_1759), .B (n_1707), .Y (n_1708));
NAND2X1 g14_dup(.A (n_1751), .B (n1850gat), .Y (n_1707));
NAND3X1 g8811(.A (n_1830), .B (n_1718), .C (n_1719), .Y (n_1720));
INVX1 g8816(.A (n_2094), .Y (n_1715));
NAND2X1 g8819(.A (n_1824), .B (n3077gat), .Y (n_1718));
NAND2X2 g8820(.A (n3068gat), .B (n_1651), .Y (n_1719));
NAND2X1 g8821(.A (n_1729), .B (n_1732), .Y (n_1733));
AOI21X1 g8822(.A0 (n_705), .A1 (n_1721), .B0 (n_1728), .Y (n_1729));
NAND2X1 g8823(.A (n_1498), .B (n_1497), .Y (n_1721));
NAND2X1 g8824(.A (n_1726), .B (n_1727), .Y (n_1728));
OR2X1 g8825(.A (n_1721), .B (n_1725), .Y (n_1726));
NAND2X1 g57(.A (n_2101), .B (n_1724), .Y (n_1725));
NOR2X1 g58(.A (n327gat), .B (n384gat), .Y (n_1724));
NAND2X1 g8827(.A (n_1872), .B (n3078gat), .Y (n_1727));
AOI21X1 g56(.A0 (n_1208), .A1 (n_1730), .B0 (n_1731), .Y (n_1732));
AND2X1 g59(.A (n384gat), .B (n327gat), .Y (n_1730));
AND2X1 g64(.A (n_1871), .B (n3069gat), .Y (n_1731));
INVX1 g60(.A (n_2101), .Y (n_1734));
CLKBUFX1 g8837(.A (n_1749), .Y (n_1748));
INVX2 g8838(.A (n_2072), .Y (n_1749));
NAND4X1 g8839(.A (n_1753), .B (n_1756), .C (n_1757), .D (n_1758), .Y(n_1761));
NOR2X1 g8840(.A (n_1580), .B (n_1752), .Y (n_1753));
NAND2X1 g8841(.A (n_1751), .B (n1850gat), .Y (n_1752));
INVX2 g8842(.A (n_1562), .Y (n_1751));
NAND2X2 g8843(.A (n_1754), .B (n_1755), .Y (n_1756));
INVX2 g8844(.A (n1880gat), .Y (n_1754));
INVX1 g8845(.A (n1763gat), .Y (n_1755));
INVX1 g8846(.A (n_1366), .Y (n_1757));
INVX1 g8848(.A (n_1758), .Y (n_1759));
INVX2 g8849(.A (n1899gat), .Y (n_1758));
INVX1 g8850(.A (n_1759), .Y (n_1241));
INVX1 g8854(.A (n1767gat), .Y (n_1766));
NAND2X1 g8855(.A (n_1761), .B (n_1784), .Y (n_1770));
AND2X1 g8856(.A (n_880), .B (n_1777), .Y (n_1995));
NAND4X1 g8858(.A (n_199), .B (n_1963), .C (n2037gat), .D (n2095gat),.Y (n_1771));
AOI21X1 g36_dup(.A0 (n_2021), .A1 (n_1775), .B0 (n_1776), .Y(n_1777));
NOR2X1 g8860(.A (n_1774), .B (n_412), .Y (n_1775));
NAND2X1 g8861(.A (n_63), .B (n_175), .Y (n_1774));
NOR2X1 g8862(.A (n_627), .B (n_2021), .Y (n_1776));
AOI21X1 g8863(.A0 (n_2027), .A1 (n_1775), .B0 (n_1776), .Y (n_1779));
NAND2X2 g8864(.A (n_1888), .B (n_2030), .Y (n_1784));
NAND2X2 g8868(.A (n_1756), .B (n2102gat), .Y (n_2030));
NAND2X1 g8869(.A (n_1787), .B (n_1789), .Y (n_1790));
AOI21X1 g8870(.A0 (n_1786), .A1 (n830gat), .B0 (n_444), .Y (n_1787));
INVX1 g8871(.A (n_1785), .Y (n_1786));
NAND2X1 g8872(.A (n_2004), .B (n_367), .Y (n_1785));
AOI21X1 g8873(.A0 (n_387), .A1 (n830gat), .B0 (n_1788), .Y (n_1789));
NOR2X1 g8874(.A (n830gat), .B (n_344), .Y (n_1788));
NAND2X1 g17(.A (n_1792), .B (n_1793), .Y (n_1794));
NAND2X2 g8877(.A (n_791), .B (n_515), .Y (n_1792));
OR2X1 g8878(.A (n_1345), .B (n_1363), .Y (n_1793));
INVX2 g8879(.A (n_1801), .Y (n_1802));
NAND3X1 g8880(.A (n_1797), .B (n_1798), .C (n_1800), .Y (n_1801));
INVX1 g8881(.A (n_1796), .Y (n_1797));
NAND2X2 g8882(.A (n_789), .B (n_598), .Y (n_1796));
NOR2X1 g8883(.A (n_1771), .B (n_1289), .Y (n_1798));
INVX1 g8884(.A (n_1799), .Y (n_1800));
NOR2X1 g8885(.A (n_314), .B (n_788), .Y (n_1799));
NAND3X1 g8886(.A (n_1807), .B (n_1810), .C (n_1811), .Y (n_1812));
NAND3X1 g8887(.A (n_1803), .B (n_1878), .C (n463gat), .Y (n_1807));
NAND2X1 g39(.A (n_547), .B (n_1571), .Y (n_1803));
NAND2X1 g8890(.A (n_1808), .B (n_1809), .Y (n_1810));
INVX1 g38(.A (n_1803), .Y (n_1808));
NOR2X1 g8891(.A (n463gat), .B (n_1877), .Y (n_1809));
AOI22X1 g37(.A0 (n3082gat), .A1 (n_1872), .B0 (n_1871), .B1(n3073gat), .Y (n_1811));
NOR2X1 g8892(.A (n_1816), .B (n_1818), .Y (n_1819));
NAND2X1 g8893(.A (n_1905), .B (n_1646), .Y (n_1816));
OR2X1 g8896(.A (n_63), .B (n_4), .Y (n_1814));
INVX1 g8897(.A (n_1904), .Y (n_1818));
NAND3X1 g8900(.A (n_1821), .B (n_1825), .C (n_1828), .Y (n_1829));
NAND2X1 g8901(.A (n_1651), .B (n3066gat), .Y (n_1821));
NAND2X1 g22(.A (n_1824), .B (n3075gat), .Y (n_1825));
INVX4 g8902(.A (n_1823), .Y (n_1824));
NAND2X2 g8903(.A (n_1658), .B (n3095gat), .Y (n_1823));
INVX1 g8904(.A (n_1827), .Y (n_1828));
INVX2 g8905(.A (n_1826), .Y (n_1827));
NAND2X1 g8906(.A (n_1715), .B (n_1749), .Y (n_1826));
INVX4 g8907(.A (n_1827), .Y (n_1830));
NAND4X1 g8908(.A (n_1981), .B (n_2043), .C (n_197), .D (n919gat), .Y(n_1834));
AND2X1 g8909(.A (n_1852), .B (n_2002), .Y (n_1981));
NAND2X1 g8913(.A (n_197), .B (n_2035), .Y (n_1837));
OR2X1 g46(.A (n2407gat), .B (n_1814), .Y (n_1842));
NAND2X1 g8917(.A (n_1892), .B (n_398), .Y (n_1843));
NOR2X1 g8922(.A (n_1920), .B (n_1637), .Y (n_1851));
INVX1 g8923(.A (n2454gat), .Y (n_1852));
NAND2X1 g8925(.A (n_1851), .B (n_1852), .Y (n_2051));
NAND2X1 g8926(.A (n_2116), .B (n_1860), .Y (n_1862));
NAND3X1 g8927(.A (n_1857), .B (n_342), .C (n_1859), .Y (n_1860));
INVX1 g8928(.A (n_1699), .Y (n_1857));
NOR2X1 g8929(.A (n_130), .B (n_1902), .Y (n_1859));
NAND2X1 g8931(.A (n_1515), .B (n_1453), .Y (n_2116));
NAND2X1 g8932(.A (n_1870), .B (n_1873), .Y (n_1874));
NAND2X1 g8933(.A (n_1864), .B (n_2101), .Y (n_1870));
OAI21X1 g8934(.A0 (n_2055), .A1 (n388gat), .B0 (n_1571), .Y (n_1864));
AOI22X1 g8940(.A0 (n3072gat), .A1 (n_1871), .B0 (n_1872), .B1(n3081gat), .Y (n_1873));
CLKBUFX1 g8941(.A (n_2100), .Y (n_1871));
CLKBUFX1 g8942(.A (n_2097), .Y (n_1872));
INVX1 g8943(.A (n_1871), .Y (n_1875));
INVX1 g8944(.A (n_1877), .Y (n_1878));
INVX1 g8945(.A (n_2101), .Y (n_1877));
NAND2X1 g14(.A (n_1882), .B (n_1927), .Y (n_1884));
NOR2X1 g15(.A (n_2044), .B (n_1881), .Y (n_1882));
INVX1 g8948(.A (n402gat), .Y (n_1881));
NOR2X1 g8950(.A (n_1885), .B (n_1887), .Y (n_1888));
NAND2X1 g8951(.A (n_1758), .B (n_1581), .Y (n_1885));
NAND3X1 g8952(.A (n_1886), .B (n_1548), .C (n_1562), .Y (n_1887));
INVX2 g8953(.A (n1850gat), .Y (n_1886));
AND2X1 g43(.A (n_2041), .B (n_1647), .Y (n_1889));
NOR2X1 g8955(.A (n_1894), .B (n_1895), .Y (n_1896));
NAND4X1 g36(.A (n_1902), .B (n_2083), .C (n_1510), .D (n_1893), .Y(n_1894));
INVX1 g8956(.A (n_1892), .Y (n_1893));
INVX2 g8957(.A (n_1891), .Y (n_1892));
INVX1 g8958(.A (n_1926), .Y (n_1891));
INVX1 g8960(.A (n_1819), .Y (n_1895));
INVX1 g8961(.A (n_1893), .Y (n_1898));
NAND4X1 g8963(.A (n_1903), .B (n_1906), .C (n_1907), .D (n_1908), .Y(n_1909));
AND2X1 g8964(.A (n_2083), .B (n_1902), .Y (n_1903));
INVX2 g8966(.A (n_1901), .Y (n_1902));
NOR2X1 g8967(.A (n919gat), .B (n_2043), .Y (n_1901));
AND2X1 g8968(.A (n_1904), .B (n_1905), .Y (n_1906));
NAND2X1 g8969(.A (n_1784), .B (n_1761), .Y (n_1904));
NAND2X2 g8970(.A (n_638), .B (n_1766), .Y (n_1905));
INVX1 g8971(.A (n_1842), .Y (n_1907));
INVX1 g8972(.A (n_1843), .Y (n_1908));
NAND2X1 g21(.A (n_1913), .B (n_1915), .Y (n_1916));
OAI21X1 g8973(.A0 (n_1396), .A1 (n_1912), .B0 (n470gat), .Y (n_1913));
AOI21X1 g8975(.A0 (n_0), .A1 (n256gat), .B0 (n156gat), .Y (n_1912));
NAND2X1 g8977(.A (n_1914), .B (n_549), .Y (n_1915));
NOR2X1 g8978(.A (n470gat), .B (n_1912), .Y (n_1914));
NAND2X1 g8979(.A (n156gat), .B (n_549), .Y (n_1917));
NAND3X1 g8980(.A (n_1918), .B (n_1919), .C (n_1923), .Y (n_1924));
NAND2X1 g8981(.A (n_385), .B (n842gat), .Y (n_1918));
OR2X1 g8982(.A (n842gat), .B (n_1785), .Y (n_1919));
AOI21X1 g8983(.A0 (n_1922), .A1 (n842gat), .B0 (n_436), .Y (n_1923));
INVX1 g8984(.A (n_1920), .Y (n_1922));
NAND2X1 g8986(.A (n919gat), .B (n_2002), .Y (n_1920));
NAND2X1 g8987(.A (n_1926), .B (n_1927), .Y (n_1928));
NOR2X1 g8988(.A (n402gat), .B (n_2044), .Y (n_1926));
INVX2 g8990(.A (n919gat), .Y (n_1927));
NAND4X1 g8991(.A (n_1930), .B (n_1932), .C (n_1933), .D (n_1935), .Y(n_1936));
AOI21X1 g8992(.A0 (n_1889), .A1 (n_1896), .B0 (n_1929), .Y (n_1930));
INVX1 g8993(.A (n_2088), .Y (n_1929));
NOR2X1 g8994(.A (n_1931), .B (n_1621), .Y (n_1932));
NAND2X1 g47_dup(.A (n_1326), .B (n_1909), .Y (n_1931));
AND2X1 g8995(.A (n_1344), .B (n_1421), .Y (n_1933));
NOR2X1 g45(.A (n_1253), .B (n_1934), .Y (n_1935));
INVX1 g48(.A (n_1342), .Y (n_1934));
NAND2X1 g8996(.A (n_1326), .B (n_1909), .Y (n_1937));
NAND2X2 g8997(.A (n_1154), .B (n_1158), .Y (n_1938));
NAND2X1 g6967_dup(.A (n_1154), .B (n_1158), .Y (n_1939));
XOR2X1 g20(.A (n_1947), .B (n_1949), .Y (n_1950));
INVX1 g9005(.A (n256gat), .Y (n_1947));
NOR2X1 g9006(.A (n_1948), .B (n_1396), .Y (n_1949));
OR2X1 g9007(.A (n152gat), .B (n156gat), .Y (n_1948));
NOR2X1 g9008(.A (n_1396), .B (n156gat), .Y (n_1951));
NAND4X1 g9014(.A (n_1959), .B (n_1961), .C (n_1962), .D (n_1965), .Y(n_1966));
CLKBUFX1 g50(.A (n_1958), .Y (n_1959));
NOR2X1 g9015(.A (n_1937), .B (n_1957), .Y (n_1958));
INVX1 g9016(.A (n_1420), .Y (n_1957));
CLKBUFX1 g9017(.A (n_1960), .Y (n_1961));
AOI21X1 g9018(.A0 (n_1896), .A1 (n_1889), .B0 (n_1794), .Y (n_1960));
AND2X1 g9019(.A (n_1421), .B (n_2088), .Y (n_1962));
AND2X1 g9020(.A (n_1963), .B (n_1964), .Y (n_1965));
NAND2X1 g9021(.A (n_786), .B (n_281), .Y (n_1963));
AND2X1 g9022(.A (n2169gat), .B (n1312gat), .Y (n_1964));
NAND3X1 g9023(.A (n_1958), .B (n_1962), .C (n_1960), .Y (n_1967));
INVX2 g9041(.A (n777gat), .Y (n_1990));
INVX2 g9043(.A (n_1995), .Y (n_1992));
CLKBUFX1 g9044(.A (n_1995), .Y (n_1994));
INVX1 g9049(.A (n_2004), .Y (n_2003));
INVX2 g9050(.A (n_2002), .Y (n_2004));
CLKBUFX2 g9053(.A (n_2008), .Y (n_2007));
CLKBUFX2 g9054(.A (n_2004), .Y (n_2008));
INVX1 g9059(.A (n_1373), .Y (n_2014));
INVX1 g9063(.A (n_2021), .Y (n_2019));
INVX1 g9065(.A (n_2024), .Y (n_2022));
INVX4 g9069(.A (n_2027), .Y (n_2024));
CLKBUFX3 g9070(.A (n_2021), .Y (n_2027));
CLKBUFX3 g9071(.A (n_2029), .Y (n_2021));
INVX2 g9072(.A (n_2015), .Y (n_2029));
CLKBUFX3 g9073(.A (n_2030), .Y (n_2015));
INVX1 g9074(.A (n_2032), .Y (n_2031));
CLKBUFX1 g9075(.A (n_2033), .Y (n_2032));
INVX1 g9077(.A (n_2041), .Y (n_2035));
CLKBUFX1 g9083(.A (n_2042), .Y (n_2041));
INVX2 g9084(.A (n_2043), .Y (n_2042));
CLKBUFX3 g9085(.A (n_2044), .Y (n_2043));
INVX2 g9086(.A (n398gat), .Y (n_2044));
INVX1 g9088(.A (n_2048), .Y (n_2046));
CLKBUFX1 g9090(.A (n_2049), .Y (n_2048));
INVX1 g9091(.A (n2622gat), .Y (n_2049));
INVX1 g9092(.A (n_2051), .Y (n_2050));
INVX1 g9096(.A (n_2056), .Y (n_2055));
CLKBUFX1 g9097(.A (n_2051), .Y (n_2056));
INVX1 g9099(.A (n_2063), .Y (n_2059));
CLKBUFX1 g9103(.A (n_2064), .Y (n_2063));
CLKBUFX1 g9104(.A (n_2065), .Y (n_2064));
INVX1 g9105(.A (n2630gat), .Y (n_2065));
CLKBUFX1 g9106(.A (n_2067), .Y (n_2066));
NOR2X1 g9107(.A (n_2068), .B (n_2071), .Y (n_2072));
NAND2X1 g18_dup(.A (n_1550), .B (n_1834), .Y (n_2068));
NAND2X1 g17_dup(.A (n_2069), .B (n_2070), .Y (n_2071));
NAND2X2 g9108(.A (n_1552), .B (n_457), .Y (n_2069));
NAND2X1 g9109(.A (n_1851), .B (n_1852), .Y (n_2070));
NAND2X1 g9110(.A (n_2069), .B (n_2070), .Y (n_2119));
NAND2X1 g18(.A (n_1550), .B (n_1834), .Y (n_2074));
XOR2X1 g9111(.A (n1197gat), .B (n3116gat), .Y (n_2082));
MX2X1 g9112(.A (n_2076), .B (n_2079), .S0 (n_2080), .Y (n3116gat));
MX2X1 g9113(.A (n_1092), .B (n_2075), .S0 (n_1091), .Y (n_2076));
INVX1 g9114(.A (n_1092), .Y (n_2075));
NAND2X1 g9115(.A (n_2078), .B (n_1084), .Y (n_2079));
NAND2X1 g9116(.A (n_2077), .B (n_2075), .Y (n_2078));
INVX1 g41(.A (n_1091), .Y (n_2077));
AOI21X1 g9117(.A0 (n_1009), .A1 (n1045gat), .B0 (n_1034), .Y(n_2080));
NAND4X1 g9118(.A (n_2086), .B (n_2087), .C (n_382), .D (n_343), .Y(n_2088));
NOR2X1 g9119(.A (n_2084), .B (n_2085), .Y (n_2086));
INVX1 g9120(.A (n_2083), .Y (n_2084));
NAND2X2 g9121(.A (n_2042), .B (n_2004), .Y (n_2083));
NAND2X1 g9122(.A (n_1770), .B (n_1905), .Y (n_2085));
AND2X1 g9123(.A (n_1337), .B (n_1510), .Y (n_2087));
NAND2X2 g9124(.A (n_2089), .B (n_2095), .Y (n_2096));
OR2X1 g9125(.A (n_2119), .B (n_2074), .Y (n_2089));
INVX1 g9126(.A (n_2094), .Y (n_2095));
NAND2X1 g9127(.A (n_2090), .B (n_2093), .Y (n_2094));
NOR2X1 g9128(.A (n_1485), .B (n_1486), .Y (n_2090));
NAND2X1 g9129(.A (n_2091), .B (n_1378), .Y (n_2093));
INVX1 g9130(.A (n_1376), .Y (n_2091));
NOR2X1 g9132(.A (n_2097), .B (n_2100), .Y (n_2101));
NOR2X1 g9133(.A (n_1589), .B (n_1591), .Y (n_2097));
AND2X1 g9134(.A (n_2098), .B (n_2099), .Y (n_2100));
NOR2X1 g9135(.A (n_320), .B (n_1669), .Y (n_2098));
AND2X1 g9136(.A (n_116), .B (n_173), .Y (n_2099));
NAND3X1 g9137(.A (n_2106), .B (n_2107), .C (n_2108), .Y (n_2109));
NAND2X1 g9138(.A (n_2102), .B (n_2104), .Y (n_2106));
NAND2X1 g9139(.A (n_1277), .B (n_1167), .Y (n_2102));
CLKBUFX1 g9141(.A (n_2103), .Y (n_2104));
NAND2X1 g9142(.A (n_527), .B (n_487), .Y (n_2103));
OAI21X1 g9143(.A0 (n_1661), .A1 (n_1660), .B0 (n1389gat), .Y(n_2107));
NOR2X1 g9144(.A (n_1664), .B (n_1283), .Y (n_2108));
AOI21X1 g9149(.A0 (n_1397), .A1 (n_1399), .B0 (n_1402), .Y (n_2117));
AOI21X1 g8567_dup(.A0 (n_1397), .A1 (n_1399), .B0 (n_1402), .Y(n_2118));
endmodule
