module des_area(desOut, desIn, kcy1, kcy2, kcy3, decrypt, roundSel, clk, d_out_1, q_in_1, d_out_2, q_in_2, d_out_3, q_in_3, d_out_4, q_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, q_in_7, d_out_8, q_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, d_out_12, q_in_12, d_out_13, q_in_13, d_out_14, q_in_14, d_out_15, q_in_15, d_out_16, q_in_16, d_out_17, q_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, q_in_20, d_out_21, q_in_21, d_out_22, q_in_22, d_out_23, q_in_23, d_out_24, q_in_24, d_out_25, q_in_25, d_out_26, q_in_26, d_out_27, q_in_27, d_out_28, q_in_28, d_out_29, q_in_29, d_out_30, q_in_30, d_out_31, q_in_31, d_out_32, q_in_32, d_out_33, q_in_33, d_out_34, q_in_34, d_out_35, q_in_35, d_out_36, q_in_36, d_out_37, q_in_37, d_out_38, q_in_38, d_out_39, q_in_39, d_out_40, q_in_40, d_out_41, q_in_41, d_out_42, q_in_42, d_out_43, q_in_43, d_out_44, q_in_44, d_out_45, q_in_45, d_out_46, q_in_46, d_out_47, q_in_47, d_out_48, q_in_48, d_out_49, qn_in_49, d_out_50, q_in_50, d_out_51, qn_in_51, d_out_52, q_in_52, d_out_53, q_in_53, d_out_54, q_in_54, d_out_55, q_in_55, d_out_56, q_in_56, d_out_57, q_in_57, d_out_58, q_in_58, d_out_59, qn_in_59, d_out_60, q_in_60, d_out_61, q_in_61, d_out_62, q_in_62, d_out_63, q_in_63, d_out_64, q_in_64, d_out_65, q_in_65, d_out_66, q_in_66, d_out_67, q_in_67, d_out_68, q_in_68, d_out_69, q_in_69, d_out_70, q_in_70, d_out_71, q_in_71, d_out_72, q_in_72, d_out_73, q_in_73, d_out_74, q_in_74, d_out_75, q_in_75, d_out_76, q_in_76, d_out_77, q_in_77, d_out_78, q_in_78, d_out_79, q_in_79, d_out_80, q_in_80, d_out_81, q_in_81, d_out_82, q_in_82, d_out_83, q_in_83, d_out_84, q_in_84, d_out_85, q_in_85, d_out_86, q_in_86, d_out_87, q_in_87, d_out_88, q_in_88, d_out_89, q_in_89, d_out_90, q_in_90, d_out_91, q_in_91, d_out_92, q_in_92, d_out_93, q_in_93, d_out_94, q_in_94, d_out_95, q_in_95, d_out_96, q_in_96, d_out_97, q_in_97, d_out_98, q_in_98, d_out_99, q_in_99, d_out_100, q_in_100, d_out_101, q_in_101, d_out_102, q_in_102, d_out_103, q_in_103, d_out_104, q_in_104, d_out_105, q_in_105, d_out_106, q_in_106, d_out_107, q_in_107, d_out_108, q_in_108, d_out_109, q_in_109, d_out_110, q_in_110, d_out_111, q_in_111, d_out_112, q_in_112, d_out_113, q_in_113, d_out_114, q_in_114, d_out_115, q_in_115, d_out_116, q_in_116, d_out_117, q_in_117, d_out_118, q_in_118, d_out_119, qn_in_119, d_out_120, q_in_120, d_out_121, q_in_121, d_out_122, q_in_122, d_out_123, q_in_123, d_out_124, q_in_124, d_out_125, q_in_125, d_out_126, q_in_126, d_out_127, q_in_127, d_out_128, q_in_128);
input q_in_124;
input q_in_123;
input q_in_122;
input q_in_87;
input q_in_86;
input q_in_85;
input q_in_84;
input q_in_121;
input q_in_81;
input qn_in_49;
input q_in_120;
input qn_in_119;
input q_in_118;
input q_in_117;
input q_in_79;
input q_in_78;
input q_in_77;
input q_in_115;
input q_in_76;
input q_in_116;
input q_in_114;
input q_in_113;
input q_in_112;
input q_in_111;
input q_in_110;
input q_in_109;
input q_in_108;
input q_in_107;
input q_in_106;
input q_in_105;
input q_in_104;
input q_in_103;
input q_in_102;
input q_in_101;
input q_in_100;
input q_in_99;
input q_in_98;
input q_in_97;
input q_in_96;
input q_in_95;
input q_in_94;
input q_in_93;
input q_in_92;
input q_in_91;
input q_in_90;
input q_in_89;
input q_in_88;
input q_in_64;
input q_in_63;
input q_in_62;
input q_in_61;
input q_in_60;
input qn_in_59;
input q_in_128;
input q_in_127;
input q_in_58;
input q_in_57;
input q_in_56;
input q_in_55;
input q_in_54;
input q_in_53;
input q_in_52;
input qn_in_51;
input q_in_83;
input q_in_82;
input q_in_50;
input q_in_80;
input q_in_48;
input q_in_47;
input q_in_46;
input q_in_45;
input q_in_44;
input q_in_43;
input q_in_42;
input q_in_41;
input q_in_40;
input q_in_39;
input q_in_38;
input q_in_37;
input q_in_36;
input q_in_35;
input q_in_34;
input q_in_33;
input q_in_32;
input q_in_31;
input q_in_30;
input q_in_29;
input q_in_28;
input q_in_27;
input q_in_26;
input q_in_25;
input q_in_24;
input q_in_23;
input q_in_22;
input q_in_21;
input q_in_20;
input q_in_19;
input q_in_18;
input q_in_17;
input q_in_16;
input q_in_15;
input q_in_14;
input q_in_13;
input q_in_12;
input q_in_11;
input q_in_10;
input q_in_9;
input q_in_8;
input q_in_7;
input q_in_6;
input q_in_5;
input q_in_4;
input q_in_3;
input q_in_2;
input q_in_1;
input q_in_75;
input q_in_74;
input q_in_73;
input q_in_72;
input q_in_71;
input q_in_70;
input q_in_69;
input q_in_68;
input q_in_67;
input q_in_66;
input q_in_65;
input q_in_126;
input q_in_125;
input [5:0] roundSel;
input decrypt, clk;
input [55:0] kcy1, kcy2, kcy3;
input [63:0] desIn;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_121;
output d_out_81;
output d_out_80;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_115;
output d_out_76;
output d_out_116;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_111;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_64;
output d_out_63;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_128;
output d_out_127;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_83;
output d_out_82;
output d_out_50;
output d_out_49;
output d_out_48;
output d_out_47;
output d_out_46;
output d_out_45;
output d_out_44;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_30;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_5;
output d_out_4;
output d_out_3;
output d_out_2;
output d_out_1;
output d_out_75;
output d_out_74;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_126;
output d_out_125;
output [63:0] desOut;
wire n_7908;
wire n_7900, n_7901, n_7902, n_7903, n_7904, n_7905, n_7906, n_7907;
wire n_7890, n_7891, n_7892, n_7893, n_7894, n_7897, n_7898, n_7899;
wire n_7869, n_7871, n_7884, n_7885, n_7886, n_7887, n_7888, n_7889;
wire n_7821, n_7824, n_7846, n_7854, n_7857, n_7858, n_7859, n_7867;
wire n_7807, n_7808, n_7812, n_7813, n_7815, n_7816, n_7819, n_7820;
wire n_7799, n_7800, n_7801, n_7802, n_7803, n_7804, n_7805, n_7806;
wire n_7790, n_7791, n_7793, n_7794, n_7795, n_7796, n_7797, n_7798;
wire n_7782, n_7783, n_7784, n_7785, n_7786, n_7787, n_7788, n_7789;
wire n_7774, n_7775, n_7776, n_7777, n_7778, n_7779, n_7780, n_7781;
wire n_7754, n_7755, n_7756, n_7757, n_7758, n_7760, n_7762, n_7763;
wire n_7728, n_7732, n_7733, n_7735, n_7738, n_7740, n_7741, n_7753;
wire n_7704, n_7705, n_7706, n_7707, n_7709, n_7711, n_7712, n_7714;
wire n_7683, n_7684, n_7685, n_7686, n_7688, n_7700, n_7701, n_7702;
wire n_7675, n_7676, n_7677, n_7678, n_7679, n_7680, n_7681, n_7682;
wire n_7655, n_7656, n_7660, n_7661, n_7662, n_7663, n_7664, n_7674;
wire n_7636, n_7637, n_7648, n_7649, n_7650, n_7651, n_7652, n_7653;
wire n_7614, n_7615, n_7627, n_7631, n_7632, n_7633, n_7634, n_7635;
wire n_7600, n_7603, n_7604, n_7605, n_7606, n_7607, n_7608, n_7612;
wire n_7588, n_7589, n_7590, n_7594, n_7596, n_7597, n_7598, n_7599;
wire n_7579, n_7580, n_7581, n_7582, n_7583, n_7585, n_7586, n_7587;
wire n_7542, n_7543, n_7544, n_7546, n_7556, n_7559, n_7563, n_7568;
wire n_7532, n_7535, n_7536, n_7537, n_7538, n_7539, n_7540, n_7541;
wire n_7522, n_7525, n_7526, n_7527, n_7528, n_7529, n_7530, n_7531;
wire n_7511, n_7512, n_7513, n_7516, n_7517, n_7518, n_7520, n_7521;
wire n_7503, n_7504, n_7505, n_7506, n_7507, n_7508, n_7509, n_7510;
wire n_7495, n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502;
wire n_7487, n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494;
wire n_7469, n_7470, n_7479, n_7480, n_7481, n_7483, n_7485, n_7486;
wire n_7460, n_7461, n_7462, n_7463, n_7464, n_7465, n_7466, n_7467;
wire n_7448, n_7449, n_7450, n_7451, n_7453, n_7454, n_7455, n_7458;
wire n_7437, n_7440, n_7441, n_7442, n_7443, n_7445, n_7446, n_7447;
wire n_7428, n_7429, n_7430, n_7431, n_7432, n_7434, n_7435, n_7436;
wire n_7419, n_7420, n_7421, n_7422, n_7423, n_7424, n_7426, n_7427;
wire n_7411, n_7412, n_7413, n_7414, n_7415, n_7416, n_7417, n_7418;
wire n_7403, n_7404, n_7405, n_7406, n_7407, n_7408, n_7409, n_7410;
wire n_7380, n_7381, n_7382, n_7397, n_7399, n_7400, n_7401, n_7402;
wire n_7372, n_7373, n_7374, n_7375, n_7376, n_7377, n_7378, n_7379;
wire n_7360, n_7362, n_7363, n_7364, n_7367, n_7368, n_7369, n_7371;
wire n_7350, n_7351, n_7352, n_7353, n_7354, n_7357, n_7358, n_7359;
wire n_7342, n_7343, n_7344, n_7345, n_7346, n_7347, n_7348, n_7349;
wire n_7334, n_7335, n_7336, n_7337, n_7338, n_7339, n_7340, n_7341;
wire n_7319, n_7320, n_7321, n_7322, n_7323, n_7331, n_7332, n_7333;
wire n_7305, n_7307, n_7308, n_7309, n_7311, n_7314, n_7317, n_7318;
wire n_7294, n_7298, n_7299, n_7300, n_7301, n_7302, n_7303, n_7304;
wire n_7250, n_7251, n_7252, n_7253, n_7284, n_7285, n_7289, n_7290;
wire n_7233, n_7237, n_7239, n_7244, n_7245, n_7247, n_7248, n_7249;
wire n_7221, n_7222, n_7224, n_7225, n_7226, n_7227, n_7228, n_7231;
wire n_7199, n_7200, n_7201, n_7216, n_7217, n_7218, n_7219, n_7220;
wire n_7191, n_7192, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198;
wire n_7182, n_7184, n_7185, n_7186, n_7187, n_7188, n_7189, n_7190;
wire n_7174, n_7175, n_7176, n_7177, n_7178, n_7179, n_7180, n_7181;
wire n_7166, n_7167, n_7168, n_7169, n_7170, n_7171, n_7172, n_7173;
wire n_7153, n_7154, n_7156, n_7157, n_7158, n_7159, n_7161, n_7163;
wire n_7145, n_7146, n_7147, n_7148, n_7149, n_7150, n_7151, n_7152;
wire n_7128, n_7129, n_7130, n_7131, n_7133, n_7141, n_7142, n_7144;
wire n_7119, n_7120, n_7121, n_7122, n_7124, n_7125, n_7126, n_7127;
wire n_7095, n_7110, n_7111, n_7112, n_7113, n_7114, n_7117, n_7118;
wire n_7082, n_7086, n_7087, n_7088, n_7090, n_7091, n_7092, n_7093;
wire n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081;
wire n_7050, n_7061, n_7062, n_7068, n_7069, n_7071, n_7072, n_7073;
wire n_7040, n_7041, n_7042, n_7043, n_7044, n_7045, n_7048, n_7049;
wire n_7020, n_7021, n_7022, n_7023, n_7024, n_7026, n_7028, n_7037;
wire n_6997, n_6998, n_6999, n_7002, n_7004, n_7006, n_7018, n_7019;
wire n_6987, n_6988, n_6989, n_6990, n_6991, n_6992, n_6993, n_6994;
wire n_6975, n_6976, n_6978, n_6980, n_6983, n_6984, n_6985, n_6986;
wire n_6963, n_6964, n_6965, n_6966, n_6968, n_6969, n_6972, n_6974;
wire n_6943, n_6944, n_6956, n_6957, n_6959, n_6960, n_6961, n_6962;
wire n_6923, n_6928, n_6930, n_6931, n_6935, n_6936, n_6940, n_6942;
wire n_6904, n_6905, n_6906, n_6909, n_6911, n_6912, n_6913, n_6914;
wire n_6880, n_6881, n_6882, n_6886, n_6888, n_6890, n_6891, n_6903;
wire n_6868, n_6869, n_6872, n_6873, n_6874, n_6875, n_6876, n_6878;
wire n_6847, n_6848, n_6851, n_6852, n_6853, n_6857, n_6865, n_6866;
wire n_6838, n_6840, n_6841, n_6842, n_6843, n_6844, n_6845, n_6846;
wire n_6827, n_6828, n_6829, n_6830, n_6831, n_6832, n_6833, n_6837;
wire n_6818, n_6819, n_6820, n_6821, n_6822, n_6823, n_6824, n_6826;
wire n_6797, n_6799, n_6800, n_6801, n_6802, n_6805, n_6816, n_6817;
wire n_6786, n_6788, n_6789, n_6790, n_6792, n_6794, n_6795, n_6796;
wire n_6775, n_6776, n_6777, n_6779, n_6780, n_6781, n_6782, n_6783;
wire n_6749, n_6750, n_6751, n_6752, n_6753, n_6757, n_6758, n_6759;
wire n_6738, n_6740, n_6741, n_6742, n_6743, n_6744, n_6746, n_6748;
wire n_6703, n_6705, n_6706, n_6707, n_6725, n_6726, n_6727, n_6728;
wire n_6692, n_6693, n_6694, n_6696, n_6697, n_6698, n_6699, n_6700;
wire n_6676, n_6677, n_6679, n_6680, n_6684, n_6686, n_6689, n_6690;
wire n_6643, n_6647, n_6648, n_6660, n_6661, n_6673, n_6674, n_6675;
wire n_6614, n_6615, n_6621, n_6635, n_6636, n_6638, n_6639, n_6640;
wire n_6604, n_6605, n_6607, n_6609, n_6610, n_6611, n_6612, n_6613;
wire n_6594, n_6596, n_6597, n_6598, n_6599, n_6600, n_6602, n_6603;
wire n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592, n_6593;
wire n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6585;
wire n_6567, n_6570, n_6572, n_6573, n_6574, n_6575, n_6576, n_6577;
wire n_6540, n_6541, n_6558, n_6559, n_6560, n_6562, n_6563, n_6564;
wire n_6532, n_6533, n_6534, n_6535, n_6536, n_6537, n_6538, n_6539;
wire n_6502, n_6504, n_6511, n_6526, n_6528, n_6529, n_6530, n_6531;
wire n_6481, n_6485, n_6486, n_6488, n_6491, n_6495, n_6500, n_6501;
wire n_6473, n_6474, n_6475, n_6476, n_6477, n_6478, n_6479, n_6480;
wire n_6464, n_6466, n_6467, n_6468, n_6469, n_6470, n_6471, n_6472;
wire n_6441, n_6450, n_6451, n_6454, n_6457, n_6458, n_6461, n_6463;
wire n_6420, n_6421, n_6430, n_6431, n_6432, n_6435, n_6436, n_6437;
wire n_6406, n_6412, n_6414, n_6415, n_6416, n_6417, n_6418, n_6419;
wire n_6393, n_6394, n_6395, n_6400, n_6402, n_6403, n_6404, n_6405;
wire n_6384, n_6385, n_6386, n_6387, n_6388, n_6389, n_6390, n_6391;
wire n_6375, n_6376, n_6377, n_6378, n_6379, n_6381, n_6382, n_6383;
wire n_6360, n_6361, n_6362, n_6363, n_6371, n_6372, n_6373, n_6374;
wire n_6347, n_6350, n_6351, n_6352, n_6354, n_6355, n_6358, n_6359;
wire n_6335, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344;
wire n_6326, n_6327, n_6328, n_6329, n_6331, n_6332, n_6333, n_6334;
wire n_6316, n_6317, n_6320, n_6321, n_6322, n_6323, n_6324, n_6325;
wire n_6297, n_6298, n_6299, n_6301, n_6302, n_6306, n_6307, n_6311;
wire n_6285, n_6286, n_6287, n_6288, n_6289, n_6290, n_6291, n_6296;
wire n_6276, n_6277, n_6278, n_6279, n_6281, n_6282, n_6283, n_6284;
wire n_6267, n_6268, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275;
wire n_6242, n_6243, n_6244, n_6262, n_6263, n_6264, n_6265, n_6266;
wire n_6222, n_6224, n_6225, n_6226, n_6227, n_6228, n_6229, n_6241;
wire n_6208, n_6209, n_6212, n_6215, n_6216, n_6217, n_6220, n_6221;
wire n_6191, n_6192, n_6195, n_6197, n_6198, n_6199, n_6206, n_6207;
wire n_6181, n_6182, n_6183, n_6184, n_6186, n_6187, n_6188, n_6190;
wire n_6171, n_6172, n_6174, n_6175, n_6176, n_6178, n_6179, n_6180;
wire n_6161, n_6162, n_6163, n_6164, n_6165, n_6167, n_6168, n_6169;
wire n_6136, n_6137, n_6151, n_6153, n_6154, n_6156, n_6159, n_6160;
wire n_6117, n_6118, n_6119, n_6120, n_6121, n_6129, n_6130, n_6132;
wire n_6096, n_6097, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105;
wire n_6086, n_6088, n_6089, n_6090, n_6091, n_6092, n_6094, n_6095;
wire n_6062, n_6065, n_6070, n_6081, n_6082, n_6083, n_6084, n_6085;
wire n_6048, n_6049, n_6050, n_6052, n_6053, n_6056, n_6058, n_6060;
wire n_6022, n_6023, n_6025, n_6027, n_6040, n_6043, n_6044, n_6047;
wire n_6013, n_6014, n_6015, n_6016, n_6017, n_6018, n_6019, n_6020;
wire n_5993, n_5995, n_5996, n_6007, n_6009, n_6010, n_6011, n_6012;
wire n_5968, n_5969, n_5970, n_5971, n_5974, n_5975, n_5977, n_5992;
wire n_5927, n_5929, n_5931, n_5935, n_5938, n_5948, n_5966, n_5967;
wire n_5892, n_5895, n_5897, n_5898, n_5908, n_5912, n_5921, n_5924;
wire n_5713, n_5722, n_5726, n_5732, n_5835, n_5836, n_5838, n_5891;
wire n_5697, n_5698, n_5699, n_5703, n_5704, n_5707, n_5708, n_5711;
wire n_5684, n_5686, n_5687, n_5690, n_5691, n_5694, n_5695, n_5696;
wire n_5667, n_5668, n_5669, n_5676, n_5677, n_5678, n_5680, n_5681;
wire n_5651, n_5652, n_5655, n_5658, n_5659, n_5662, n_5663, n_5666;
wire n_5639, n_5640, n_5641, n_5642, n_5645, n_5646, n_5647, n_5648;
wire n_5616, n_5617, n_5620, n_5624, n_5627, n_5628, n_5631, n_5632;
wire n_5596, n_5597, n_5598, n_5601, n_5609, n_5610, n_5612, n_5613;
wire n_5542, n_5543, n_5544, n_5551, n_5553, n_5590, n_5591, n_5592;
wire n_5523, n_5524, n_5525, n_5526, n_5528, n_5529, n_5532, n_5540;
wire n_5467, n_5472, n_5480, n_5481, n_5483, n_5487, n_5496, n_5516;
wire n_5433, n_5440, n_5443, n_5444, n_5445, n_5447, n_5457, n_5464;
wire n_5411, n_5412, n_5417, n_5419, n_5425, n_5426, n_5428, n_5430;
wire n_5389, n_5391, n_5392, n_5400, n_5402, n_5403, n_5404, n_5407;
wire n_5370, n_5372, n_5375, n_5376, n_5377, n_5379, n_5386, n_5387;
wire n_5355, n_5356, n_5361, n_5363, n_5364, n_5365, n_5366, n_5369;
wire n_5339, n_5340, n_5345, n_5347, n_5349, n_5350, n_5351, n_5354;
wire n_5320, n_5324, n_5325, n_5327, n_5329, n_5331, n_5332, n_5333;
wire n_5302, n_5304, n_5306, n_5307, n_5308, n_5311, n_5316, n_5319;
wire n_5285, n_5287, n_5288, n_5290, n_5291, n_5293, n_5296, n_5300;
wire n_5273, n_5275, n_5277, n_5278, n_5279, n_5280, n_5283, n_5284;
wire n_5261, n_5262, n_5263, n_5265, n_5266, n_5267, n_5269, n_5272;
wire n_5243, n_5245, n_5249, n_5251, n_5252, n_5254, n_5255, n_5260;
wire n_5231, n_5234, n_5236, n_5237, n_5238, n_5239, n_5241, n_5242;
wire n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5230;
wire n_5212, n_5213, n_5214, n_5216, n_5218, n_5219, n_5220, n_5221;
wire n_5194, n_5197, n_5198, n_5201, n_5202, n_5203, n_5207, n_5209;
wire n_5181, n_5184, n_5185, n_5187, n_5188, n_5189, n_5191, n_5193;
wire n_5169, n_5170, n_5171, n_5172, n_5173, n_5176, n_5178, n_5180;
wire n_5161, n_5162, n_5163, n_5164, n_5165, n_5166, n_5167, n_5168;
wire n_5149, n_5150, n_5151, n_5154, n_5155, n_5157, n_5158, n_5160;
wire n_5134, n_5136, n_5138, n_5140, n_5141, n_5142, n_5144, n_5147;
wire n_5119, n_5121, n_5124, n_5126, n_5129, n_5131, n_5132, n_5133;
wire n_5105, n_5106, n_5108, n_5111, n_5112, n_5113, n_5114, n_5118;
wire n_5096, n_5097, n_5099, n_5100, n_5101, n_5102, n_5103, n_5104;
wire n_5077, n_5081, n_5082, n_5083, n_5084, n_5089, n_5092, n_5095;
wire n_5060, n_5062, n_5065, n_5067, n_5068, n_5070, n_5072, n_5075;
wire n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5058, n_5059;
wire n_5039, n_5040, n_5041, n_5042, n_5044, n_5045, n_5048, n_5049;
wire n_5029, n_5030, n_5032, n_5034, n_5035, n_5036, n_5037, n_5038;
wire n_5017, n_5018, n_5019, n_5020, n_5024, n_5025, n_5026, n_5028;
wire n_5005, n_5008, n_5010, n_5012, n_5013, n_5014, n_5015, n_5016;
wire n_4995, n_4996, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004;
wire n_4980, n_4981, n_4982, n_4983, n_4986, n_4988, n_4989, n_4994;
wire n_4965, n_4966, n_4967, n_4969, n_4973, n_4975, n_4976, n_4977;
wire n_4954, n_4955, n_4956, n_4957, n_4959, n_4960, n_4963, n_4964;
wire n_4942, n_4943, n_4944, n_4947, n_4948, n_4949, n_4950, n_4952;
wire n_4934, n_4935, n_4936, n_4937, n_4938, n_4939, n_4940, n_4941;
wire n_4925, n_4926, n_4927, n_4928, n_4930, n_4931, n_4932, n_4933;
wire n_4909, n_4912, n_4918, n_4919, n_4920, n_4921, n_4923, n_4924;
wire n_4894, n_4896, n_4900, n_4902, n_4903, n_4904, n_4907, n_4908;
wire n_4884, n_4885, n_4886, n_4888, n_4889, n_4891, n_4892, n_4893;
wire n_4871, n_4872, n_4873, n_4875, n_4876, n_4877, n_4880, n_4883;
wire n_4863, n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870;
wire n_4850, n_4853, n_4854, n_4856, n_4858, n_4859, n_4861, n_4862;
wire n_4841, n_4842, n_4843, n_4844, n_4845, n_4846, n_4847, n_4849;
wire n_4833, n_4834, n_4835, n_4836, n_4837, n_4838, n_4839, n_4840;
wire n_4825, n_4826, n_4827, n_4828, n_4829, n_4830, n_4831, n_4832;
wire n_4814, n_4815, n_4817, n_4818, n_4819, n_4821, n_4823, n_4824;
wire n_4803, n_4804, n_4807, n_4808, n_4809, n_4810, n_4812, n_4813;
wire n_4788, n_4791, n_4795, n_4796, n_4797, n_4799, n_4800, n_4801;
wire n_4778, n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4787;
wire n_4768, n_4769, n_4770, n_4772, n_4773, n_4774, n_4775, n_4777;
wire n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766, n_4767;
wire n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758, n_4759;
wire n_4739, n_4740, n_4741, n_4743, n_4744, n_4745, n_4747, n_4750;
wire n_4729, n_4730, n_4732, n_4733, n_4734, n_4736, n_4737, n_4738;
wire n_4719, n_4720, n_4721, n_4723, n_4724, n_4726, n_4727, n_4728;
wire n_4706, n_4708, n_4709, n_4710, n_4711, n_4714, n_4717, n_4718;
wire n_4698, n_4699, n_4700, n_4701, n_4702, n_4703, n_4704, n_4705;
wire n_4689, n_4690, n_4691, n_4692, n_4694, n_4695, n_4696, n_4697;
wire n_4679, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686, n_4687;
wire n_4670, n_4671, n_4672, n_4673, n_4675, n_4676, n_4677, n_4678;
wire n_4661, n_4662, n_4663, n_4665, n_4666, n_4667, n_4668, n_4669;
wire n_4651, n_4652, n_4653, n_4655, n_4656, n_4657, n_4658, n_4660;
wire n_4642, n_4644, n_4645, n_4646, n_4647, n_4648, n_4649, n_4650;
wire n_4632, n_4633, n_4634, n_4635, n_4637, n_4638, n_4639, n_4641;
wire n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4630, n_4631;
wire n_4613, n_4615, n_4616, n_4617, n_4619, n_4620, n_4621, n_4622;
wire n_4603, n_4604, n_4605, n_4606, n_4608, n_4609, n_4610, n_4612;
wire n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602;
wire n_4584, n_4585, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594;
wire n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582;
wire n_4558, n_4561, n_4562, n_4569, n_4570, n_4572, n_4573, n_4574;
wire n_4543, n_4544, n_4545, n_4546, n_4548, n_4549, n_4551, n_4554;
wire n_4533, n_4534, n_4536, n_4537, n_4539, n_4540, n_4541, n_4542;
wire n_4524, n_4525, n_4526, n_4527, n_4528, n_4529, n_4531, n_4532;
wire n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4521, n_4522;
wire n_4501, n_4503, n_4504, n_4508, n_4509, n_4510, n_4511, n_4513;
wire n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498, n_4499;
wire n_4482, n_4485, n_4486, n_4487, n_4488, n_4489, n_4490, n_4491;
wire n_4473, n_4474, n_4476, n_4477, n_4478, n_4479, n_4480, n_4481;
wire n_4464, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471, n_4472;
wire n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4462;
wire n_4443, n_4446, n_4447, n_4449, n_4450, n_4451, n_4452, n_4453;
wire n_4434, n_4435, n_4436, n_4438, n_4439, n_4440, n_4441, n_4442;
wire n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433;
wire n_4414, n_4418, n_4419, n_4420, n_4421, n_4423, n_4424, n_4425;
wire n_4404, n_4405, n_4406, n_4408, n_4409, n_4410, n_4412, n_4413;
wire n_4392, n_4393, n_4394, n_4395, n_4398, n_4399, n_4400, n_4403;
wire n_4381, n_4384, n_4386, n_4387, n_4388, n_4389, n_4390, n_4391;
wire n_4350, n_4356, n_4365, n_4366, n_4368, n_4375, n_4378, n_4380;
wire n_4341, n_4342, n_4343, n_4344, n_4345, n_4346, n_4348, n_4349;
wire n_4333, n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340;
wire n_4323, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330, n_4332;
wire n_4313, n_4314, n_4315, n_4316, n_4317, n_4319, n_4320, n_4322;
wire n_4302, n_4306, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312;
wire n_4286, n_4287, n_4289, n_4293, n_4294, n_4296, n_4300, n_4301;
wire n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4284, n_4285;
wire n_4269, n_4270, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276;
wire n_4257, n_4260, n_4261, n_4262, n_4263, n_4264, n_4267, n_4268;
wire n_4245, n_4247, n_4249, n_4250, n_4252, n_4253, n_4255, n_4256;
wire n_4236, n_4237, n_4238, n_4239, n_4241, n_4242, n_4243, n_4244;
wire n_4223, n_4226, n_4227, n_4228, n_4230, n_4231, n_4233, n_4235;
wire n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220, n_4222;
wire n_4203, n_4204, n_4206, n_4207, n_4210, n_4211, n_4212, n_4213;
wire n_4189, n_4191, n_4193, n_4195, n_4197, n_4198, n_4199, n_4202;
wire n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4187, n_4188;
wire n_4145, n_4158, n_4159, n_4161, n_4164, n_4172, n_4176, n_4177;
wire n_4119, n_4120, n_4124, n_4125, n_4126, n_4133, n_4134, n_4142;
wire n_4107, n_4108, n_4109, n_4111, n_4114, n_4116, n_4117, n_4118;
wire n_4095, n_4096, n_4097, n_4098, n_4099, n_4104, n_4105, n_4106;
wire n_4082, n_4083, n_4088, n_4090, n_4091, n_4092, n_4093, n_4094;
wire n_4069, n_4073, n_4074, n_4075, n_4077, n_4078, n_4079, n_4080;
wire n_4061, n_4062, n_4063, n_4064, n_4065, n_4066, n_4067, n_4068;
wire n_4052, n_4054, n_4055, n_4056, n_4057, n_4058, n_4059, n_4060;
wire n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4049, n_4050;
wire n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041;
wire n_4014, n_4022, n_4025, n_4027, n_4028, n_4029, n_4030, n_4031;
wire n_3982, n_3983, n_3984, n_3985, n_3988, n_3994, n_4012, n_4013;
wire n_3972, n_3973, n_3974, n_3975, n_3976, n_3977, n_3978, n_3980;
wire n_3962, n_3965, n_3966, n_3967, n_3968, n_3969, n_3970, n_3971;
wire n_3948, n_3950, n_3953, n_3954, n_3956, n_3957, n_3958, n_3960;
wire n_3932, n_3934, n_3938, n_3941, n_3942, n_3945, n_3946, n_3947;
wire n_3909, n_3913, n_3919, n_3924, n_3926, n_3929, n_3930, n_3931;
wire n_3890, n_3891, n_3892, n_3893, n_3894, n_3896, n_3897, n_3899;
wire n_3872, n_3873, n_3875, n_3876, n_3879, n_3883, n_3885, n_3887;
wire n_3855, n_3860, n_3861, n_3863, n_3864, n_3865, n_3866, n_3870;
wire n_3829, n_3830, n_3831, n_3832, n_3834, n_3844, n_3850, n_3851;
wire n_3814, n_3815, n_3816, n_3817, n_3818, n_3821, n_3824, n_3827;
wire n_3776, n_3780, n_3786, n_3787, n_3797, n_3798, n_3805, n_3806;
wire n_3759, n_3764, n_3766, n_3768, n_3771, n_3772, n_3774, n_3775;
wire n_3747, n_3748, n_3751, n_3752, n_3754, n_3755, n_3756, n_3758;
wire n_3734, n_3736, n_3737, n_3738, n_3742, n_3744, n_3745, n_3746;
wire n_3721, n_3724, n_3725, n_3729, n_3730, n_3731, n_3732, n_3733;
wire n_3704, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3720;
wire n_3680, n_3681, n_3683, n_3685, n_3691, n_3692, n_3693, n_3695;
wire n_3667, n_3668, n_3669, n_3670, n_3673, n_3675, n_3677, n_3678;
wire n_3645, n_3650, n_3651, n_3654, n_3658, n_3664, n_3665, n_3666;
wire n_3631, n_3634, n_3635, n_3637, n_3638, n_3639, n_3640, n_3641;
wire n_3613, n_3614, n_3617, n_3624, n_3625, n_3628, n_3629, n_3630;
wire n_3593, n_3596, n_3601, n_3602, n_3603, n_3604, n_3608, n_3612;
wire n_3576, n_3578, n_3585, n_3586, n_3587, n_3588, n_3589, n_3592;
wire n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3570, n_3571;
wire n_3550, n_3552, n_3553, n_3554, n_3557, n_3558, n_3560, n_3561;
wire n_3535, n_3536, n_3537, n_3540, n_3541, n_3544, n_3548, n_3549;
wire n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3534;
wire n_3512, n_3513, n_3514, n_3515, n_3516, n_3521, n_3522, n_3524;
wire n_3503, n_3504, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511;
wire n_3485, n_3487, n_3491, n_3492, n_3493, n_3494, n_3498, n_3501;
wire n_3471, n_3472, n_3473, n_3478, n_3479, n_3480, n_3481, n_3483;
wire n_3459, n_3460, n_3462, n_3463, n_3465, n_3466, n_3467, n_3468;
wire n_3446, n_3451, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458;
wire n_3429, n_3430, n_3432, n_3436, n_3440, n_3442, n_3444, n_3445;
wire n_3419, n_3420, n_3421, n_3422, n_3423, n_3425, n_3426, n_3428;
wire n_3405, n_3406, n_3410, n_3411, n_3414, n_3416, n_3417, n_3418;
wire n_3395, n_3397, n_3398, n_3399, n_3400, n_3401, n_3403, n_3404;
wire n_3382, n_3383, n_3387, n_3390, n_3391, n_3392, n_3393, n_3394;
wire n_3358, n_3361, n_3372, n_3377, n_3378, n_3379, n_3380, n_3381;
wire n_3346, n_3349, n_3351, n_3352, n_3354, n_3355, n_3356, n_3357;
wire n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3344, n_3345;
wire n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3329, n_3336;
wire n_3311, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319;
wire n_3301, n_3302, n_3303, n_3304, n_3305, n_3308, n_3309, n_3310;
wire n_3275, n_3276, n_3280, n_3281, n_3282, n_3284, n_3285, n_3287;
wire n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273;
wire n_3247, n_3248, n_3251, n_3252, n_3255, n_3257, n_3258, n_3262;
wire n_3233, n_3234, n_3235, n_3238, n_3240, n_3243, n_3244, n_3245;
wire n_3211, n_3221, n_3223, n_3226, n_3227, n_3228, n_3229, n_3232;
wire n_3201, n_3202, n_3203, n_3204, n_3207, n_3208, n_3209, n_3210;
wire n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, n_3200;
wire n_3183, n_3185, n_3186, n_3188, n_3189, n_3190, n_3191, n_3192;
wire n_3173, n_3174, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181;
wire n_3161, n_3162, n_3164, n_3166, n_3167, n_3168, n_3170, n_3171;
wire n_3151, n_3152, n_3153, n_3154, n_3155, n_3158, n_3159, n_3160;
wire n_3140, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3149;
wire n_3129, n_3130, n_3132, n_3133, n_3134, n_3135, n_3138, n_3139;
wire n_3119, n_3120, n_3121, n_3122, n_3123, n_3125, n_3126, n_3128;
wire n_3107, n_3109, n_3110, n_3112, n_3114, n_3115, n_3116, n_3117;
wire n_3085, n_3090, n_3093, n_3101, n_3103, n_3104, n_3105, n_3106;
wire n_3070, n_3071, n_3074, n_3076, n_3078, n_3080, n_3081, n_3084;
wire n_3057, n_3058, n_3059, n_3060, n_3061, n_3065, n_3067, n_3068;
wire n_3047, n_3048, n_3049, n_3050, n_3051, n_3053, n_3054, n_3056;
wire n_3036, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045;
wire n_3021, n_3026, n_3027, n_3028, n_3029, n_3030, n_3033, n_3035;
wire n_3009, n_3010, n_3011, n_3013, n_3014, n_3015, n_3016, n_3019;
wire n_2997, n_2998, n_2999, n_3000, n_3002, n_3006, n_3007, n_3008;
wire n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995;
wire n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987;
wire n_2965, n_2966, n_2969, n_2970, n_2973, n_2974, n_2977, n_2979;
wire n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2962, n_2964;
wire n_2944, n_2946, n_2947, n_2949, n_2950, n_2952, n_2953, n_2954;
wire n_2930, n_2931, n_2932, n_2935, n_2936, n_2939, n_2941, n_2943;
wire n_2918, n_2921, n_2923, n_2925, n_2926, n_2927, n_2928, n_2929;
wire n_2909, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917;
wire n_2898, n_2899, n_2900, n_2902, n_2903, n_2905, n_2907, n_2908;
wire n_2888, n_2889, n_2891, n_2892, n_2893, n_2895, n_2896, n_2897;
wire n_2874, n_2876, n_2878, n_2879, n_2881, n_2882, n_2883, n_2886;
wire n_2863, n_2864, n_2865, n_2867, n_2868, n_2870, n_2871, n_2872;
wire n_2852, n_2854, n_2855, n_2856, n_2857, n_2859, n_2860, n_2862;
wire n_2840, n_2841, n_2842, n_2843, n_2845, n_2847, n_2848, n_2850;
wire n_2831, n_2832, n_2833, n_2834, n_2836, n_2837, n_2838, n_2839;
wire n_2822, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830;
wire n_2811, n_2812, n_2813, n_2814, n_2815, n_2817, n_2818, n_2819;
wire n_2800, n_2801, n_2802, n_2805, n_2806, n_2807, n_2809, n_2810;
wire n_2790, n_2792, n_2793, n_2794, n_2795, n_2797, n_2798, n_2799;
wire n_2781, n_2782, n_2783, n_2785, n_2786, n_2787, n_2788, n_2789;
wire n_2766, n_2767, n_2769, n_2770, n_2774, n_2776, n_2777, n_2778;
wire n_2753, n_2757, n_2759, n_2761, n_2762, n_2763, n_2764, n_2765;
wire n_2743, n_2744, n_2746, n_2747, n_2748, n_2749, n_2751, n_2752;
wire n_2729, n_2734, n_2735, n_2736, n_2737, n_2738, n_2740, n_2742;
wire n_2719, n_2720, n_2721, n_2723, n_2725, n_2726, n_2727, n_2728;
wire n_2708, n_2709, n_2711, n_2712, n_2713, n_2715, n_2716, n_2717;
wire n_2694, n_2695, n_2699, n_2700, n_2701, n_2702, n_2704, n_2705;
wire n_2682, n_2684, n_2685, n_2686, n_2688, n_2689, n_2692, n_2693;
wire n_2670, n_2671, n_2672, n_2673, n_2674, n_2676, n_2678, n_2680;
wire n_2660, n_2661, n_2662, n_2664, n_2665, n_2666, n_2667, n_2668;
wire n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658;
wire n_2639, n_2640, n_2642, n_2643, n_2644, n_2645, n_2649, n_2650;
wire n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638;
wire n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630;
wire n_2614, n_2615, n_2616, n_2617, n_2619, n_2620, n_2621, n_2622;
wire n_2605, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613;
wire n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2603, n_2604;
wire n_2587, n_2588, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595;
wire n_2578, n_2579, n_2580, n_2581, n_2582, n_2584, n_2585, n_2586;
wire n_2568, n_2569, n_2570, n_2572, n_2573, n_2575, n_2576, n_2577;
wire n_2557, n_2558, n_2559, n_2561, n_2562, n_2564, n_2565, n_2566;
wire n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2555, n_2556;
wire n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546;
wire n_2530, n_2531, n_2532, n_2534, n_2535, n_2536, n_2537, n_2538;
wire n_2517, n_2520, n_2521, n_2522, n_2523, n_2526, n_2528, n_2529;
wire n_2506, n_2507, n_2509, n_2510, n_2511, n_2512, n_2514, n_2516;
wire n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505;
wire n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496;
wire n_2479, n_2480, n_2482, n_2483, n_2484, n_2486, n_2487, n_2488;
wire n_2469, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477;
wire n_2460, n_2461, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468;
wire n_2449, n_2451, n_2453, n_2454, n_2455, n_2456, n_2457, n_2459;
wire n_2439, n_2440, n_2441, n_2443, n_2444, n_2446, n_2447, n_2448;
wire n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438;
wire n_2419, n_2420, n_2422, n_2423, n_2425, n_2427, n_2429, n_2430;
wire n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2415, n_2417;
wire n_2399, n_2400, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407;
wire n_2390, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398;
wire n_2381, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389;
wire n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380;
wire n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2371;
wire n_2353, n_2354, n_2355, n_2356, n_2357, n_2359, n_2361, n_2362;
wire n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351;
wire n_2331, n_2332, n_2334, n_2337, n_2339, n_2340, n_2341, n_2343;
wire n_2318, n_2319, n_2322, n_2324, n_2325, n_2326, n_2329, n_2330;
wire n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317;
wire n_2293, n_2294, n_2298, n_2304, n_2305, n_2306, n_2307, n_2309;
wire n_2281, n_2282, n_2283, n_2284, n_2286, n_2287, n_2289, n_2291;
wire n_2267, n_2269, n_2271, n_2273, n_2275, n_2276, n_2278, n_2280;
wire n_2256, n_2257, n_2258, n_2261, n_2263, n_2264, n_2265, n_2266;
wire n_2246, n_2247, n_2248, n_2249, n_2250, n_2252, n_2253, n_2254;
wire n_2234, n_2236, n_2237, n_2238, n_2239, n_2241, n_2242, n_2245;
wire n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2232, n_2233;
wire n_2215, n_2216, n_2217, n_2218, n_2219, n_2221, n_2222, n_2223;
wire n_2206, n_2207, n_2208, n_2209, n_2211, n_2212, n_2213, n_2214;
wire n_2196, n_2198, n_2199, n_2200, n_2201, n_2203, n_2204, n_2205;
wire n_2184, n_2185, n_2188, n_2190, n_2191, n_2193, n_2194, n_2195;
wire n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183;
wire n_2166, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175;
wire n_2154, n_2155, n_2157, n_2158, n_2159, n_2162, n_2163, n_2165;
wire n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152;
wire n_2135, n_2136, n_2137, n_2138, n_2139, n_2141, n_2143, n_2144;
wire n_2124, n_2125, n_2126, n_2129, n_2130, n_2131, n_2133, n_2134;
wire n_2114, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123;
wire n_2104, n_2105, n_2107, n_2108, n_2109, n_2110, n_2112, n_2113;
wire n_2095, n_2096, n_2097, n_2098, n_2100, n_2101, n_2102, n_2103;
wire n_2084, n_2086, n_2087, n_2089, n_2090, n_2091, n_2092, n_2094;
wire n_2073, n_2074, n_2075, n_2076, n_2078, n_2079, n_2081, n_2083;
wire n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072;
wire n_2055, n_2056, n_2057, n_2058, n_2060, n_2061, n_2063, n_2064;
wire n_2045, n_2046, n_2047, n_2049, n_2050, n_2052, n_2053, n_2054;
wire n_2036, n_2037, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
wire n_2025, n_2027, n_2028, n_2029, n_2030, n_2032, n_2034, n_2035;
wire n_2016, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
wire n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015;
wire n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2007;
wire n_1988, n_1989, n_1991, n_1993, n_1994, n_1995, n_1996, n_1997;
wire n_1977, n_1979, n_1980, n_1982, n_1984, n_1985, n_1986, n_1987;
wire n_1968, n_1969, n_1970, n_1971, n_1972, n_1974, n_1975, n_1976;
wire n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1967;
wire n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957;
wire n_1941, n_1942, n_1943, n_1944, n_1946, n_1947, n_1948, n_1949;
wire n_1930, n_1931, n_1933, n_1935, n_1936, n_1937, n_1939, n_1940;
wire n_1920, n_1921, n_1922, n_1923, n_1924, n_1926, n_1928, n_1929;
wire n_1911, n_1912, n_1913, n_1914, n_1915, n_1917, n_1918, n_1919;
wire n_1885, n_1886, n_1887, n_1888, n_1893, n_1896, n_1897, n_1902;
wire n_1876, n_1877, n_1878, n_1879, n_1880, n_1882, n_1883, n_1884;
wire n_1861, n_1862, n_1863, n_1865, n_1868, n_1869, n_1870, n_1872;
wire n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1858, n_1860;
wire n_1841, n_1842, n_1843, n_1846, n_1847, n_1848, n_1849, n_1850;
wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1830, n_1831, n_1832;
wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
wire n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1814, n_1815;
wire n_1797, n_1798, n_1799, n_1800, n_1802, n_1803, n_1805, n_1806;
wire n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796;
wire n_1779, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
wire n_1768, n_1769, n_1770, n_1771, n_1773, n_1776, n_1777, n_1778;
wire n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1766, n_1767;
wire n_1749, n_1750, n_1751, n_1753, n_1754, n_1755, n_1757, n_1758;
wire n_1739, n_1740, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747;
wire n_1729, n_1730, n_1732, n_1733, n_1734, n_1735, n_1737, n_1738;
wire n_1720, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728;
wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1719;
wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701;
wire n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692;
wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1684;
wire n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1675;
wire n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666;
wire n_1650, n_1651, n_1652, n_1654, n_1655, n_1656, n_1657, n_1658;
wire n_1640, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1649;
wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1638, n_1639;
wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
wire n_1613, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
wire n_1604, n_1605, n_1606, n_1607, n_1608, n_1610, n_1611, n_1612;
wire n_1595, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603;
wire n_1586, n_1587, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594;
wire n_1577, n_1578, n_1579, n_1580, n_1582, n_1583, n_1584, n_1585;
wire n_1568, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576;
wire n_1556, n_1560, n_1561, n_1562, n_1563, n_1564, n_1566, n_1567;
wire n_1545, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554;
wire n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544;
wire n_1527, n_1528, n_1530, n_1531, n_1532, n_1533, n_1534, n_1536;
wire n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1525, n_1526;
wire n_1509, n_1510, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
wire n_1498, n_1499, n_1500, n_1501, n_1502, n_1506, n_1507, n_1508;
wire n_1488, n_1489, n_1490, n_1491, n_1493, n_1495, n_1496, n_1497;
wire n_1478, n_1480, n_1481, n_1482, n_1484, n_1485, n_1486, n_1487;
wire n_1459, n_1464, n_1465, n_1466, n_1469, n_1470, n_1472, n_1475;
wire n_1436, n_1437, n_1442, n_1443, n_1445, n_1449, n_1454, n_1455;
wire n_1422, n_1423, n_1424, n_1427, n_1428, n_1429, n_1433, n_1435;
wire n_1411, n_1413, n_1414, n_1415, n_1416, n_1418, n_1419, n_1420;
wire n_1399, n_1402, n_1403, n_1404, n_1405, n_1406, n_1408, n_1409;
wire n_1389, n_1390, n_1391, n_1393, n_1395, n_1396, n_1397, n_1398;
wire n_1379, n_1380, n_1381, n_1382, n_1384, n_1385, n_1387, n_1388;
wire n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378;
wire n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370;
wire n_1353, n_1355, n_1356, n_1358, n_1359, n_1360, n_1361, n_1362;
wire n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1343, n_1344;
wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1334, n_1335;
wire n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326;
wire n_1302, n_1305, n_1310, n_1311, n_1312, n_1314, n_1316, n_1317;
wire n_1281, n_1284, n_1286, n_1290, n_1291, n_1292, n_1294, n_1300;
wire n_1268, n_1269, n_1271, n_1272, n_1276, n_1277, n_1279, n_1280;
wire n_1253, n_1255, n_1256, n_1258, n_1259, n_1260, n_1264, n_1267;
wire n_1227, n_1228, n_1229, n_1232, n_1233, n_1237, n_1241, n_1251;
wire n_1212, n_1213, n_1215, n_1216, n_1218, n_1219, n_1221, n_1225;
wire n_1195, n_1198, n_1200, n_1201, n_1204, n_1206, n_1208, n_1209;
wire n_1182, n_1183, n_1184, n_1188, n_1190, n_1192, n_1193, n_1194;
wire n_1172, n_1173, n_1174, n_1176, n_1177, n_1178, n_1180, n_1181;
wire n_1163, n_1164, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171;
wire n_1154, n_1155, n_1156, n_1157, n_1158, n_1160, n_1161, n_1162;
wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153;
wire n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145;
wire n_1129, n_1130, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137;
wire n_1109, n_1113, n_1115, n_1116, n_1125, n_1126, n_1127, n_1128;
wire n_1094, n_1099, n_1100, n_1102, n_1103, n_1104, n_1106, n_1107;
wire n_1075, n_1076, n_1081, n_1082, n_1085, n_1088, n_1089, n_1093;
wire n_1056, n_1061, n_1063, n_1064, n_1065, n_1068, n_1070, n_1071;
wire n_1046, n_1047, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054;
wire n_1031, n_1033, n_1034, n_1035, n_1036, n_1038, n_1041, n_1043;
wire n_1015, n_1018, n_1024, n_1025, n_1026, n_1027, n_1028, n_1030;
wire n_999, n_1002, n_1003, n_1004, n_1005, n_1007, n_1013, n_1014;
wire n_988, n_990, n_992, n_993, n_995, n_996, n_997, n_998;
wire n_972, n_973, n_977, n_979, n_980, n_981, n_983, n_985;
wire n_963, n_964, n_965, n_966, n_967, n_968, n_970, n_971;
wire n_951, n_953, n_954, n_955, n_956, n_957, n_958, n_962;
wire n_938, n_939, n_941, n_942, n_943, n_947, n_948, n_950;
wire n_927, n_928, n_929, n_931, n_932, n_934, n_935, n_937;
wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
wire n_902, n_905, n_908, n_909, n_912, n_914, n_915, n_918;
wire n_886, n_887, n_888, n_889, n_891, n_898, n_899, n_901;
wire n_877, n_878, n_879, n_880, n_881, n_883, n_884, n_885;
wire n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_876;
wire n_859, n_860, n_861, n_863, n_864, n_865, n_866, n_867;
wire n_848, n_849, n_852, n_853, n_854, n_855, n_856, n_858;
wire n_836, n_837, n_838, n_839, n_840, n_842, n_843, n_846;
wire n_826, n_827, n_828, n_829, n_831, n_833, n_834, n_835;
wire n_814, n_815, n_817, n_818, n_820, n_821, n_822, n_825;
wire n_798, n_801, n_803, n_808, n_809, n_810, n_811, n_812;
wire n_789, n_790, n_791, n_792, n_793, n_794, n_796, n_797;
wire n_778, n_779, n_781, n_783, n_784, n_785, n_786, n_788;
wire n_767, n_768, n_770, n_772, n_773, n_774, n_775, n_777;
wire n_758, n_759, n_760, n_761, n_763, n_764, n_765, n_766;
wire n_748, n_750, n_751, n_752, n_753, n_754, n_755, n_756;
wire n_736, n_737, n_739, n_741, n_742, n_743, n_744, n_746;
wire n_726, n_728, n_729, n_730, n_731, n_732, n_733, n_735;
wire n_716, n_717, n_719, n_720, n_721, n_722, n_724, n_725;
wire n_701, n_702, n_707, n_709, n_710, n_711, n_714, n_715;
wire n_690, n_692, n_693, n_695, n_696, n_697, n_698, n_700;
wire n_665, n_666, n_675, n_676, n_680, n_684, n_685, n_689;
wire n_652, n_654, n_655, n_657, n_658, n_659, n_662, n_664;
wire n_633, n_634, n_636, n_637, n_639, n_644, n_646, n_649;
wire n_621, n_622, n_623, n_625, n_626, n_627, n_630, n_632;
wire n_611, n_612, n_613, n_614, n_615, n_617, n_618, n_619;
wire n_589, n_592, n_593, n_595, n_601, n_602, n_606, n_610;
wire n_568, n_569, n_570, n_571, n_573, n_574, n_576, n_586;
wire n_549, n_552, n_553, n_556, n_559, n_562, n_563, n_565;
wire n_533, n_534, n_536, n_538, n_539, n_542, n_544, n_548;
wire n_522, n_524, n_525, n_527, n_528, n_529, n_530, n_532;
wire n_509, n_510, n_511, n_512, n_515, n_518, n_520, n_521;
wire n_498, n_500, n_502, n_503, n_504, n_506, n_507, n_508;
wire n_483, n_485, n_487, n_488, n_490, n_493, n_494, n_497;
wire n_467, n_469, n_471, n_472, n_473, n_475, n_476, n_477;
wire n_452, n_454, n_455, n_459, n_460, n_463, n_464, n_466;
wire n_443, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
wire n_430, n_431, n_432, n_434, n_437, n_438, n_439, n_440;
wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_429;
wire n_411, n_413, n_414, n_415, n_416, n_418, n_419, n_420;
wire n_399, n_400, n_401, n_402, n_404, n_405, n_406, n_408;
wire n_387, n_388, n_390, n_391, n_392, n_393, n_397, n_398;
wire n_373, n_375, n_376, n_377, n_379, n_380, n_381, n_386;
wire n_362, n_364, n_365, n_367, n_369, n_370, n_371, n_372;
wire n_346, n_349, n_351, n_355, n_356, n_358, n_359, n_360;
wire n_329, n_332, n_333, n_337, n_338, n_339, n_340, n_341;
wire n_302, n_303, n_315, n_316, n_318, n_320, n_321, n_324;
wire n_281, n_282, n_283, n_290, n_295, n_296, n_297, n_299;
wire n_266, n_269, n_274, n_275, n_276, n_277, n_278, n_280;
wire n_248, n_249, n_253, n_256, n_259, n_260, n_262, n_265;
wire n_233, n_234, n_235, n_239, n_240, n_241, n_243, n_245;
wire n_221, n_223, n_225, n_226, n_227, n_229, n_231, n_232;
wire n_198, n_199, n_200, n_204, n_207, n_215, n_217, n_219;
wire n_177, n_180, n_181, n_183, n_187, n_189, n_191, n_192;
wire n_158, n_159, n_162, n_164, n_170, n_171, n_172, n_174;
wire n_136, n_139, n_140, n_145, n_149, n_155, n_156, n_157;
wire n_126, n_127, n_128, n_129, n_131, n_132, n_133, n_135;
wire n_104, n_105, n_106, n_109, n_113, n_117, n_123, n_124;
wire n_92, n_93, n_95, n_96, n_97, n_99, n_102, n_103;
wire n_83, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
wire n_74, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
wire n_64, n_65, n_66, n_67, n_69, n_70, n_72, n_73;
wire n_52, n_53, n_54, n_56, n_60, n_61, n_62, n_63;
wire n_43, n_45, n_46, n_47, n_48, n_49, n_50, n_51;
wire n_34, n_35, n_37, n_38, n_39, n_40, n_41, n_42;
wire n_24, n_25, n_26, n_27, n_30, n_31, n_32, n_33;
wire n_11, n_12, n_14, n_15, n_17, n_18, n_19, n_23;
wire n_0, n_1, n_5, n_6, n_7, n_8, n_9, n_10;
wire R_118, R_119, R_120, R_121, R_122, R_123, R_124, R_125;
wire R_110, R_111, R_112, R_113, R_114, R_115, R_116, R_117;
wire R_102, R_103, R_104, R_105, R_106, R_107, R_108, R_109;
wire R, R_95, R_96, R_97, R_98, R_99, R_100, R_101;
wire L_87, L_88, L_89, L_90, L_91, L_92, L_93, L_94;
wire L_79, L_80, L_81, L_82, L_83, L_84, L_85, L_86;
wire L_71, L_72, L_73, L_74, L_75, L_76, L_77, L_78;
wire L, L_64, L_65, L_66, L_67, L_68, L_69, L_70;
wire FP_R_56, FP_R_57, FP_R_58, FP_R_59, FP_R_60, FP_R_61, FP_R_62, FP_R_63;
wire FP_R_48, FP_R_49, FP_R_50, FP_R_51, FP_R_52, FP_R_53, FP_R_54, FP_R_55;
wire FP_R_40, FP_R_41, FP_R_42, FP_R_43, FP_R_44, FP_R_45, FP_R_46, FP_R_47;
wire FP_R_32, FP_R_33, FP_R_34, FP_R_35, FP_R_36, FP_R_37, FP_R_38, FP_R_39;
wire FP_R_24, FP_R_25, FP_R_26, FP_R_27, FP_R_28, FP_R_29, FP_R_30, FP_R_31;
wire FP_R_16, FP_R_17, FP_R_18, FP_R_19, FP_R_20, FP_R_21, FP_R_22, FP_R_23;
wire FP_R_8, FP_R_9, FP_R_10, FP_R_11, FP_R_12, FP_R_13, FP_R_14, FP_R_15;
wire FP_R, FP_R_1, FP_R_2, FP_R_3, FP_R_4, FP_R_5, FP_R_6, FP_R_7;
wire [63:0] desOut;
wire [5:0] roundSel;
wire decrypt, clk;
wire [55:0] kcy1, kcy2, kcy3;
wire [63:0] desIn;
CLKBUFX1 gbuf_d_1(.A(desOut[0]), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(FP_R_39));
CLKBUFX1 gbuf_d_2(.A(desOut[0]), .Y(d_out_2));
CLKBUFX1 gbuf_q_2(.A(q_in_2), .Y(R_101));
CLKBUFX1 gbuf_d_3(.A(desOut[20]), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(FP_R_53));
CLKBUFX1 gbuf_d_4(.A(n_7631), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(R_115));
CLKBUFX1 gbuf_d_5(.A(desOut[22]), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(FP_R_61));
CLKBUFX1 gbuf_d_6(.A(desOut[54]), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(R_119));
CLKBUFX1 gbuf_d_7(.A(desOut[54]), .Y(d_out_7));
CLKBUFX1 gbuf_q_7(.A(q_in_7), .Y(FP_R_57));
CLKBUFX1 gbuf_d_8(.A(desOut[22]), .Y(d_out_8));
CLKBUFX1 gbuf_q_8(.A(q_in_8), .Y(R_123));
CLKBUFX1 gbuf_d_9(.A(desOut[52]), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(FP_R_49));
CLKBUFX1 gbuf_d_10(.A(desOut[52]), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(R_111));
CLKBUFX1 gbuf_d_11(.A(desOut[30]), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(FP_R_60));
CLKBUFX1 gbuf_d_12(.A(desOut[30]), .Y(d_out_12));
CLKBUFX1 gbuf_q_12(.A(q_in_12), .Y(R_122));
CLKBUFX1 gbuf_d_13(.A(desOut[32]), .Y(d_out_13));
CLKBUFX1 gbuf_q_13(.A(q_in_13), .Y(FP_R_35));
CLKBUFX1 gbuf_d_14(.A(desOut[32]), .Y(d_out_14));
CLKBUFX1 gbuf_q_14(.A(q_in_14), .Y(R_97));
CLKBUFX1 gbuf_d_15(.A(desOut[42]), .Y(d_out_15));
CLKBUFX1 gbuf_q_15(.A(q_in_15), .Y(FP_R_42));
CLKBUFX1 gbuf_d_16(.A(desOut[42]), .Y(d_out_16));
CLKBUFX1 gbuf_q_16(.A(q_in_16), .Y(R_104));
CLKBUFX1 gbuf_d_17(.A(desOut[44]), .Y(d_out_17));
CLKBUFX1 gbuf_q_17(.A(q_in_17), .Y(R_112));
CLKBUFX1 gbuf_d_18(.A(desOut[14]), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(R_124));
CLKBUFX1 gbuf_d_19(.A(desOut[38]), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(FP_R_59));
CLKBUFX1 gbuf_d_20(.A(desOut[38]), .Y(d_out_20));
CLKBUFX1 gbuf_q_20(.A(q_in_20), .Y(R_121));
CLKBUFX1 gbuf_d_21(.A(desOut[24]), .Y(d_out_21));
CLKBUFX1 gbuf_q_21(.A(q_in_21), .Y(FP_R_36));
CLKBUFX1 gbuf_d_22(.A(desOut[44]), .Y(d_out_22));
CLKBUFX1 gbuf_q_22(.A(q_in_22), .Y(FP_R_50));
CLKBUFX1 gbuf_d_23(.A(desOut[14]), .Y(d_out_23));
CLKBUFX1 gbuf_q_23(.A(q_in_23), .Y(FP_R_62));
CLKBUFX1 gbuf_d_24(.A(desOut[36]), .Y(d_out_24));
CLKBUFX1 gbuf_q_24(.A(q_in_24), .Y(R_113));
CLKBUFX1 gbuf_d_25(.A(desOut[24]), .Y(d_out_25));
CLKBUFX1 gbuf_q_25(.A(q_in_25), .Y(R_98));
CLKBUFX1 gbuf_d_26(.A(n_7546), .Y(d_out_26));
CLKBUFX1 gbuf_q_26(.A(q_in_26), .Y(FP_R_51));
NAND2X2 g13479(.A (n_7762), .B (n_7763), .Y (desOut[54]));
NAND2X2 g13481(.A (n_5551), .B (n_5524), .Y (desOut[22]));
NAND2X2 g13526(.A (n_5544), .B (n_5553), .Y (desOut[52]));
CLKBUFX1 gbuf_d_27(.A(desOut[48]), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(FP_R_33));
CLKBUFX1 gbuf_d_28(.A(desOut[8]), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(R_100));
CLKBUFX1 gbuf_d_29(.A(desOut[62]), .Y(d_out_29));
CLKBUFX1 gbuf_q_29(.A(q_in_29), .Y(FP_R_56));
CLKBUFX1 gbuf_d_30(.A(desOut[26]), .Y(d_out_30));
CLKBUFX1 gbuf_q_30(.A(q_in_30), .Y(FP_R_44));
CLKBUFX1 gbuf_d_31(.A(desOut[48]), .Y(d_out_31));
CLKBUFX1 gbuf_q_31(.A(q_in_31), .Y(R_95));
CLKBUFX1 gbuf_d_32(.A(desOut[26]), .Y(d_out_32));
CLKBUFX1 gbuf_q_32(.A(q_in_32), .Y(R_106));
CLKBUFX1 gbuf_d_33(.A(n_7627), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(R_118));
CLKBUFX1 gbuf_d_34(.A(desOut[28]), .Y(d_out_34));
CLKBUFX1 gbuf_q_34(.A(q_in_34), .Y(FP_R_52));
CLKBUFX1 gbuf_d_35(.A(desOut[28]), .Y(d_out_35));
CLKBUFX1 gbuf_q_35(.A(q_in_35), .Y(R_114));
CLKBUFX1 gbuf_d_36(.A(desOut[8]), .Y(d_out_36));
CLKBUFX1 gbuf_q_36(.A(q_in_36), .Y(FP_R_38));
CLKBUFX1 gbuf_d_37(.A(desOut[16]), .Y(d_out_37));
CLKBUFX1 gbuf_q_37(.A(q_in_37), .Y(FP_R_37));
CLKBUFX1 gbuf_d_38(.A(desOut[18]), .Y(d_out_38));
CLKBUFX1 gbuf_q_38(.A(q_in_38), .Y(FP_R_45));
CLKBUFX1 gbuf_d_39(.A(desOut[12]), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(FP_R_54));
CLKBUFX1 gbuf_d_40(.A(desOut[34]), .Y(d_out_40));
CLKBUFX1 gbuf_q_40(.A(q_in_40), .Y(FP_R_43));
CLKBUFX1 gbuf_d_41(.A(desOut[46]), .Y(d_out_41));
CLKBUFX1 gbuf_q_41(.A(q_in_41), .Y(FP_R_58));
CLKBUFX1 gbuf_d_42(.A(desOut[12]), .Y(d_out_42));
CLKBUFX1 gbuf_q_42(.A(q_in_42), .Y(R_116));
CLKBUFX1 gbuf_d_43(.A(desOut[18]), .Y(d_out_43));
CLKBUFX1 gbuf_q_43(.A(q_in_43), .Y(R_107));
CLKBUFX1 gbuf_d_44(.A(desOut[34]), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(R_105));
CLKBUFX1 gbuf_d_45(.A(n_6880), .Y(d_out_45));
CLKBUFX1 gbuf_q_45(.A(q_in_45), .Y(R_99));
CLKBUFX1 gbuf_d_46(.A(desOut[46]), .Y(d_out_46));
CLKBUFX1 gbuf_q_46(.A(q_in_46), .Y(R_120));
CLKBUFX1 gbuf_d_47(.A(desOut[4]), .Y(d_out_47));
CLKBUFX1 gbuf_q_47(.A(q_in_47), .Y(FP_R_55));
CLKBUFX1 gbuf_d_48(.A(desOut[4]), .Y(d_out_48));
CLKBUFX1 gbuf_q_48(.A(q_in_48), .Y(R_117));
CLKBUFX1 gbuf_d_49(.A(desOut[10]), .Y(d_out_49));
CLKBUFX1 gbuf_qn_49(.A(qn_in_49), .Y(FP_R_46));
CLKBUFX1 gbuf_d_50(.A(n_7660), .Y(d_out_50));
CLKBUFX1 gbuf_q_50(.A(q_in_50), .Y(R_108));
NAND2X2 g13480(.A (n_5525), .B (n_5542), .Y (desOut[24]));
NAND2X2 g13453(.A (n_5496), .B (n_5540), .Y (desOut[42]));
CLKBUFX1 gbuf_d_51(.A(desOut[40]), .Y(d_out_51));
CLKBUFX1 gbuf_qn_51(.A(qn_in_51), .Y(FP_R_34));
CLKBUFX1 gbuf_d_52(.A(desOut[56]), .Y(d_out_52));
CLKBUFX1 gbuf_q_52(.A(q_in_52), .Y(FP_R_32));
CLKBUFX1 gbuf_d_53(.A(desOut[56]), .Y(d_out_53));
CLKBUFX1 gbuf_q_53(.A(q_in_53), .Y(R));
CLKBUFX1 gbuf_d_54(.A(desOut[50]), .Y(d_out_54));
CLKBUFX1 gbuf_q_54(.A(q_in_54), .Y(FP_R_41));
CLKBUFX1 gbuf_d_55(.A(desOut[50]), .Y(d_out_55));
CLKBUFX1 gbuf_q_55(.A(q_in_55), .Y(R_103));
CLKBUFX1 gbuf_d_56(.A(desOut[6]), .Y(d_out_56));
CLKBUFX1 gbuf_q_56(.A(q_in_56), .Y(FP_R_63));
CLKBUFX1 gbuf_d_57(.A(desOut[6]), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(R_125));
CLKBUFX1 gbuf_d_58(.A(desOut[40]), .Y(d_out_58));
CLKBUFX1 gbuf_q_58(.A(q_in_58), .Y(R_96));
NAND2X1 g13537(.A (n_5529), .B (n_3720), .Y (n_5553));
NAND2X2 g13484(.A (n_5481), .B (n_5516), .Y (desOut[12]));
NAND2X1 g13495(.A (n_7199), .B (n_5526), .Y (n_7763));
NAND2X2 g13498(.A (n_6394), .B (n_5523), .Y (n_5551));
CLKBUFX1 gbuf_d_59(.A(desOut[2]), .Y(d_out_59));
CLKBUFX1 gbuf_qn_59(.A(qn_in_59), .Y(FP_R_47));
CLKBUFX1 gbuf_d_60(.A(desOut[2]), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(R_109));
CLKBUFX1 gbuf_d_61(.A(desOut[58]), .Y(d_out_61));
CLKBUFX1 gbuf_q_61(.A(q_in_61), .Y(FP_R_40));
CLKBUFX1 gbuf_d_62(.A(n_7688), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(R_102));
CLKBUFX1 gbuf_d_63(.A(desOut[60]), .Y(d_out_63));
CLKBUFX1 gbuf_q_63(.A(q_in_63), .Y(FP_R_48));
CLKBUFX1 gbuf_d_64(.A(desOut[60]), .Y(d_out_64));
CLKBUFX1 gbuf_q_64(.A(q_in_64), .Y(R_110));
NAND2X1 g13535(.A (n_5528), .B (n_3721), .Y (n_5544));
NAND2X1 g13547(.A (n_5483), .B (n_3670), .Y (n_5543));
NAND2X1 g13497(.A (n_5487), .B (n_3724), .Y (n_5542));
NAND2X1 g13471(.A (n_5472), .B (n_3664), .Y (n_5540));
NAND2X1 g13545(.A (n_6324), .B (n_3669), .Y (n_5532));
NAND2X2 g13558(.A (n_5464), .B (n_5457), .Y (desOut[60]));
INVX1 g13572(.A (n_5528), .Y (n_5529));
OR4X1 g13496(.A (n_5526), .B (n_7193), .C (n_7201), .D (n_7200), .Y(n_7762));
NAND2X1 g13499(.A (n_6378), .B (n_3725), .Y (n_5525));
OR4X1 g13500(.A (n_5523), .B (n_6390), .C (n_5304), .D (n_6395), .Y(n_5524));
NAND2X1 g13504(.A (n_5467), .B (n_3629), .Y (n_5516));
NAND2X1 g13470(.A (n_6333), .B (n_3665), .Y (n_5496));
INVX1 g13551(.A (n_6378), .Y (n_5487));
INVX1 g13568(.A (n_6324), .Y (n_5483));
NAND4X1 g13573(.A (n_7907), .B (n_7908), .C (n_5411), .D (n_5249), .Y(n_5528));
NAND2X1 g13503(.A (n_6789), .B (n_3630), .Y (n_5481));
NAND2X2 g13595(.A (n_7159), .B (n_3675), .Y (n_5480));
INVX1 g13521(.A (n_6333), .Y (n_5472));
INVX1 g13553(.A (n_6789), .Y (n_5467));
NAND2X1 g13566(.A (n_6912), .B (n_3667), .Y (n_5464));
OAI21X1 g13563(.A0 (n_5386), .A1 (n_5077), .B0 (n_5445), .Y (n_6090));
NAND4X1 g13564(.A (n_3666), .B (n_6905), .C (n_6913), .D (n_6914), .Y(n_5457));
NAND2X1 g13609(.A (n_5412), .B (n_5275), .Y (n_5447));
AOI22X1 g13579(.A0 (n_6966), .A1 (n_7544), .B0 (n_5279), .B1(n_7465), .Y (n_5444));
AOI21X1 g13581(.A0 (n_5327), .A1 (n_6786), .B0 (n_5392), .Y (n_5443));
NAND2X1 g13593(.A (n_5387), .B (n_5428), .Y (n_5440));
NAND2X1 g13617(.A (n_5403), .B (n_5445), .Y (n_5698));
AOI22X1 g13532(.A0 (n_6965), .A1 (n_7650), .B0 (n_4960), .B1(n_7464), .Y (n_5433));
OAI21X1 g13571(.A0 (n_5329), .A1 (n_4624), .B0 (n_5426), .Y (n_5430));
AOI21X1 g13580(.A0 (n_5332), .A1 (n_5419), .B0 (n_5319), .Y (n_5425));
NOR2X1 g13612(.A (n_5040), .B (n_5363), .Y (n_5417));
NAND2X1 g13615(.A (n_5377), .B (n_3899), .Y (n_7907));
OAI21X1 g13630(.A0 (n_5339), .A1 (n_4686), .B0 (n_6966), .Y (n_5412));
NOR2X1 g13635(.A (n_4862), .B (n_5379), .Y (n_5411));
NAND2X1 g13669(.A (n_7424), .B (n_6327), .Y (n_5407));
OAI21X1 g13680(.A0 (n_5287), .A1 (n_7173), .B0 (n_5260), .Y (n_5403));
INVX1 g13685(.A (n_5376), .Y (n_5402));
NAND4X1 g13596(.A (n_7537), .B (n_7538), .C (n_5262), .D (n_5272), .Y(n_5400));
AOI22X1 g13605(.A0 (n_5285), .A1 (n_5428), .B0 (n_4429), .B1(n_5144), .Y (n_6089));
NAND4X1 g13620(.A (n_6013), .B (n_5167), .C (n_6014), .D (n_5171), .Y(n_5392));
NAND2X1 g13621(.A (n_5350), .B (n_4356), .Y (n_5391));
NOR2X1 g13627(.A (n_4630), .B (n_5347), .Y (n_5389));
NAND3X1 g13632(.A (n_7529), .B (n_7530), .C (n_5102), .Y (n_5387));
NAND4X1 g13634(.A (n_5680), .B (n_5224), .C (n_5681), .D (n_5254), .Y(n_5386));
AOI21X1 g13665(.A0 (n_7599), .A1 (n_7600), .B0 (n_3899), .Y (n_5379));
NAND4X1 g13681(.A (n_7525), .B (n_4667), .C (n_5099), .D (n_7526), .Y(n_5377));
NAND3X1 g13686(.A (n_5703), .B (n_5704), .C (n_5243), .Y (n_5376));
NOR2X1 g13687(.A (n_4925), .B (n_5302), .Y (n_5375));
NAND2X1 g13689(.A (n_5291), .B (n_7375), .Y (n_5372));
NAND2X1 g13726(.A (n_5290), .B (n_5361), .Y (n_5370));
OAI21X1 g13728(.A0 (n_5284), .A1 (n_4817), .B0 (n_7367), .Y (n_5369));
NAND4X1 g13597(.A (n_5252), .B (n_5131), .C (n_5230), .D (n_4903), .Y(n_7650));
NAND4X1 g13603(.A (n_6868), .B (n_5365), .C (n_6869), .D (n_4924), .Y(n_5366));
OAI21X1 g13623(.A0 (n_5273), .A1 (n_4779), .B0 (n_6209), .Y (n_5364));
AOI21X1 g13628(.A0 (n_4821), .A1 (n_5266), .B0 (n_5419), .Y (n_5363));
NAND4X1 g13637(.A (n_7777), .B (n_7778), .C (n_5209), .D (n_4896), .Y(n_7544));
NAND2X1 g13654(.A (n_5261), .B (n_5265), .Y (n_5356));
NAND3X1 g13657(.A (n_5048), .B (n_5150), .C (n_5219), .Y (n_5355));
AOI21X1 g13659(.A0 (n_4489), .A1 (n_7225), .B0 (n_5263), .Y (n_5354));
NAND2X1 g13661(.A (n_5278), .B (n_7142), .Y (n_5686));
NAND3X1 g13668(.A (n_5201), .B (n_5216), .C (n_5213), .Y (n_5351));
NAND4X1 g13670(.A (n_5035), .B (n_5049), .C (n_5118), .D (n_4818), .Y(n_5350));
NAND4X1 g13672(.A (n_5283), .B (n_5154), .C (n_4954), .D (n_5025), .Y(n_5349));
AOI21X1 g13674(.A0 (n_5197), .A1 (n_5191), .B0 (n_6195), .Y (n_5347));
NOR2X1 g13683(.A (n_5054), .B (n_5277), .Y (n_5345));
NAND3X1 g13706(.A (n_7587), .B (n_7588), .C (n_5068), .Y (n_5340));
NAND3X1 g13709(.A (n_5255), .B (n_5176), .C (n_4581), .Y (n_5339));
NAND3X1 g13613(.A (n_7755), .B (n_4799), .C (n_7756), .Y (n_5333));
NAND4X1 g13624(.A (n_7795), .B (n_7796), .C (n_5038), .D (n_4726), .Y(n_5332));
NAND3X1 g13626(.A (n_4965), .B (n_5227), .C (n_4927), .Y (n_5331));
NAND4X1 g13641(.A (n_7539), .B (n_4631), .C (n_7540), .D (n_4315), .Y(n_5329));
NAND4X1 g13643(.A (n_5155), .B (n_5104), .C (n_5119), .D (n_4655), .Y(n_5327));
NAND4X1 g13644(.A (n_7884), .B (n_6088), .C (n_7885), .D (n_4697), .Y(n_7556));
NAND3X1 g13645(.A (n_5238), .B (n_5198), .C (n_5053), .Y (n_5325));
NAND4X1 g13646(.A (n_5251), .B (n_4800), .C (n_5030), .D (n_4940), .Y(n_5324));
NAND3X1 g13656(.A (n_5097), .B (n_4348), .C (n_5147), .Y (n_5320));
AOI21X1 g13667(.A0 (n_5138), .A1 (n_5100), .B0 (n_4554), .Y (n_5319));
NAND3X1 g13694(.A (n_5178), .B (n_4975), .C (n_4888), .Y (n_5316));
NOR2X1 g13699(.A (n_5222), .B (n_5311), .Y (n_5699));
NAND3X1 g13707(.A (n_5032), .B (n_5072), .C (n_5028), .Y (n_5308));
NAND2X1 g13708(.A (n_4900), .B (n_5207), .Y (n_5307));
AOI21X1 g13713(.A0 (n_5114), .A1 (n_7489), .B0 (n_5404), .Y (n_5306));
INVX1 g13718(.A (n_6391), .Y (n_5304));
NAND3X1 g13720(.A (n_6104), .B (n_6105), .C (n_6993), .Y (n_5302));
NAND2X1 g13729(.A (n_7788), .B (n_7789), .Y (n_5300));
NAND3X1 g13736(.A (n_4891), .B (n_4889), .C (n_5106), .Y (n_5296));
NOR2X1 g13737(.A (n_4518), .B (n_5226), .Y (n_7529));
NAND2X1 g13744(.A (n_5237), .B (n_7173), .Y (n_5293));
NAND3X1 g13746(.A (n_7775), .B (n_7776), .C (n_6451), .Y (n_5291));
NAND2X1 g13747(.A (n_5234), .B (n_4956), .Y (n_5290));
OAI21X1 g13782(.A0 (n_5149), .A1 (n_7490), .B0 (n_5184), .Y (n_5288));
NOR2X1 g13802(.A (n_4703), .B (n_5236), .Y (n_5287));
NAND2X1 g13813(.A (n_5228), .B (n_6151), .Y (n_7538));
NAND2X1 g13653(.A (n_5231), .B (n_4767), .Y (n_5285));
NAND2X1 g13918(.A (n_5060), .B (n_5169), .Y (n_5284));
NAND2X1 g13924(.A (n_4210), .B (n_5160), .Y (n_5283));
OAI21X1 g13676(.A0 (n_4986), .A1 (n_4658), .B0 (n_4554), .Y (n_7908));
NOR2X1 g13691(.A (n_4989), .B (n_5279), .Y (n_5280));
NAND2X1 g13695(.A (n_5136), .B (n_4723), .Y (n_5278));
NAND4X1 g13698(.A (n_5590), .B (n_4350), .C (n_4740), .D (n_5034), .Y(n_5277));
OAI21X1 g13703(.A0 (n_5016), .A1 (n_4950), .B0 (n_7464), .Y (n_5275));
NAND4X1 g13705(.A (n_5895), .B (n_5092), .C (n_4918), .D (n_4529), .Y(n_5273));
NAND2X1 g13714(.A (n_5141), .B (n_6151), .Y (n_5272));
OAI21X1 g13721(.A0 (n_4943), .A1 (n_7122), .B0 (n_4850), .Y (n_5269));
NAND2X1 g13725(.A (n_5103), .B (n_5142), .Y (n_5267));
AOI21X1 g13727(.A0 (n_4967), .A1 (n_5121), .B0 (n_4973), .Y (n_5266));
NOR2X1 g13730(.A (n_4595), .B (n_5126), .Y (n_5265));
AOI21X1 g13740(.A0 (n_4980), .A1 (n_4434), .B0 (n_7122), .Y (n_5263));
NAND3X1 g13742(.A (n_5601), .B (n_6151), .C (n_5203), .Y (n_5262));
NOR2X1 g13750(.A (n_4760), .B (n_5173), .Y (n_5261));
NAND2X1 g13752(.A (n_5075), .B (n_7170), .Y (n_5260));
OAI21X1 g13757(.A0 (n_5058), .A1 (n_4682), .B0 (n_6999), .Y (n_6013));
NAND2X1 g13773(.A (n_5083), .B (n_7237), .Y (n_5255));
NAND2X1 g13776(.A (n_5084), .B (n_7171), .Y (n_5254));
NOR2X1 g13778(.A (n_4868), .B (n_5105), .Y (n_6011));
OAI21X1 g13785(.A0 (n_5005), .A1 (n_7740), .B0 (n_7237), .Y (n_5252));
NAND2X1 g13790(.A (n_5112), .B (n_5938), .Y (n_5251));
NAND2X1 g13804(.A (n_5095), .B (n_5121), .Y (n_5249));
AOI21X1 g13806(.A0 (n_4672), .A1 (n_4854), .B0 (n_5165), .Y (n_6014));
AOI21X1 g13874(.A0 (n_4982), .A1 (n_5041), .B0 (n_3994), .Y (n_5245));
NOR2X1 g13882(.A (n_5164), .B (n_4741), .Y (n_5243));
NAND2X1 g13883(.A (n_5163), .B (n_4727), .Y (n_5242));
NAND2X1 g13897(.A (n_5168), .B (n_7322), .Y (n_5241));
NAND2X1 g13911(.A (n_5036), .B (n_4784), .Y (n_5239));
NAND2X1 g13913(.A (n_5020), .B (n_7237), .Y (n_5238));
NAND2X1 g13914(.A (n_4625), .B (n_5180), .Y (n_5237));
NAND2X1 g13917(.A (n_4549), .B (n_5052), .Y (n_5236));
NOR2X1 g13991(.A (n_4590), .B (n_5000), .Y (n_5234));
OAI21X1 g13693(.A0 (n_4764), .A1 (n_4117), .B0 (n_5225), .Y (n_6868));
OAI21X1 g13716(.A0 (n_4756), .A1 (n_4477), .B0 (n_5935), .Y (n_7755));
OAI21X1 g13717(.A0 (n_4935), .A1 (n_4963), .B0 (n_5214), .Y (n_5231));
OAI21X1 g13722(.A0 (n_4762), .A1 (n_4750), .B0 (n_7463), .Y (n_5230));
AOI21X1 g13731(.A0 (n_4937), .A1 (n_4902), .B0 (n_4584), .Y (n_7777));
NAND2X1 g14119(.A (n_4995), .B (n_5044), .Y (n_5228));
NOR2X1 g13738(.A (n_5065), .B (n_5002), .Y (n_5227));
OAI21X1 g13743(.A0 (n_4928), .A1 (n_5225), .B0 (n_5224), .Y (n_5226));
OAI21X1 g14141(.A0 (n_4145), .A1 (n_4645), .B0 (n_5003), .Y (n_5223));
NAND2X1 g13753(.A (n_4977), .B (n_5220), .Y (n_5222));
NAND2X1 g13755(.A (n_5051), .B (n_5220), .Y (n_5221));
OAI21X1 g13758(.A0 (n_4919), .A1 (n_4183), .B0 (n_3994), .Y (n_5219));
AOI21X1 g13762(.A0 (n_4912), .A1 (n_4761), .B0 (n_4575), .Y (n_5218));
NOR2X1 g13764(.A (n_4930), .B (n_4947), .Y (n_5216));
NAND2X1 g13765(.A (n_4949), .B (n_5214), .Y (n_5680));
NOR2X1 g13766(.A (n_4944), .B (n_4718), .Y (n_5213));
NAND2X1 g13771(.A (n_4941), .B (n_7142), .Y (n_5212));
OAI21X1 g13774(.A0 (n_4695), .A1 (n_4831), .B0 (n_7237), .Y (n_5209));
OAI21X1 g13775(.A0 (n_4886), .A1 (n_4314), .B0 (n_5931), .Y (n_5207));
OAI21X1 g13777(.A0 (n_4670), .A1 (n_4892), .B0 (n_5938), .Y (n_7788));
OAI21X1 g13783(.A0 (n_4827), .A1 (n_5113), .B0 (n_5203), .Y (n_7537));
OAI21X1 g13784(.A0 (n_4830), .A1 (n_5089), .B0 (n_4498), .Y (n_5202));
NOR2X1 g13788(.A (n_4966), .B (n_4734), .Y (n_5201));
OAI21X1 g13789(.A0 (n_4840), .A1 (n_4311), .B0 (n_5948), .Y (n_7756));
OAI21X1 g13791(.A0 (n_4833), .A1 (n_4828), .B0 (n_7465), .Y (n_5198));
AOI21X1 g13794(.A0 (n_4845), .A1 (n_7709), .B0 (n_4622), .Y (n_5197));
OAI21X1 g13796(.A0 (n_5194), .A1 (n_4525), .B0 (n_5166), .Y (n_5703));
OAI21X1 g13798(.A0 (n_4842), .A1 (n_7170), .B0 (n_4628), .Y (n_5193));
AOI22X1 g13809(.A0 (n_4826), .A1 (n_7714), .B0 (n_4849), .B1(n_4558), .Y (n_5191));
NAND3X1 g13816(.A (n_5188), .B (n_4788), .C (n_4485), .Y (n_5189));
NAND2X1 g13818(.A (n_4681), .B (n_5133), .Y (n_5187));
INVX1 g13843(.A (n_5096), .Y (n_7525));
AOI21X1 g13846(.A0 (n_4824), .A1 (n_5184), .B0 (n_4727), .Y (n_5185));
NAND2X1 g13853(.A (n_5012), .B (n_5931), .Y (n_7587));
NAND2X1 g13862(.A (n_4876), .B (n_5180), .Y (n_5181));
NAND2X1 g13898(.A (n_5056), .B (n_5214), .Y (n_5178));
NAND2X1 g13909(.A (n_5029), .B (n_4443), .Y (n_5176));
NAND2X1 g13910(.A (n_7531), .B (n_7532), .Y (n_5279));
OAI21X1 g13922(.A0 (n_6373), .A1 (n_7322), .B0 (n_4663), .Y (n_5173));
NOR2X1 g13925(.A (n_4511), .B (n_4933), .Y (n_5172));
NAND2X1 g13932(.A (n_4191), .B (n_4791), .Y (n_5171));
NAND2X1 g13956(.A (n_4782), .B (n_4106), .Y (n_5170));
NAND2X1 g13967(.A (n_4783), .B (n_7321), .Y (n_5169));
NAND2X1 g13968(.A (n_4804), .B (n_5062), .Y (n_5168));
NAND2X1 g13969(.A (n_5166), .B (n_4639), .Y (n_5167));
NOR2X1 g13970(.A (n_4813), .B (n_7543), .Y (n_5165));
NOR3X1 g13974(.A (n_4509), .B (n_4784), .C (n_4591), .Y (n_5164));
NAND2X1 g13975(.A (n_4775), .B (n_6094), .Y (n_5163));
NAND2X1 g13976(.A (n_4981), .B (n_4430), .Y (n_5162));
NOR2X1 g13977(.A (n_4747), .B (n_4809), .Y (n_5161));
NAND2X1 g13983(.A (n_4759), .B (n_7360), .Y (n_5160));
INVX1 g14001(.A (n_5157), .Y (n_5158));
NAND2X1 g14006(.A (n_4787), .B (n_7321), .Y (n_5975));
AND2X1 g14012(.A (n_4999), .B (n_4671), .Y (n_5155));
NAND3X1 g14018(.A (n_7463), .B (n_5024), .C (n_4217), .Y (n_5154));
NOR2X1 g14105(.A (n_4780), .B (n_4391), .Y (n_7775));
NAND2X1 g14107(.A (n_4825), .B (n_6207), .Y (n_5151));
INVX1 g14108(.A (n_5013), .Y (n_5150));
NOR2X1 g14142(.A (n_4653), .B (n_4810), .Y (n_5149));
AOI21X1 g14143(.A0 (n_4245), .A1 (n_4226), .B0 (n_4815), .Y (n_7776));
OAI21X1 g13745(.A0 (n_4733), .A1 (n_4425), .B0 (n_4854), .Y (n_5147));
NAND3X1 g13748(.A (n_4442), .B (n_4633), .C (n_4948), .Y (n_5144));
AOI21X1 g13749(.A0 (n_4704), .A1 (n_5948), .B0 (n_4472), .Y (n_7539));
AOI21X1 g13751(.A0 (n_4710), .A1 (n_7237), .B0 (n_4691), .Y (n_5142));
NAND3X1 g13759(.A (n_5140), .B (n_4729), .C (n_4440), .Y (n_5141));
OAI21X1 g13760(.A0 (n_4690), .A1 (n_3968), .B0 (n_5938), .Y (n_5891));
NOR2X1 g13761(.A (n_4724), .B (n_4774), .Y (n_5138));
NAND2X1 g13769(.A (n_4768), .B (n_4976), .Y (n_6869));
OAI21X1 g13770(.A0 (n_4683), .A1 (n_4517), .B0 (n_4908), .Y (n_5136));
INVX1 g14216(.A (n_5133), .Y (n_5134));
NAND3X1 g13779(.A (n_5131), .B (n_6403), .C (n_4988), .Y (n_5132));
OAI21X1 g13780(.A0 (n_4738), .A1 (n_5129), .B0 (n_4554), .Y (n_5696));
OAI21X1 g13786(.A0 (n_4706), .A1 (n_4615), .B0 (n_7463), .Y (n_7884));
AOI21X1 g13792(.A0 (n_4673), .A1 (n_4082), .B0 (n_7321), .Y (n_5126));
NAND2X1 g13793(.A (n_4757), .B (n_6744), .Y (n_5124));
NAND2X1 g13803(.A (n_4770), .B (n_5121), .Y (n_7796));
NOR2X1 g13810(.A (n_4510), .B (n_4772), .Y (n_5119));
NAND2X1 g13812(.A (n_4847), .B (n_5166), .Y (n_5118));
AOI21X1 g13817(.A0 (n_4641), .A1 (n_4727), .B0 (n_5113), .Y (n_5114));
NAND2X1 g13823(.A (n_4837), .B (n_4077), .Y (n_5112));
NAND2X1 g13824(.A (n_5108), .B (n_7417), .Y (n_5111));
NAND2X1 g13827(.A (n_5108), .B (n_5931), .Y (n_7789));
NAND2X1 g13828(.A (n_4836), .B (n_5931), .Y (n_5106));
NAND4X1 g13829(.A (n_5104), .B (n_6103), .C (n_4519), .D (n_4521), .Y(n_5105));
NOR2X1 g13830(.A (n_4701), .B (n_7466), .Y (n_5103));
NOR2X1 g13831(.A (n_4853), .B (n_4926), .Y (n_5102));
NOR2X1 g13834(.A (n_7171), .B (n_5681), .Y (n_5311));
NAND2X1 g13837(.A (n_5100), .B (n_5099), .Y (n_5101));
NOR2X1 g13841(.A (n_5194), .B (n_5018), .Y (n_5097));
NAND2X1 g13844(.A (n_4920), .B (n_4765), .Y (n_5096));
NAND2X1 g13845(.A (n_4730), .B (n_6829), .Y (n_5095));
INVX1 g13851(.A (n_4969), .Y (n_7778));
NAND2X1 g13858(.A (n_4834), .B (n_4705), .Y (n_5084));
NAND3X1 g13859(.A (n_4829), .B (n_4604), .C (n_4582), .Y (n_5083));
AOI21X1 g13861(.A0 (n_4638), .A1 (n_4952), .B0 (n_5010), .Y (n_5082));
NAND2X1 g13866(.A (n_4894), .B (n_4763), .Y (n_5081));
NOR2X1 g13870(.A (n_5008), .B (n_4755), .Y (n_6088));
NAND2X1 g13877(.A (n_4696), .B (n_5001), .Y (n_5077));
NAND2X1 g13879(.A (n_4865), .B (n_5365), .Y (n_5075));
NAND2X1 g13880(.A (n_4921), .B (n_7321), .Y (n_6104));
OAI21X1 g13890(.A0 (n_4642), .A1 (n_4257), .B0 (n_5010), .Y (n_5072));
AOI21X1 g13895(.A0 (n_4598), .A1 (n_5010), .B0 (n_4499), .Y (n_5070));
INVX1 g13919(.A (n_4936), .Y (n_5068));
OAI21X1 g13921(.A0 (n_4431), .A1 (n_3994), .B0 (n_4409), .Y (n_5067));
NOR2X1 g13926(.A (n_4286), .B (n_7171), .Y (n_5065));
NAND2X1 g13929(.A (n_4610), .B (n_5059), .Y (n_5974));
NAND2X1 g13930(.A (n_4602), .B (n_5059), .Y (n_5060));
NAND2X1 g13941(.A (n_4533), .B (n_4478), .Y (n_5058));
NOR2X1 g13942(.A (n_4752), .B (n_4803), .Y (n_7522));
NAND2X1 g13943(.A (n_4603), .B (n_4934), .Y (n_5056));
OR2X1 g13949(.A (n_4666), .B (n_6048), .Y (n_5055));
NAND2X1 g13951(.A (n_4478), .B (n_4739), .Y (n_5054));
NAND2X1 g13957(.A (n_4605), .B (n_5015), .Y (n_5053));
NAND2X1 g13958(.A (n_4606), .B (n_4551), .Y (n_5052));
NAND2X1 g13959(.A (n_4592), .B (n_4460), .Y (n_5051));
NAND3X1 g13962(.A (n_4380), .B (n_4908), .C (n_4428), .Y (n_5687));
NAND2X1 g13972(.A (n_4609), .B (n_4955), .Y (n_5049));
NOR2X1 g13978(.A (n_4679), .B (n_4651), .Y (n_5048));
NAND2X1 g13982(.A (n_4561), .B (n_4652), .Y (n_7599));
AND2X1 g13985(.A (n_5044), .B (n_4777), .Y (n_5045));
NAND3X1 g13989(.A (n_5042), .B (n_4250), .C (n_5041), .Y (n_5601));
NOR3X1 g13999(.A (n_7142), .B (n_4423), .C (n_4861), .Y (n_5040));
NOR3X1 g14000(.A (n_4599), .B (n_7709), .C (n_4133), .Y (n_5039));
NOR2X1 g14002(.A (n_5038), .B (n_5121), .Y (n_5157));
NAND2X1 g14005(.A (n_5188), .B (n_6451), .Y (n_5037));
NAND2X1 g14011(.A (n_4983), .B (n_4846), .Y (n_5036));
AND2X1 g14013(.A (n_5034), .B (n_4478), .Y (n_5035));
NOR2X1 g14014(.A (n_4648), .B (n_4942), .Y (n_5032));
NAND4X1 g14019(.A (n_4923), .B (n_4665), .C (n_6048), .D (n_4161), .Y(n_5180));
INVX1 g14023(.A (n_4904), .Y (n_5030));
NAND2X1 g14025(.A (n_5004), .B (n_4832), .Y (n_5029));
NAND2X1 g14026(.A (n_4600), .B (n_7714), .Y (n_5028));
NOR3X1 g14048(.A (n_7251), .B (n_4902), .C (n_4795), .Y (n_5026));
NAND2X1 g14049(.A (n_5024), .B (n_4856), .Y (n_5025));
INVX1 g14057(.A (n_4884), .Y (n_5892));
NAND2X1 g14061(.A (n_4597), .B (n_7714), .Y (n_5597));
NAND2X1 g14076(.A (n_4293), .B (n_4616), .Y (n_5020));
INVX1 g14079(.A (n_5018), .Y (n_5019));
NAND2X1 g14082(.A (n_4808), .B (n_5203), .Y (n_5017));
NOR2X1 g14084(.A (n_5015), .B (n_4694), .Y (n_5016));
NOR2X1 g14104(.A (n_4646), .B (n_4527), .Y (n_5014));
OAI21X1 g14109(.A0 (n_4414), .A1 (n_3844), .B0 (n_4412), .Y (n_5013));
NAND2X1 g14113(.A (n_4612), .B (n_4871), .Y (n_5012));
INVX1 g14116(.A (n_5008), .Y (n_6872));
NAND2X1 g14134(.A (n_5004), .B (n_7542), .Y (n_5005));
NAND2X1 g14153(.A (n_4430), .B (n_4996), .Y (n_5003));
NAND3X1 g13754(.A (n_5001), .B (n_4508), .C (n_4543), .Y (n_5002));
INVX1 g14198(.A (n_4999), .Y (n_5000));
NAND2X1 g14217(.A (n_4996), .B (n_3994), .Y (n_5133));
NAND2X1 g14225(.A (n_4647), .B (n_4996), .Y (n_4995));
NAND2X1 g14237(.A (n_4238), .B (n_7228), .Y (n_4994));
AOI22X1 g13797(.A0 (n_4536), .A1 (n_4554), .B0 (n_4279), .B1(n_4572), .Y (n_7795));
AOI21X1 g13800(.A0 (n_4832), .A1 (n_4988), .B0 (n_7465), .Y (n_4989));
NAND3X1 g13805(.A (n_4745), .B (n_5099), .C (n_4773), .Y (n_4986));
INVX1 g14368(.A (n_4981), .Y (n_4982));
AOI21X1 g13821(.A0 (n_4491), .A1 (n_7228), .B0 (n_6676), .Y (n_4980));
NAND3X1 g13832(.A (n_4875), .B (n_4976), .C (n_4309), .Y (n_4977));
NAND2X1 g13835(.A (n_7171), .B (n_4893), .Y (n_4975));
NOR2X1 g13836(.A (n_4744), .B (n_4973), .Y (n_5697));
NAND2X1 g13852(.A (n_6403), .B (n_7467), .Y (n_4969));
NAND3X1 g13855(.A (n_4675), .B (n_4438), .C (n_4124), .Y (n_4967));
NAND2X1 g13857(.A (n_4753), .B (n_4769), .Y (n_4966));
NOR2X1 g13863(.A (n_4841), .B (n_4880), .Y (n_4965));
NAND2X1 g13865(.A (n_4963), .B (n_4551), .Y (n_4964));
NOR2X1 g13867(.A (n_4702), .B (n_4877), .Y (n_7530));
NAND2X1 g13868(.A (n_6403), .B (n_4758), .Y (n_4960));
NOR2X1 g13869(.A (n_4708), .B (n_4626), .Y (n_4959));
NAND3X1 g13876(.A (n_4902), .B (n_7237), .C (n_4447), .Y (n_4957));
OAI21X1 g13881(.A0 (n_4436), .A1 (n_4273), .B0 (n_4955), .Y (n_4956));
NAND3X1 g13884(.A (n_5015), .B (n_4164), .C (n_4447), .Y (n_4954));
INVX1 g13888(.A (n_4950), .Y (n_7885));
NAND2X1 g13892(.A (n_4684), .B (n_4948), .Y (n_4949));
AOI21X1 g13894(.A0 (n_4737), .A1 (n_4657), .B0 (n_4554), .Y (n_4947));
NAND2X1 g13900(.A (n_4720), .B (n_4721), .Y (n_4944));
AOI21X1 g13903(.A0 (n_4432), .A1 (n_7714), .B0 (n_4942), .Y (n_4943));
NAND2X1 g13904(.A (n_4662), .B (n_4717), .Y (n_4941));
AOI21X1 g13906(.A0 (n_4433), .A1 (n_7426), .B0 (n_4801), .Y (n_4940));
INVX1 g13907(.A (n_4938), .Y (n_4939));
NAND2X1 g13912(.A (n_4546), .B (n_4700), .Y (n_4937));
AOI21X1 g13920(.A0 (n_4471), .A1 (n_4198), .B0 (n_7426), .Y (n_4936));
OAI21X1 g13923(.A0 (n_4632), .A1 (n_4934), .B0 (n_4468), .Y (n_4935));
AOI21X1 g13927(.A0 (n_4263), .A1 (n_4732), .B0 (n_4854), .Y (n_4933));
NAND2X1 g13936(.A (n_4931), .B (n_4736), .Y (n_4932));
NOR2X1 g13937(.A (n_4380), .B (n_4907), .Y (n_4930));
NOR2X1 g13944(.A (n_4613), .B (n_4864), .Y (n_4928));
INVX1 g13945(.A (n_4926), .Y (n_4927));
NOR2X1 g13947(.A (n_4601), .B (n_4245), .Y (n_4925));
NAND3X1 g13950(.A (n_4923), .B (n_7171), .C (n_4873), .Y (n_4924));
NOR2X1 g13955(.A (n_4819), .B (n_4525), .Y (n_6012));
NAND3X1 g13963(.A (n_7774), .B (n_4106), .C (n_4222), .Y (n_4921));
NAND3X1 g13971(.A (n_4126), .B (n_4542), .C (n_4661), .Y (n_4920));
NAND2X1 g13979(.A (n_5044), .B (n_4040), .Y (n_4919));
OAI21X1 g13987(.A0 (n_4280), .A1 (n_4281), .B0 (n_3994), .Y (n_4918));
NAND3X1 g13998(.A (n_4542), .B (n_6823), .C (n_4719), .Y (n_5100));
NOR2X1 g14004(.A (n_4486), .B (n_4399), .Y (n_4912));
NOR2X1 g14009(.A (n_4908), .B (n_4907), .Y (n_4909));
NAND2X1 g14024(.A (n_4885), .B (n_4835), .Y (n_4904));
NAND4X1 g14027(.A (n_4902), .B (n_7251), .C (n_3938), .D (n_4068), .Y(n_4903));
NAND3X1 g14029(.A (n_4449), .B (n_5948), .C (n_7413), .Y (n_4900));
NAND2X1 g14030(.A (n_5938), .B (n_4462), .Y (n_7540));
NAND2X1 g14032(.A (n_4902), .B (n_4711), .Y (n_4896));
NAND2X1 g14034(.A (n_7362), .B (n_4474), .Y (n_7532));
INVX1 g14038(.A (n_4893), .Y (n_4894));
NAND2X1 g14041(.A (n_4839), .B (n_4870), .Y (n_4892));
NAND2X1 g14042(.A (n_7426), .B (n_4458), .Y (n_4891));
NAND3X1 g14043(.A (n_5931), .B (n_4366), .C (n_4302), .Y (n_4889));
NAND2X1 g14047(.A (n_4627), .B (n_4863), .Y (n_4888));
NAND2X1 g14055(.A (n_7362), .B (n_4617), .Y (n_7531));
NAND2X1 g14056(.A (n_4631), .B (n_4885), .Y (n_4886));
NAND2X1 g14058(.A (n_4623), .B (n_4883), .Y (n_4884));
INVX1 g14059(.A (n_4699), .Y (n_7588));
INVX2 g14064(.A (n_4880), .Y (n_5681));
NAND3X1 g14071(.A (n_4875), .B (n_7170), .C (n_4873), .Y (n_4876));
NAND2X1 g14072(.A (n_4871), .B (n_4870), .Y (n_4872));
NAND2X1 g14073(.A (n_5948), .B (n_4455), .Y (n_4869));
AOI21X1 g14074(.A0 (n_4424), .A1 (n_4332), .B0 (n_4345), .Y (n_4868));
NAND2X1 g14075(.A (n_4660), .B (n_4866), .Y (n_4867));
NOR2X1 g14077(.A (n_4864), .B (n_4863), .Y (n_4865));
NOR3X1 g14080(.A (n_3851), .B (n_4854), .C (n_4608), .Y (n_5018));
NOR3X1 g14083(.A (n_4908), .B (n_3899), .C (n_4861), .Y (n_4862));
NAND3X1 g14092(.A (n_4621), .B (n_4596), .C (n_4650), .Y (n_4859));
NAND2X1 g14097(.A (n_7362), .B (n_4856), .Y (n_4858));
NAND2X1 g14100(.A (n_4534), .B (n_4854), .Y (n_5590));
NOR3X1 g14101(.A (n_7900), .B (n_4743), .C (n_4159), .Y (n_4853));
NAND3X1 g14103(.A (n_4660), .B (n_7322), .C (n_4226), .Y (n_6105));
NAND2X1 g14112(.A (n_4531), .B (n_4849), .Y (n_4850));
NOR2X1 g14117(.A (n_4569), .B (n_7360), .Y (n_5008));
OAI21X1 g14120(.A0 (n_4813), .A1 (n_3983), .B0 (n_4846), .Y (n_4847));
NAND2X1 g14121(.A (n_4494), .B (n_4599), .Y (n_4845));
NAND2X1 g14123(.A (n_4419), .B (n_6451), .Y (n_4844));
NAND2X1 g14124(.A (n_4513), .B (n_6062), .Y (n_4843));
NOR2X1 g14127(.A (n_4841), .B (n_6100), .Y (n_4842));
NAND2X1 g14128(.A (n_4470), .B (n_4839), .Y (n_4840));
NAND2X1 g14129(.A (n_4079), .B (n_4838), .Y (n_5108));
AOI21X1 g14130(.A0 (n_4476), .A1 (n_7413), .B0 (n_4469), .Y (n_4837));
NAND2X1 g14131(.A (n_3972), .B (n_4835), .Y (n_4836));
NAND2X1 g14135(.A (n_4464), .B (n_4537), .Y (n_4834));
NAND2X1 g14136(.A (n_4394), .B (n_4832), .Y (n_4833));
NAND2X2 g14137(.A (n_4496), .B (n_5034), .Y (n_5194));
NAND2X1 g14138(.A (n_4453), .B (n_4709), .Y (n_4831));
NAND2X1 g14139(.A (n_4497), .B (n_4088), .Y (n_4830));
AOI21X1 g14140(.A0 (n_7358), .A1 (n_4828), .B0 (n_4388), .Y (n_4829));
NAND2X1 g14144(.A (n_4532), .B (n_4203), .Y (n_4827));
NAND2X1 g14145(.A (n_4058), .B (n_4493), .Y (n_4826));
NAND2X1 g14152(.A (n_4145), .B (n_4247), .Y (n_4825));
NAND2X1 g14154(.A (n_4823), .B (n_4410), .Y (n_4824));
NAND2X1 g14158(.A (n_4271), .B (n_4854), .Y (n_7543));
NAND2X1 g14163(.A (n_5129), .B (n_4554), .Y (n_4821));
INVX1 g14165(.A (n_4983), .Y (n_4819));
NAND2X1 g14183(.A (n_4337), .B (n_4812), .Y (n_4818));
INVX1 g14186(.A (n_7317), .Y (n_4817));
NOR2X1 g14197(.A (n_4814), .B (n_4421), .Y (n_4815));
NAND2X1 g14199(.A (n_4813), .B (n_4812), .Y (n_4999));
NAND2X1 g14208(.A (n_7735), .B (n_4593), .Y (n_4810));
INVX1 g14233(.A (n_4808), .Y (n_4809));
NAND3X1 g14242(.A (n_4637), .B (n_4570), .C (n_4046), .Y (n_4807));
INVX1 g14269(.A (n_4803), .Y (n_4804));
NAND2X1 g14295(.A (n_4619), .B (n_4797), .Y (n_4800));
NAND2X1 g14323(.A (n_4180), .B (n_4797), .Y (n_4799));
OR2X1 g14335(.A (n_7362), .B (n_4795), .Y (n_4796));
AND2X1 g13819(.A (n_7111), .B (n_6677), .Y (n_5598));
AOI21X1 g14369(.A0 (n_4177), .A1 (n_4381), .B0 (n_4405), .Y (n_4981));
NAND2X1 g14374(.A (n_4178), .B (n_4589), .Y (n_4791));
NAND2X1 g14378(.A (n_4426), .B (n_7320), .Y (n_4788));
NAND2X1 g14381(.A (n_4386), .B (n_4514), .Y (n_4787));
NAND3X1 g13825(.A (n_6786), .B (n_4333), .C (n_4784), .Y (n_5704));
NAND2X1 g14384(.A (n_4418), .B (n_4082), .Y (n_4783));
AOI21X1 g14389(.A0 (n_4635), .A1 (n_4781), .B0 (n_4049), .Y (n_4782));
NAND2X1 g14394(.A (n_4264), .B (n_6532), .Y (n_4780));
NAND2X1 g14399(.A (n_4096), .B (n_4406), .Y (n_4779));
INVX1 g14400(.A (n_4777), .Y (n_4778));
INVX1 g14405(.A (n_4996), .Y (n_4775));
NAND2X1 g13840(.A (n_5099), .B (n_4773), .Y (n_4774));
AOI21X1 g13842(.A0 (n_4338), .A1 (n_4260), .B0 (n_4784), .Y (n_4772));
NAND2X1 g13854(.A (n_4769), .B (n_6740), .Y (n_4770));
NAND2X1 g13860(.A (n_4767), .B (n_4934), .Y (n_4768));
NAND2X1 g13864(.A (n_4349), .B (n_4765), .Y (n_4766));
NAND2X1 g13873(.A (n_4696), .B (n_4763), .Y (n_4764));
NAND2X1 g13875(.A (n_4692), .B (n_4694), .Y (n_4762));
INVX1 g14537(.A (n_4760), .Y (n_4761));
NAND2X1 g14550(.A (n_4573), .B (n_4068), .Y (n_4759));
NAND2X1 g13889(.A (n_4685), .B (n_4758), .Y (n_4950));
NAND2X1 g13902(.A (n_4368), .B (n_4907), .Y (n_4757));
OAI21X1 g13905(.A0 (n_4457), .A1 (n_4212), .B0 (n_4754), .Y (n_4756));
INVX1 g14623(.A (n_5004), .Y (n_4755));
OAI21X1 g13908(.A0 (n_4449), .A1 (n_4669), .B0 (n_4754), .Y (n_4938));
NAND3X1 g14634(.A (n_4323), .B (n_4125), .C (n_6830), .Y (n_4753));
INVX1 g14635(.A (n_6993), .Y (n_4752));
OAI21X1 g13915(.A0 (n_7360), .A1 (n_4539), .B0 (n_4296), .Y (n_4750));
OR2X1 g14690(.A (n_7488), .B (n_5203), .Y (n_4747));
NAND2X1 g13931(.A (n_4561), .B (n_4339), .Y (n_4745));
INVX1 g13934(.A (n_4769), .Y (n_4744));
NOR2X1 g13946(.A (n_4743), .B (n_4307), .Y (n_4926));
INVX1 g13952(.A (n_4740), .Y (n_4741));
NAND2X1 g13960(.A (n_4737), .B (n_4736), .Y (n_4738));
INVX1 g13964(.A (n_4773), .Y (n_4734));
NAND2X1 g13966(.A (n_4478), .B (n_4732), .Y (n_4733));
NAND2X1 g13973(.A (n_6744), .B (n_4562), .Y (n_7526));
INVX1 g13980(.A (n_4973), .Y (n_4730));
NAND4X1 g13986(.A (n_4728), .B (n_4727), .C (n_3844), .D (n_4045), .Y(n_5140));
NAND4X1 g13988(.A (n_4728), .B (n_4727), .C (n_6007), .D (n_4405), .Y(n_4729));
NAND2X1 g13993(.A (n_4380), .B (n_4487), .Y (n_4726));
INVX1 g13996(.A (n_4723), .Y (n_4724));
NAND3X1 g14010(.A (n_6822), .B (n_4554), .C (n_3982), .Y (n_4721));
NAND3X1 g14015(.A (n_4561), .B (n_4554), .C (n_4719), .Y (n_4720));
INVX1 g14016(.A (n_4717), .Y (n_4718));
NAND2X1 g14028(.A (n_4711), .B (n_7362), .Y (n_5131));
NAND2X1 g14031(.A (n_4709), .B (n_4473), .Y (n_4710));
NOR3X1 g14033(.A (n_3896), .B (n_7800), .C (n_5935), .Y (n_4708));
NAND2X1 g14035(.A (n_4446), .B (n_4832), .Y (n_4706));
NAND2X1 g14037(.A (n_4301), .B (n_4467), .Y (n_4963));
NAND2X1 g14039(.A (n_6009), .B (n_4705), .Y (n_4893));
NAND2X1 g14040(.A (n_4392), .B (n_4698), .Y (n_4704));
NOR2X1 g14044(.A (n_4459), .B (n_4158), .Y (n_4703));
NOR2X1 g14046(.A (n_4158), .B (n_4763), .Y (n_4702));
INVX1 g14052(.A (n_4700), .Y (n_4701));
NAND2X1 g14060(.A (n_4698), .B (n_4885), .Y (n_4699));
NAND2X1 g14062(.A (n_7237), .B (n_4310), .Y (n_4697));
NOR2X1 g14065(.A (n_4545), .B (n_4307), .Y (n_4880));
INVX1 g14067(.A (n_4696), .Y (n_4877));
NAND2X1 g14085(.A (n_4293), .B (n_4694), .Y (n_4695));
INVX1 g14087(.A (n_4692), .Y (n_4691));
NAND2X1 g14090(.A (n_4389), .B (n_4714), .Y (n_4690));
NAND3X1 g14091(.A (n_7712), .B (n_4037), .C (n_4676), .Y (n_4689));
NAND2X1 g14093(.A (n_4284), .B (n_4327), .Y (n_4687));
INVX1 g14094(.A (n_4685), .Y (n_4686));
NOR2X1 g14098(.A (n_4548), .B (n_4441), .Y (n_4684));
OAI21X1 g14102(.A0 (n_6823), .A1 (n_3978), .B0 (n_4427), .Y (n_4683));
NAND2X1 g14106(.A (n_4335), .B (n_4739), .Y (n_4682));
AOI21X1 g14110(.A0 (n_7488), .A1 (n_4528), .B0 (n_4679), .Y (n_4681));
NAND3X1 g14111(.A (n_4677), .B (n_4252), .C (n_4676), .Y (n_4678));
NAND2X1 g14118(.A (n_4329), .B (n_6823), .Y (n_4675));
AOI21X1 g14122(.A0 (n_6441), .A1 (n_4223), .B0 (n_4420), .Y (n_4673));
NAND2X1 g14126(.A (n_4244), .B (n_4671), .Y (n_4672));
NAND2X1 g14133(.A (n_4313), .B (n_4669), .Y (n_4670));
NAND2X1 g14148(.A (n_3870), .B (n_4644), .Y (n_4668));
NAND2X1 g14161(.A (n_6823), .B (n_4213), .Y (n_4667));
NAND2X1 g14164(.A (n_4665), .B (n_4275), .Y (n_4666));
NAND2X1 g14181(.A (n_3988), .B (n_4226), .Y (n_4663));
NAND2X1 g14185(.A (n_4719), .B (n_4661), .Y (n_4662));
INVX1 g14194(.A (n_4657), .Y (n_4658));
NAND2X1 g14196(.A (n_7323), .B (n_4634), .Y (n_4656));
NAND2X1 g14200(.A (n_4813), .B (n_4277), .Y (n_4655));
NAND2X1 g14209(.A (n_4249), .B (n_5092), .Y (n_4653));
NOR2X1 g14213(.A (n_4323), .B (n_3978), .Y (n_4652));
INVX1 g14214(.A (n_5184), .Y (n_4651));
NOR2X1 g14218(.A (n_7227), .B (n_4650), .Y (n_4942));
INVX1 g14219(.A (n_4648), .Y (n_4649));
NOR2X1 g14224(.A (n_4647), .B (n_5092), .Y (n_5113));
NOR3X1 g14226(.A (n_4495), .B (n_4526), .C (n_4195), .Y (n_4646));
NAND2X1 g14234(.A (n_4098), .B (n_4645), .Y (n_4808));
NAND2X1 g14243(.A (n_4644), .B (n_4322), .Y (n_5038));
NAND2X1 g14248(.A (n_4088), .B (n_6478), .Y (n_4642));
NAND2X1 g14255(.A (n_4249), .B (n_7735), .Y (n_4641));
NAND2X1 g14267(.A (n_4637), .B (n_4095), .Y (n_4638));
NOR2X1 g14270(.A (n_6441), .B (n_4398), .Y (n_4803));
NAND2X1 g14273(.A (n_4632), .B (n_4873), .Y (n_4633));
INVX1 g14277(.A (n_4631), .Y (n_4801));
NOR2X1 g14287(.A (n_7228), .B (n_4219), .Y (n_4630));
NAND3X1 g14293(.A (n_6047), .B (n_4627), .C (n_4665), .Y (n_4628));
INVX1 g14296(.A (n_4835), .Y (n_4626));
NAND2X1 g14299(.A (n_4551), .B (n_4873), .Y (n_4625));
INVX1 g14302(.A (n_4623), .Y (n_4624));
INVX1 g14305(.A (n_4621), .Y (n_4622));
NOR2X1 g14329(.A (n_4619), .B (n_4198), .Y (n_4620));
INVX1 g14351(.A (n_4615), .Y (n_4616));
NAND3X1 g14367(.A (n_3897), .B (n_4366), .C (n_4180), .Y (n_4612));
NAND2X1 g14380(.A (n_6478), .B (n_4239), .Y (n_5089));
NAND2X1 g14382(.A (n_4220), .B (n_4390), .Y (n_4610));
NAND2X1 g14383(.A (n_4268), .B (n_4608), .Y (n_4609));
NAND2X1 g14386(.A (n_4216), .B (n_4118), .Y (n_4606));
NAND2X1 g14390(.A (n_4206), .B (n_4604), .Y (n_4605));
NOR2X1 g14391(.A (n_4215), .B (n_4065), .Y (n_4603));
INVX1 g14392(.A (n_4601), .Y (n_4602));
NAND2X1 g14395(.A (n_4253), .B (n_4599), .Y (n_4600));
NAND2X1 g14397(.A (n_4242), .B (n_4490), .Y (n_4598));
NAND2X1 g14398(.A (n_4231), .B (n_4596), .Y (n_4597));
NAND3X1 g14401(.A (n_4054), .B (n_4727), .C (n_4403), .Y (n_4777));
NAND4X1 g13833(.A (n_4976), .B (n_4875), .C (n_3965), .D (n_4665), .Y(n_5220));
NOR2X1 g14403(.A (n_4594), .B (n_4576), .Y (n_4595));
INVX2 g14406(.A (n_4593), .Y (n_4996));
NOR2X1 g14412(.A (n_4551), .B (n_7170), .Y (n_4592));
INVX1 g14437(.A (n_4812), .Y (n_4591));
INVX1 g14462(.A (n_4589), .Y (n_4590));
NOR2X1 g14509(.A (n_7228), .B (n_4094), .Y (n_4585));
NOR2X1 g14538(.A (n_4027), .B (n_4289), .Y (n_4760));
NAND2X2 g14543(.A (n_6888), .B (n_6095), .Y (n_5188));
INVX1 g14561(.A (n_4395), .Y (n_5024));
NOR3X1 g13887(.A (n_4582), .B (n_7464), .C (n_6402), .Y (n_4584));
NAND2X1 g14622(.A (n_4580), .B (n_4540), .Y (n_4581));
NAND2X2 g14624(.A (n_4580), .B (n_4068), .Y (n_5004));
NOR2X1 g14628(.A (n_4365), .B (n_4059), .Y (n_4579));
AND2X1 g14660(.A (n_7712), .B (n_7121), .Y (n_4578));
INVX1 g14695(.A (n_4576), .Y (n_4577));
INVX1 g14699(.A (n_4574), .Y (n_4575));
NOR2X1 g14706(.A (n_7359), .B (n_7760), .Y (n_4573));
NAND4X1 g13935(.A (n_4278), .B (n_4482), .C (n_4572), .D (n_3870), .Y(n_4769));
NAND2X1 g14735(.A (n_7359), .B (n_7462), .Y (n_4569));
NAND3X1 g13948(.A (n_4025), .B (n_4214), .C (n_3965), .Y (n_5224));
NAND4X1 g13953(.A (n_4813), .B (n_4955), .C (n_4050), .D (n_3984), .Y(n_4740));
NAND2X1 g13965(.A (n_4480), .B (n_4562), .Y (n_4773));
NOR2X1 g13981(.A (n_4736), .B (n_4561), .Y (n_4973));
NAND2X1 g13997(.A (n_4541), .B (n_6746), .Y (n_4723));
NAND2X1 g14017(.A (n_4554), .B (n_6942), .Y (n_4717));
INVX2 g15104(.A (n_7362), .Y (n_4902));
INVX1 g15116(.A (n_6402), .Y (n_5015));
INVX2 g15194(.A (n_7228), .Y (n_5010));
NAND2X1 g14036(.A (n_4551), .B (n_4306), .Y (n_4767));
NAND2X1 g14045(.A (n_4544), .B (n_4548), .Y (n_4549));
NAND2X1 g14050(.A (n_7359), .B (n_7741), .Y (n_4988));
NAND2X1 g14051(.A (n_4443), .B (n_7741), .Y (n_4546));
NAND2X1 g14053(.A (n_7463), .B (n_4294), .Y (n_4700));
NAND4X1 g14068(.A (n_4013), .B (n_6047), .C (n_4012), .D (n_4285), .Y(n_4696));
NAND2X1 g14069(.A (n_4545), .B (n_4309), .Y (n_5001));
NAND2X1 g14070(.A (n_4300), .B (n_4544), .Y (n_5365));
NAND2X1 g14078(.A (n_4545), .B (n_4548), .Y (n_4543));
NAND3X1 g14081(.A (n_4542), .B (n_4541), .C (n_4719), .Y (n_4765));
NAND4X1 g14088(.A (n_7359), .B (n_7248), .C (n_4540), .D (n_6817), .Y(n_4692));
NAND2X1 g14095(.A (n_4539), .B (n_6707), .Y (n_4685));
NAND2X1 g14096(.A (n_4539), .B (n_7741), .Y (n_4758));
NAND2X1 g14099(.A (n_4537), .B (n_4308), .Y (n_4948));
OAI21X1 g14115(.A0 (n_4480), .A1 (n_7706), .B0 (n_4516), .Y (n_4536));
NAND2X1 g14150(.A (n_4533), .B (n_4435), .Y (n_4534));
NAND2X1 g14155(.A (n_4430), .B (n_4255), .Y (n_4532));
NAND2X1 g14159(.A (n_4501), .B (n_4728), .Y (n_5042));
NOR2X1 g14160(.A (n_7121), .B (n_4488), .Y (n_4531));
NAND2X1 g14162(.A (n_7492), .B (n_4528), .Y (n_4529));
NOR2X1 g14170(.A (n_4526), .B (n_4108), .Y (n_4527));
INVX1 g14172(.A (n_4524), .Y (n_4525));
INVX1 g14175(.A (n_4521), .Y (n_4522));
NAND2X1 g14179(.A (n_4345), .B (n_4107), .Y (n_6103));
NAND2X1 g14180(.A (n_4337), .B (n_4261), .Y (n_4519));
NOR2X1 g14182(.A (n_4285), .B (n_4274), .Y (n_4518));
NOR2X1 g14184(.A (n_4516), .B (n_4541), .Y (n_4517));
NAND2X1 g14189(.A (n_4514), .B (n_4269), .Y (n_4515));
NAND2X1 g14190(.A (n_3988), .B (n_4105), .Y (n_4513));
NOR2X1 g14191(.A (n_4813), .B (n_4276), .Y (n_4511));
NAND2X1 g14195(.A (n_4541), .B (n_4204), .Y (n_4657));
NOR2X1 g14201(.A (n_4509), .B (n_4272), .Y (n_4510));
NAND2X1 g14204(.A (n_4743), .B (n_4065), .Y (n_4508));
NAND2X1 g14215(.A (n_4647), .B (n_7479), .Y (n_5184));
NOR2X1 g14220(.A (n_4504), .B (n_4256), .Y (n_4648));
NAND3X1 g14221(.A (n_3919), .B (n_7492), .C (n_4439), .Y (n_5044));
NAND2X1 g14222(.A (n_3994), .B (n_4247), .Y (n_4503));
NAND2X1 g14223(.A (n_4501), .B (n_7492), .Y (n_5895));
NOR2X1 g14229(.A (n_4498), .B (n_4599), .Y (n_4499));
NAND2X1 g14230(.A (n_7228), .B (n_4326), .Y (n_4497));
NAND4X1 g14231(.A (n_4495), .B (n_3984), .C (n_4344), .D (n_4340), .Y(n_4496));
NAND4X1 g14232(.A (n_4677), .B (n_3945), .C (n_6476), .D (n_6464), .Y(n_4952));
NAND2X1 g14235(.A (n_4378), .B (n_4492), .Y (n_4494));
NAND2X1 g14236(.A (n_4677), .B (n_4492), .Y (n_4493));
NAND2X1 g14238(.A (n_4091), .B (n_4490), .Y (n_4491));
NAND2X1 g14239(.A (n_4188), .B (n_4488), .Y (n_4489));
INVX1 g14240(.A (n_4487), .Y (n_4907));
NAND2X1 g14249(.A (n_4514), .B (n_4227), .Y (n_4866));
INVX1 g14251(.A (n_4485), .Y (n_4486));
NAND3X1 g14257(.A (n_4126), .B (n_4482), .C (n_3924), .Y (n_4931));
NOR2X1 g14258(.A (n_4480), .B (n_4479), .Y (n_4481));
INVX1 g14263(.A (n_4478), .Y (n_4639));
NAND2X1 g14265(.A (n_4495), .B (n_4271), .Y (n_4846));
NAND2X1 g14272(.A (n_3962), .B (n_4477), .Y (n_4838));
NAND4X1 g14278(.A (n_4476), .B (n_4212), .C (n_7612), .D (n_4312), .Y(n_4631));
INVX1 g14282(.A (n_4473), .Y (n_4474));
INVX1 g14285(.A (n_4471), .Y (n_4472));
NAND2X1 g14288(.A (n_4619), .B (n_4469), .Y (n_4470));
NAND2X1 g14289(.A (n_7890), .B (n_4319), .Y (n_4468));
INVX1 g14290(.A (n_4467), .Y (n_4863));
NAND2X1 g14292(.A (n_4875), .B (n_4320), .Y (n_4466));
NAND4X1 g14297(.A (n_4476), .B (n_4212), .C (n_7605), .D (n_3787), .Y(n_4835));
NAND2X1 g14301(.A (n_4539), .B (n_4317), .Y (n_7542));
NAND2X1 g14303(.A (n_4456), .B (n_4197), .Y (n_4623));
NAND2X1 g14306(.A (n_6674), .B (n_4676), .Y (n_4621));
NAND2X1 g14309(.A (n_3887), .B (n_4119), .Y (n_4464));
INVX1 g14313(.A (n_4885), .Y (n_4462));
INVX1 g14321(.A (n_4459), .Y (n_4460));
INVX1 g14324(.A (n_4457), .Y (n_4458));
NAND2X1 g14330(.A (n_4456), .B (n_4074), .Y (n_4871));
NAND2X1 g14331(.A (n_3834), .B (n_4451), .Y (n_4870));
INVX1 g14332(.A (n_4714), .Y (n_4455));
INVX1 g14338(.A (n_4694), .Y (n_4617));
NAND2X1 g14340(.A (n_6472), .B (n_4676), .Y (n_4454));
NAND2X1 g14342(.A (n_4539), .B (n_7239), .Y (n_4453));
NAND2X1 g14344(.A (n_7417), .B (n_4451), .Y (n_4452));
NAND3X1 g14345(.A (n_4449), .B (n_5938), .C (n_3941), .Y (n_4450));
INVX1 g14347(.A (n_4446), .Y (n_4447));
NOR2X1 g14352(.A (n_4539), .B (n_7253), .Y (n_4615));
NOR2X1 g14356(.A (n_4443), .B (n_4057), .Y (n_4856));
INVX1 g14360(.A (n_4441), .Y (n_4442));
INVX1 g14363(.A (n_4286), .Y (n_4613));
NAND3X1 g14366(.A (n_7491), .B (n_4727), .C (n_4439), .Y (n_4440));
NAND3X1 g14372(.A (n_3870), .B (n_4323), .C (n_4380), .Y (n_4438));
NAND2X1 g14379(.A (n_4062), .B (n_4435), .Y (n_4436));
NOR2X1 g14387(.A (n_4114), .B (n_4218), .Y (n_4434));
NAND2X1 g14388(.A (n_7753), .B (n_7754), .Y (n_4433));
NOR2X1 g14393(.A (n_3873), .B (n_4105), .Y (n_4601));
NAND2X1 g14396(.A (n_4029), .B (n_4596), .Y (n_4432));
AOI21X1 g14402(.A0 (n_4430), .A1 (n_4439), .B0 (n_4189), .Y (n_4431));
NAND2X2 g14407(.A (n_3855), .B (n_4176), .Y (n_4593));
AND2X1 g14410(.A (n_7171), .B (n_5428), .Y (n_4429));
INVX1 g14413(.A (n_4427), .Y (n_4428));
NAND2X1 g14423(.A (n_4375), .B (n_4193), .Y (n_4426));
INVX1 g14424(.A (n_4424), .Y (n_4425));
INVX1 g14426(.A (n_4661), .Y (n_4423));
NOR2X1 g14438(.A (n_4036), .B (n_4047), .Y (n_4812));
INVX1 g14445(.A (n_4420), .Y (n_4421));
NAND2X1 g14447(.A (n_4594), .B (n_4400), .Y (n_4419));
NAND2X1 g14457(.A (n_3988), .B (n_6891), .Y (n_4418));
NAND2X1 g14463(.A (n_4340), .B (n_4262), .Y (n_4589));
NAND2X1 g14464(.A (n_5203), .B (n_4408), .Y (n_4414));
INVX1 g14465(.A (n_6478), .Y (n_4413));
NAND2X1 g14469(.A (n_7488), .B (n_4404), .Y (n_4412));
INVX1 g14481(.A (n_5092), .Y (n_4410));
NAND2X1 g14484(.A (n_4282), .B (n_4408), .Y (n_4409));
NAND2X1 g14496(.A (n_4405), .B (n_4404), .Y (n_4406));
NAND2X1 g14499(.A (n_4647), .B (n_4403), .Y (n_5041));
INVX1 g14517(.A (n_4230), .Y (n_5129));
NAND2X1 g14532(.A (n_6530), .B (n_4400), .Y (n_6040));
NAND2X1 g14533(.A (n_4245), .B (n_6888), .Y (n_5062));
INVX1 g14534(.A (n_4398), .Y (n_4399));
NOR2X1 g14557(.A (n_4285), .B (n_4545), .Y (n_6100));
NAND2X1 g14562(.A (n_7359), .B (n_6965), .Y (n_4395));
NAND2X1 g14565(.A (n_4540), .B (n_4539), .Y (n_4394));
INVX1 g14575(.A (n_4392), .Y (n_4393));
INVX1 g14578(.A (n_4390), .Y (n_4391));
INVX1 g14597(.A (n_4389), .Y (n_4797));
NOR2X1 g14601(.A (n_4179), .B (n_5624), .Y (n_4388));
AND2X1 g14617(.A (n_4180), .B (n_5938), .Y (n_4387));
NAND2X1 g14629(.A (n_6450), .B (n_4400), .Y (n_4386));
INVX1 g14678(.A (n_4408), .Y (n_4384));
NAND2X1 g14696(.A (n_4325), .B (n_7320), .Y (n_4576));
NOR2X1 g14700(.A (n_7322), .B (n_7367), .Y (n_4574));
INVX1 g14713(.A (n_4403), .Y (n_4381));
NAND2X1 g13938(.A (n_4380), .B (n_6942), .Y (n_5099));
AND2X1 g14734(.A (n_4378), .B (n_7711), .Y (n_4570));
NOR2X1 g14737(.A (n_6816), .B (n_7358), .Y (n_4580));
INVX1 g14743(.A (n_4375), .Y (n_6095));
INVX4 g14793(.A (n_4554), .Y (n_4908));
INVX4 g14799(.A (n_4554), .Y (n_5121));
NAND2X1 g13961(.A (n_4480), .B (n_6942), .Y (n_4368));
INVX1 g14843(.A (n_4366), .Y (n_4365));
INVX1 g14871(.A (n_4627), .Y (n_4923));
INVX2 g14913(.A (n_4955), .Y (n_4784));
INVX1 g15034(.A (n_5428), .Y (n_5445));
INVX1 g15093(.A (n_4356), .Y (n_5361));
INVX4 g15146(.A (n_3994), .Y (n_5203));
INVX1 g15214(.A (n_4660), .Y (n_4635));
NAND2X1 g14149(.A (n_4526), .B (n_4336), .Y (n_4350));
NAND2X1 g14151(.A (n_3926), .B (n_4346), .Y (n_5104));
NAND2X1 g14156(.A (n_4561), .B (n_4322), .Y (n_4349));
NAND2X1 g14157(.A (n_5166), .B (n_4341), .Y (n_4348));
NAND2X1 g14168(.A (n_4337), .B (n_4346), .Y (n_4983));
NAND4X1 g14169(.A (n_4345), .B (n_3913), .C (n_3768), .D (n_4343), .Y(n_4739));
NAND4X1 g14171(.A (n_4342), .B (n_3913), .C (n_4344), .D (n_4343), .Y(n_5034));
NAND2X1 g14174(.A (n_4342), .B (n_4341), .Y (n_4524));
NAND3X1 g14176(.A (n_3913), .B (n_4340), .C (n_4334), .Y (n_4521));
INVX1 g14177(.A (n_4736), .Y (n_4339));
NAND2X1 g14202(.A (n_4337), .B (n_4336), .Y (n_4338));
NAND3X1 g14203(.A (n_4034), .B (n_4334), .C (n_3985), .Y (n_4335));
NAND2X1 g14205(.A (n_4533), .B (n_4332), .Y (n_4333));
INVX1 g14227(.A (n_4562), .Y (n_4330));
NOR2X1 g14241(.A (n_4022), .B (n_4328), .Y (n_4487));
NAND2X1 g14246(.A (n_4328), .B (n_4063), .Y (n_4329));
NOR2X1 g14247(.A (n_4326), .B (n_4095), .Y (n_4327));
NAND2X1 g14252(.A (n_4325), .B (n_4083), .Y (n_4485));
NAND2X1 g14254(.A (n_6441), .B (n_4634), .Y (n_6062));
NAND2X2 g14256(.A (n_4323), .B (n_4322), .Y (n_4737));
NAND2X2 g14264(.A (n_4035), .B (n_4109), .Y (n_4478));
NAND2X1 g14266(.A (n_4337), .B (n_4341), .Y (n_4671));
NAND4X1 g14271(.A (n_3967), .B (n_3934), .C (n_7614), .D (n_4064), .Y(n_4754));
NAND2X2 g14274(.A (n_4320), .B (n_4316), .Y (n_4934));
NOR2X1 g14275(.A (n_4319), .B (n_4075), .Y (n_4841));
INVX2 g14280(.A (n_4832), .Y (n_4711));
NAND2X1 g14283(.A (n_7248), .B (n_4828), .Y (n_4473));
NAND2X1 g14284(.A (n_6400), .B (n_4317), .Y (n_4709));
NAND2X1 g14286(.A (n_4456), .B (n_4080), .Y (n_4471));
NAND2X1 g14291(.A (n_4316), .B (n_4066), .Y (n_4467));
NAND2X1 g14294(.A (n_4476), .B (n_4314), .Y (n_4315));
NAND2X1 g14298(.A (n_4312), .B (n_4069), .Y (n_4313));
NAND2X1 g14304(.A (n_3962), .B (n_4311), .Y (n_4698));
INVX1 g14307(.A (n_4582), .Y (n_4310));
INVX1 g14311(.A (n_4309), .Y (n_4705));
NAND4X1 g14315(.A (n_4476), .B (n_4073), .C (n_7614), .D (n_4312), .Y(n_4885));
INVX1 g14316(.A (n_4308), .Y (n_4763));
INVX1 g14318(.A (n_4306), .Y (n_4307));
NAND2X1 g14322(.A (n_6047), .B (n_4065), .Y (n_4459));
NAND2X1 g14325(.A (n_4302), .B (n_3962), .Y (n_4457));
INVX1 g14326(.A (n_4300), .Y (n_4301));
NAND4X1 g14333(.A (n_7680), .B (n_4060), .C (n_7606), .D (n_7681), .Y(n_4714));
NAND2X1 g14334(.A (n_4212), .B (n_4302), .Y (n_4669));
NOR2X1 g14336(.A (n_4014), .B (n_4287), .Y (n_4864));
NAND2X2 g14339(.A (n_4067), .B (n_7239), .Y (n_4694));
NAND2X1 g14343(.A (n_4056), .B (n_7358), .Y (n_4296));
NAND2X2 g14346(.A (n_4456), .B (n_4314), .Y (n_4883));
INVX1 g14349(.A (n_4294), .Y (n_4446));
INVX1 g14353(.A (n_6707), .Y (n_4293));
INVX1 g14358(.A (n_4548), .Y (n_6009));
NOR2X1 g14361(.A (n_3929), .B (n_4287), .Y (n_4441));
NAND3X1 g14364(.A (n_4285), .B (n_3931), .C (n_4120), .Y (n_4286));
NOR2X1 g14373(.A (n_3975), .B (n_4090), .Y (n_4284));
AOI21X1 g14377(.A0 (n_4282), .A1 (n_4041), .B0 (n_4281), .Y (n_6094));
NOR2X1 g14408(.A (n_7492), .B (n_6615), .Y (n_4280));
NAND2X1 g14414(.A (n_3870), .B (n_6660), .Y (n_4427));
NOR2X1 g14417(.A (n_4278), .B (n_6743), .Y (n_4279));
INVX1 g14419(.A (n_4276), .Y (n_4277));
INVX1 g14421(.A (n_4274), .Y (n_4275));
NAND2X1 g14425(.A (n_4342), .B (n_4267), .Y (n_4424));
INVX1 g14427(.A (n_4111), .Y (n_4661));
INVX1 g14429(.A (n_4272), .Y (n_4273));
INVX1 g14435(.A (n_4271), .Y (n_4732));
NOR2X1 g14444(.A (n_6988), .B (n_4269), .Y (n_4270));
NOR2X1 g14446(.A (n_6985), .B (n_6890), .Y (n_4420));
NAND2X1 g14450(.A (n_3850), .B (n_4267), .Y (n_4268));
NAND2X1 g14455(.A (n_6531), .B (n_4211), .Y (n_4264));
NAND2X1 g14456(.A (n_4343), .B (n_4262), .Y (n_4263));
INVX1 g14459(.A (n_4261), .Y (n_4608));
NAND2X1 g14461(.A (n_4342), .B (n_4243), .Y (n_4260));
INVX1 g14467(.A (n_4256), .Y (n_4257));
NOR2X1 g14470(.A (n_6822), .B (n_4022), .Y (n_4644));
NAND2X2 g14482(.A (n_6007), .B (n_4052), .Y (n_5092));
NOR2X1 g14483(.A (n_4282), .B (n_4042), .Y (n_4679));
NAND2X1 g14488(.A (n_4252), .B (n_4236), .Y (n_4253));
NAND2X1 g14489(.A (n_6472), .B (n_6673), .Y (n_4650));
NAND2X1 g14613(.A (n_4202), .B (n_4055), .Y (n_4250));
INVX1 g14490(.A (n_4501), .Y (n_4249));
INVX1 g14494(.A (n_4247), .Y (n_4645));
NAND2X1 g14500(.A (n_4245), .B (n_4049), .Y (n_7774));
NAND2X1 g14501(.A (n_4243), .B (n_4233), .Y (n_4244));
NAND2X1 g14502(.A (n_4241), .B (n_5977), .Y (n_4242));
NAND2X1 g14508(.A (n_4252), .B (n_6673), .Y (n_4239));
AND2X1 g14511(.A (n_4237), .B (n_4236), .Y (n_4238));
NAND2X1 g14512(.A (n_4343), .B (n_4233), .Y (n_4235));
NAND2X1 g14515(.A (n_4187), .B (n_6472), .Y (n_4231));
NAND3X1 g14518(.A (n_4482), .B (n_4125), .C (n_3924), .Y (n_4230));
INVX1 g14526(.A (n_4227), .Y (n_4228));
INVX2 g14528(.A (n_4514), .Y (n_4226));
INVX1 g14535(.A (n_4223), .Y (n_4398));
NAND2X1 g14542(.A (n_6988), .B (n_4781), .Y (n_4222));
NAND2X1 g14544(.A (n_6441), .B (n_3980), .Y (n_4220));
INVX1 g14551(.A (n_4218), .Y (n_4219));
INVX1 g14566(.A (n_4604), .Y (n_4217));
NAND2X1 g14568(.A (n_4161), .B (n_4319), .Y (n_4216));
NOR2X1 g14569(.A (n_4161), .B (n_4214), .Y (n_4215));
INVX1 g14570(.A (n_4479), .Y (n_4213));
NAND2X1 g14576(.A (n_3832), .B (n_4212), .Y (n_4392));
NAND2X1 g14579(.A (n_6450), .B (n_4211), .Y (n_4390));
NOR2X1 g14580(.A (n_7464), .B (n_6966), .Y (n_4210));
INVX1 g14581(.A (n_3887), .Y (n_4873));
INVX1 g14587(.A (n_4469), .Y (n_4207));
NAND2X1 g14593(.A (n_4540), .B (n_7249), .Y (n_4206));
INVX1 g14594(.A (n_4065), .Y (n_7900));
NAND2X1 g14598(.A (n_4212), .B (n_3966), .Y (n_4389));
INVX1 g14602(.A (n_4204), .Y (n_4861));
NAND2X1 g14606(.A (n_6817), .B (n_4443), .Y (n_4795));
NAND2X1 g14608(.A (n_4202), .B (n_4282), .Y (n_4203));
NOR2X1 g14614(.A (n_6476), .B (n_4031), .Y (n_4199));
INVX1 g14618(.A (n_4197), .Y (n_4198));
INVX1 g14643(.A (n_4243), .Y (n_4195));
AND2X1 g14650(.A (n_4854), .B (n_6999), .Y (n_4191));
NOR2X1 g14655(.A (n_4055), .B (n_4182), .Y (n_4189));
INVX1 g14658(.A (n_4187), .Y (n_4188));
NOR2X1 g14675(.A (n_3844), .B (n_4182), .Y (n_4183));
INVX1 g14679(.A (n_4043), .Y (n_4408));
NAND2X1 g14705(.A (n_3897), .B (n_4180), .Y (n_4181));
NAND2X1 g14707(.A (n_7252), .B (n_7357), .Y (n_4179));
NAND2X1 g14708(.A (n_3768), .B (n_3984), .Y (n_4178));
INVX1 g14709(.A (n_4439), .Y (n_4177));
INVX1 g14712(.A (n_6615), .Y (n_4176));
INVX1 g14714(.A (n_6615), .Y (n_4403));
NOR2X1 g14729(.A (n_4055), .B (n_4727), .Y (n_4404));
INVX1 g14741(.A (n_4027), .Y (n_4400));
NAND2X1 g14744(.A (n_3988), .B (n_3764), .Y (n_4375));
INVX1 g14749(.A (n_5225), .Y (n_4976));
INVX1 g14772(.A (n_6327), .Y (n_4172));
INVX1 g14774(.A (n_6327), .Y (n_5426));
INVX2 g14783(.A (n_4323), .Y (n_4542));
INVX8 g14789(.A (n_6743), .Y (n_4554));
INVX1 g14822(.A (n_6966), .Y (n_4164));
INVX1 g14844(.A (n_4212), .Y (n_4366));
INVX2 g14866(.A (n_4551), .Y (n_4632));
INVX2 g14872(.A (n_4544), .Y (n_4627));
INVX1 g14876(.A (n_4159), .Y (n_4158));
CLKBUFX3 g14877(.A (n_4159), .Y (n_4875));
INVX2 g14955(.A (n_6151), .Y (n_5404));
INVX1 g15035(.A (n_4142), .Y (n_5428));
INVX1 g15094(.A (n_6786), .Y (n_4356));
INVX4 g15115(.A (n_6400), .Y (n_4539));
INVX1 g15160(.A (n_4498), .Y (n_4133));
INVX2 g15215(.A (n_4325), .Y (n_4660));
NAND3X1 g14178(.A (n_7604), .B (n_4126), .C (n_4125), .Y (n_4736));
INVX1 g14192(.A (n_6942), .Y (n_4124));
NOR2X1 g14228(.A (n_7706), .B (n_7604), .Y (n_4562));
NAND2X2 g14281(.A (n_4067), .B (n_4317), .Y (n_4832));
NOR2X1 g14300(.A (n_7247), .B (n_3969), .Y (n_7741));
NAND3X1 g14308(.A (n_3909), .B (n_6817), .C (n_5624), .Y (n_4582));
NOR2X1 g14312(.A (n_4120), .B (n_4119), .Y (n_4309));
NOR2X1 g14317(.A (n_4012), .B (n_4118), .Y (n_4308));
NOR2X1 g14320(.A (n_4120), .B (n_4116), .Y (n_4306));
NOR2X1 g14327(.A (n_4120), .B (n_4118), .Y (n_4300));
NOR2X1 g14328(.A (n_4537), .B (n_4116), .Y (n_4117));
NOR2X1 g14350(.A (n_7252), .B (n_7381), .Y (n_4294));
NOR2X1 g14359(.A (n_4116), .B (n_4012), .Y (n_4548));
NOR2X1 g14409(.A (n_6464), .B (n_4078), .Y (n_4114));
NAND2X1 g14418(.A (n_4126), .B (n_6661), .Y (n_4516));
NAND2X1 g14420(.A (n_4345), .B (n_3954), .Y (n_4276));
NAND2X1 g14422(.A (n_4214), .B (n_7169), .Y (n_4274));
NAND2X1 g14428(.A (n_6822), .B (n_6742), .Y (n_4111));
INVX1 g14430(.A (n_4109), .Y (n_4272));
INVX1 g14432(.A (n_4346), .Y (n_4108));
NOR2X1 g14436(.A (n_4047), .B (n_4104), .Y (n_4271));
NAND2X2 g14441(.A (n_4340), .B (n_4233), .Y (n_4435));
NOR2X1 g14442(.A (n_3984), .B (n_6385), .Y (n_4107));
INVX2 g14453(.A (n_4106), .Y (n_4105));
NOR2X1 g14460(.A (n_4104), .B (n_6385), .Y (n_4261));
NAND2X1 g14468(.A (n_4241), .B (n_3956), .Y (n_4256));
NOR2X1 g14480(.A (n_4038), .B (n_4097), .Y (n_4255));
INVX2 g14485(.A (n_4099), .Y (n_4599));
NOR2X1 g14492(.A (n_4098), .B (n_4055), .Y (n_4501));
NOR2X1 g14495(.A (n_4097), .B (n_4061), .Y (n_4247));
NAND2X1 g14497(.A (n_3919), .B (n_4039), .Y (n_4096));
INVX1 g14504(.A (n_4095), .Y (n_4490));
INVX1 g14506(.A (n_4326), .Y (n_4488));
NAND2X1 g14510(.A (n_4093), .B (n_4094), .Y (n_4492));
NAND2X2 g14514(.A (n_4093), .B (n_3976), .Y (n_4676));
NAND2X2 g14516(.A (n_4092), .B (n_4677), .Y (n_4596));
INVX1 g14520(.A (n_4090), .Y (n_4091));
INVX1 g14524(.A (n_4558), .Y (n_4088));
NAND3X1 g14527(.A (n_6986), .B (n_6531), .C (n_6994), .Y (n_4227));
NAND2X2 g14531(.A (n_6985), .B (n_6891), .Y (n_4514));
NOR2X1 g14536(.A (n_6985), .B (n_4269), .Y (n_4223));
INVX1 g14540(.A (n_4083), .Y (n_4082));
INVX1 g14545(.A (n_4080), .Y (n_7753));
NOR2X1 g14547(.A (n_3970), .B (n_4060), .Y (n_4477));
NAND2X1 g14548(.A (n_3962), .B (n_3947), .Y (n_4079));
NOR2X1 g14552(.A (n_4028), .B (n_4078), .Y (n_4218));
INVX1 g14553(.A (n_4311), .Y (n_4077));
INVX1 g14555(.A (n_4075), .Y (n_7890));
NOR2X1 g14558(.A (n_4073), .B (n_3973), .Y (n_4074));
INVX1 g14563(.A (n_4069), .Y (n_7800));
NAND2X2 g14567(.A (n_4067), .B (n_4068), .Y (n_4604));
NAND2X1 g14571(.A (n_3890), .B (n_7604), .Y (n_4479));
NOR2X1 g14588(.A (n_7606), .B (n_4073), .Y (n_4469));
NOR2X1 g14599(.A (n_4064), .B (n_3934), .Y (n_4451));
INVX1 g14603(.A (n_4063), .Y (n_4204));
NAND2X1 g14605(.A (n_4344), .B (n_4233), .Y (n_4062));
NOR2X1 g14607(.A (n_6875), .B (n_4061), .Y (n_4528));
NOR2X1 g14620(.A (n_4060), .B (n_4059), .Y (n_4197));
NAND2X1 g14621(.A (n_6476), .B (n_4030), .Y (n_4058));
INVX1 g14625(.A (n_4056), .Y (n_4057));
NOR2X1 g14638(.A (n_3855), .B (n_7492), .Y (n_4054));
NOR2X1 g14639(.A (n_4052), .B (n_4728), .Y (n_4202));
INVX1 g14644(.A (n_6385), .Y (n_4243));
INVX1 g14648(.A (n_4049), .Y (n_4193));
INVX1 g14651(.A (n_4093), .Y (n_4236));
NOR2X1 g14659(.A (n_3977), .B (n_5711), .Y (n_4187));
INVX1 g14670(.A (n_4047), .Y (n_4267));
INVX1 g14672(.A (n_4092), .Y (n_4046));
INVX1 g14676(.A (n_4044), .Y (n_4045));
NAND2X1 g14680(.A (n_4052), .B (n_7492), .Y (n_4043));
INVX1 g14681(.A (n_4041), .Y (n_4042));
INVX1 g14687(.A (n_4039), .Y (n_4040));
INVX1 g14710(.A (n_4038), .Y (n_4439));
INVX1 g14717(.A (n_6674), .Y (n_4037));
NOR2X1 g14720(.A (n_6988), .B (n_3764), .Y (n_4211));
NAND2X1 g14723(.A (n_4344), .B (n_4036), .Y (n_4332));
NOR2X1 g14725(.A (n_4035), .B (n_4034), .Y (n_4262));
INVX2 g14727(.A (n_4061), .Y (n_6007));
INVX1 g14730(.A (n_4030), .Y (n_4031));
NAND2X1 g14732(.A (n_4252), .B (n_4028), .Y (n_4029));
NAND2X1 g14742(.A (n_6988), .B (n_6985), .Y (n_4027));
INVX1 g14747(.A (n_4743), .Y (n_5214));
INVX2 g14750(.A (n_4025), .Y (n_5225));
INVX1 g14776(.A (n_6661), .Y (n_4482));
INVX1 g14778(.A (n_6661), .Y (n_4022));
CLKBUFX3 g14784(.A (n_6661), .Y (n_4323));
INVX4 g14845(.A (n_4060), .Y (n_4212));
INVX2 g14857(.A (n_4285), .Y (n_4161));
INVX2 g14863(.A (n_4214), .Y (n_4545));
INVX4 g14867(.A (n_4014), .Y (n_4551));
INVX2 g14873(.A (n_4537), .Y (n_4544));
INVX2 g14878(.A (n_4013), .Y (n_4159));
INVX1 g14883(.A (n_4319), .Y (n_4665));
INVX2 g14885(.A (n_4012), .Y (n_4316));
INVX1 g14922(.A (n_4854), .Y (n_5166));
INVX4 g14938(.A (n_4380), .Y (n_4561));
INVX4 g14940(.A (n_4278), .Y (n_4480));
INVX1 g14959(.A (n_6530), .Y (n_4594));
INVX1 g14995(.A (n_4430), .Y (n_4823));
INVX1 g15004(.A (n_7490), .Y (n_4145));
INVX1 g15019(.A (n_4814), .Y (n_5059));
AOI21X1 g15037(.A0 (n_3830), .A1 (n_3829), .B0 (n_3831), .Y (n_4142));
INVX1 g15128(.A (n_7248), .Y (n_7760));
INVX1 g15153(.A (n_4727), .Y (n_4134));
INVX2 g15163(.A (n_4849), .Y (n_4498));
INVX2 g15212(.A (n_3988), .Y (n_4245));
CLKBUFX3 g15216(.A (n_3988), .Y (n_4325));
INVX2 g15258(.A (n_4180), .Y (n_4449));
INVX1 g14415(.A (n_4328), .Y (n_4719));
NOR2X1 g14431(.A (n_3942), .B (n_3985), .Y (n_4109));
NOR2X1 g14433(.A (n_3983), .B (n_4104), .Y (n_4346));
NOR2X1 g14439(.A (n_4034), .B (n_3985), .Y (n_4336));
NAND3X1 g14440(.A (n_4343), .B (n_4035), .C (n_3984), .Y (n_4533));
NOR2X1 g14443(.A (n_3984), .B (n_3983), .Y (n_4341));
INVX1 g14448(.A (n_6748), .Y (n_3982));
NAND2X2 g14454(.A (n_6985), .B (n_3980), .Y (n_4106));
INVX1 g14471(.A (n_4322), .Y (n_3978));
NOR2X1 g14487(.A (n_3974), .B (n_7797), .Y (n_4099));
NOR2X1 g14505(.A (n_3976), .B (n_3977), .Y (n_4095));
NOR2X1 g14507(.A (n_6479), .B (n_3976), .Y (n_4326));
NOR2X1 g14519(.A (n_5711), .B (n_3872), .Y (n_3975));
NOR2X1 g14521(.A (n_3946), .B (n_3974), .Y (n_4090));
NOR2X1 g14525(.A (n_6470), .B (n_3974), .Y (n_4558));
NOR2X1 g14541(.A (n_3764), .B (n_3948), .Y (n_4083));
NOR2X1 g14546(.A (n_3971), .B (n_3973), .Y (n_4080));
NAND2X1 g14549(.A (n_4476), .B (n_3875), .Y (n_3972));
NOR2X1 g14554(.A (n_3971), .B (n_3970), .Y (n_4311));
NAND2X1 g14556(.A (n_3930), .B (n_6048), .Y (n_4075));
NOR2X1 g14564(.A (n_3971), .B (n_7681), .Y (n_4069));
INVX1 g14573(.A (n_3969), .Y (n_4828));
NOR2X1 g14577(.A (n_3962), .B (n_3973), .Y (n_3968));
INVX1 g14583(.A (n_3887), .Y (n_4066));
INVX1 g14585(.A (n_4119), .Y (n_4320));
NAND2X1 g14589(.A (n_3967), .B (n_3966), .Y (n_4839));
INVX1 g14590(.A (n_4118), .Y (n_3965));
NOR2X1 g14596(.A (n_3958), .B (n_4120), .Y (n_4065));
NAND2X1 g14600(.A (n_3962), .B (n_3966), .Y (n_7754));
NAND2X1 g14604(.A (n_7603), .B (n_3890), .Y (n_4063));
NAND2X1 g14615(.A (n_4028), .B (n_4237), .Y (n_3960));
NOR2X1 g14616(.A (n_3971), .B (n_3957), .Y (n_4314));
INVX1 g14626(.A (n_6706), .Y (n_4056));
NAND2X1 g14631(.A (n_3958), .B (n_4120), .Y (n_4287));
NAND2X2 g14632(.A (n_3957), .B (n_4059), .Y (n_4302));
INVX1 g14641(.A (n_3983), .Y (n_4050));
NOR2X1 g14649(.A (n_6454), .B (n_6985), .Y (n_4049));
NAND2X2 g14652(.A (n_5713), .B (n_6475), .Y (n_4093));
INVX1 g14653(.A (n_3976), .Y (n_3956));
NAND2X1 g14656(.A (n_3953), .B (n_7308), .Y (n_4098));
NOR2X1 g14657(.A (n_4035), .B (n_3861), .Y (n_4334));
NAND2X2 g14666(.A (n_6454), .B (n_6991), .Y (n_4269));
INVX1 g14667(.A (n_3985), .Y (n_3954));
NAND2X1 g14671(.A (n_6384), .B (n_6386), .Y (n_4047));
INVX2 g14673(.A (n_3974), .Y (n_4092));
NAND2X1 g14677(.A (n_3953), .B (n_3950), .Y (n_4044));
NOR2X1 g14682(.A (n_4097), .B (n_7492), .Y (n_4041));
NOR2X1 g14686(.A (n_3953), .B (n_3950), .Y (n_4281));
NOR2X1 g14688(.A (n_3844), .B (n_7492), .Y (n_4039));
NAND2X1 g14691(.A (n_5713), .B (n_6469), .Y (n_4094));
INVX1 g14692(.A (n_3980), .Y (n_4289));
INVX1 g14697(.A (n_3948), .Y (n_4781));
INVX1 g14703(.A (n_3973), .Y (n_3947));
NAND2X1 g14711(.A (n_3797), .B (n_6461), .Y (n_4038));
NAND2X1 g14716(.A (n_3946), .B (n_3945), .Y (n_4078));
NAND2X2 g14728(.A (n_6613), .B (n_6461), .Y (n_4061));
NOR2X1 g14731(.A (n_3946), .B (n_6471), .Y (n_4030));
NOR2X1 g14736(.A (n_3771), .B (n_3942), .Y (n_4233));
INVX1 g14745(.A (n_4059), .Y (n_3941));
INVX1 g14748(.A (n_7169), .Y (n_4743));
INVX1 g14751(.A (n_7169), .Y (n_4025));
INVX1 g14803(.A (n_4540), .Y (n_3938));
INVX2 g14814(.A (n_6817), .Y (n_4068));
INVX4 g14846(.A (n_3971), .Y (n_4060));
INVX1 g14849(.A (n_3971), .Y (n_4073));
INVX2 g14850(.A (n_3971), .Y (n_3934));
INVX4 g14859(.A (n_3958), .Y (n_4285));
INVX2 g14864(.A (n_3932), .Y (n_4214));
INVX2 g14868(.A (n_3932), .Y (n_4014));
INVX1 g14869(.A (n_3932), .Y (n_3931));
INVX2 g14874(.A (n_3930), .Y (n_4537));
INVX2 g14879(.A (n_3930), .Y (n_4013));
INVX1 g14880(.A (n_3930), .Y (n_3929));
INVX1 g14884(.A (n_4120), .Y (n_4319));
INVX4 g14886(.A (n_4120), .Y (n_4012));
INVX2 g14917(.A (n_3926), .Y (n_4955));
CLKBUFX1 g14918(.A (n_3926), .Y (n_4526));
INVX4 g14923(.A (n_4345), .Y (n_4854));
INVX2 g14932(.A (n_3924), .Y (n_4541));
INVX4 g14939(.A (n_3924), .Y (n_4380));
INVX4 g14942(.A (n_3924), .Y (n_4278));
INVX4 g14977(.A (n_4343), .Y (n_4340));
INVX1 g14984(.A (n_4405), .Y (n_4182));
INVX1 g14985(.A (n_4405), .Y (n_3919));
INVX1 g14996(.A (n_7492), .Y (n_4430));
INVX1 g15020(.A (n_7320), .Y (n_4814));
INVX2 g15061(.A (n_4036), .Y (n_3913));
INVX2 g15069(.A (n_7462), .Y (n_4443));
INVX4 g15121(.A (n_3909), .Y (n_4067));
INVX4 g15150(.A (n_6875), .Y (n_3994));
INVX4 g15154(.A (n_6876), .Y (n_4727));
INVX2 g15164(.A (n_4378), .Y (n_4849));
CLKBUFX1 g15202(.A (n_7142), .Y (n_5419));
INVX1 g15203(.A (n_7142), .Y (n_3899));
INVX4 g15217(.A (n_6988), .Y (n_3988));
INVX4 g15259(.A (n_3962), .Y (n_4180));
INVX1 g15267(.A (n_3896), .Y (n_3897));
NAND2X1 g15320(.A (n_3892), .B (n_3891), .Y (n_3894));
OR2X1 g15321(.A (n_3892), .B (n_3891), .Y (n_3893));
NAND2X2 g14416(.A (n_3821), .B (n_3890), .Y (n_4328));
INVX2 g14474(.A (n_3827), .Y (n_4322));
NOR2X1 g14522(.A (n_6985), .B (n_3876), .Y (n_4634));
NOR2X1 g14572(.A (n_7382), .B (n_6705), .Y (n_4317));
NAND2X2 g14574(.A (n_6705), .B (n_7382), .Y (n_3969));
NAND2X1 g14584(.A (n_3885), .B (n_6049), .Y (n_3887));
NAND2X2 g14586(.A (n_3883), .B (n_6050), .Y (n_4119));
NAND2X2 g14592(.A (n_3885), .B (n_6050), .Y (n_4118));
NAND2X2 g14630(.A (n_3883), .B (n_6049), .Y (n_4116));
NAND2X2 g14642(.A (n_6383), .B (n_6386), .Y (n_3983));
NAND2X2 g14654(.A (n_6583), .B (n_6474), .Y (n_3976));
NAND2X1 g14665(.A (n_3772), .B (n_6990), .Y (n_3879));
NAND2X2 g14668(.A (n_6383), .B (n_6382), .Y (n_3985));
NAND2X2 g14674(.A (n_6010), .B (n_6583), .Y (n_3974));
INVX1 g14693(.A (n_3876), .Y (n_3980));
NAND2X1 g14698(.A (n_6529), .B (n_3738), .Y (n_3948));
INVX1 g14701(.A (n_3970), .Y (n_3875));
NAND2X2 g14704(.A (n_4064), .B (n_7608), .Y (n_3973));
INVX1 g14721(.A (n_3957), .Y (n_3966));
NOR2X1 g14724(.A (n_6992), .B (n_6986), .Y (n_3873));
INVX1 g14738(.A (n_3872), .Y (n_4237));
NAND2X2 g14746(.A (n_3824), .B (n_7614), .Y (n_4059));
INVX2 g14768(.A (n_4126), .Y (n_3870));
INVX1 g14804(.A (n_6818), .Y (n_4540));
INVX1 g14806(.A (n_6818), .Y (n_5624));
INVX4 g14852(.A (n_3818), .Y (n_3971));
INVX4 g14860(.A (n_3885), .Y (n_3958));
INVX2 g14870(.A (n_3866), .Y (n_3932));
CLKBUFX3 g14881(.A (n_3866), .Y (n_3930));
INVX4 g14889(.A (n_3816), .Y (n_4120));
NAND2X1 g14891(.A (n_3863), .B (n_6215), .Y (n_3865));
OR2X1 g14892(.A (n_3863), .B (n_6215), .Y (n_3864));
INVX2 g14919(.A (n_3861), .Y (n_3926));
INVX2 g14924(.A (n_3861), .Y (n_4345));
INVX4 g14943(.A (n_3860), .Y (n_3924));
CLKBUFX3 g14978(.A (n_6384), .Y (n_4343));
CLKBUFX3 g14986(.A (n_3950), .Y (n_4405));
INVX1 g14987(.A (n_3950), .Y (n_4052));
INVX1 g14990(.A (n_4097), .Y (n_3855));
CLKBUFX3 g15000(.A (n_7492), .Y (n_4647));
INVX4 g15001(.A (n_7492), .Y (n_4728));
INVX4 g15042(.A (n_4337), .Y (n_4813));
INVX1 g15044(.A (n_3851), .Y (n_4509));
INVX1 g15045(.A (n_3851), .Y (n_3850));
INVX2 g15057(.A (n_3984), .Y (n_4034));
INVX1 g15060(.A (n_3942), .Y (n_4104));
CLKBUFX3 g15064(.A (n_3942), .Y (n_4036));
INVX4 g15123(.A (n_6816), .Y (n_3909));
INVX1 g15138(.A (n_6476), .Y (n_4028));
INVX2 g15165(.A (n_3946), .Y (n_4378));
INVX4 g15178(.A (n_3844), .Y (n_4055));
CLKBUFX1 g15182(.A (n_3953), .Y (n_4282));
INVX2 g15236(.A (n_4504), .Y (n_4637));
INVX2 g15249(.A (n_3967), .Y (n_4456));
INVX1 g15252(.A (n_4476), .Y (n_4619));
INVX4 g15260(.A (n_3834), .Y (n_3962));
INVX2 g15269(.A (n_3832), .Y (n_3896));
NOR2X1 g15287(.A (n_3830), .B (n_3829), .Y (n_3831));
NAND2X1 g14475(.A (n_6944), .B (n_6943), .Y (n_3827));
NAND2X1 g14694(.A (n_6533), .B (n_6990), .Y (n_3876));
NAND2X1 g14702(.A (n_3824), .B (n_7607), .Y (n_3970));
NAND2X2 g14722(.A (n_3737), .B (n_7607), .Y (n_3957));
NAND2X1 g14739(.A (n_3766), .B (n_6479), .Y (n_3872));
INVX1 g14763(.A (n_6944), .Y (n_3821));
INVX4 g14769(.A (n_6944), .Y (n_4126));
NAND2X2 g14853(.A (n_3712), .B (n_3746), .Y (n_3818));
CLKBUFX2 g14854(.A (n_3817), .Y (n_3883));
INVX2 g14861(.A (n_3817), .Y (n_3885));
NAND2X2 g14882(.A (n_3708), .B (n_3745), .Y (n_3866));
NAND2X2 g14890(.A (n_3707), .B (n_3744), .Y (n_3816));
NAND2X1 g14896(.A (n_3733), .B (desOut[49]), .Y (n_3815));
NAND2X1 g14902(.A (n_3731), .B (desOut[27]), .Y (n_3814));
NAND2X2 g14925(.A (n_3693), .B (n_3734), .Y (n_3861));
INVX2 g14944(.A (n_6821), .Y (n_3860));
INVX2 g14988(.A (n_7308), .Y (n_3950));
INVX1 g15038(.A (n_4035), .Y (n_4342));
CLKBUFX1 g15046(.A (n_3806), .Y (n_3851));
INVX2 g15050(.A (n_3806), .Y (n_4337));
CLKBUFX1 g15051(.A (n_3806), .Y (n_4495));
INVX2 g15059(.A (n_3805), .Y (n_3984));
INVX2 g15065(.A (n_3805), .Y (n_3942));
INVX1 g15099(.A (n_4125), .Y (n_4572));
INVX2 g15156(.A (n_3977), .Y (n_4677));
CLKBUFX3 g15158(.A (n_3977), .Y (n_4241));
INVX2 g15166(.A (n_3798), .Y (n_3946));
INVX1 g15170(.A (n_6613), .Y (n_3797));
INVX2 g15179(.A (n_6613), .Y (n_3844));
CLKBUFX1 g15183(.A (n_6614), .Y (n_3953));
CLKBUFX3 g15238(.A (n_3945), .Y (n_4504));
INVX2 g15239(.A (n_3945), .Y (n_4252));
INVX1 g15245(.A (n_6470), .Y (n_7797));
INVX1 g15250(.A (n_6640), .Y (n_3967));
INVX2 g15253(.A (n_6640), .Y (n_4476));
INVX2 g15254(.A (n_6640), .Y (n_7681));
INVX2 g15263(.A (n_6640), .Y (n_3834));
INVX1 g15270(.A (n_4312), .Y (n_3832));
INVX1 g15271(.A (n_4312), .Y (n_3787));
NAND2X1 g15298(.A (n_3729), .B (desOut[21]), .Y (n_3780));
NAND4X1 g15377(.A (n_2662), .B (n_3211), .C (n_3027), .D (n_3624), .Y(n_3892));
OAI21X1 g14862(.A0 (n_3710), .A1 (n_3709), .B0 (n_3711), .Y (n_3817));
NAND2X1 g14900(.A (n_3732), .B (n_2769), .Y (n_3776));
NAND2X1 g14901(.A (n_3730), .B (n_3709), .Y (n_3775));
NAND2X1 g14904(.A (n_3685), .B (desOut[17]), .Y (n_3774));
INVX1 g14965(.A (n_6533), .Y (n_3772));
INVX2 g15040(.A (n_3771), .Y (n_4035));
CLKBUFX2 g15052(.A (n_3771), .Y (n_3806));
INVX2 g15066(.A (n_3742), .Y (n_3805));
INVX1 g15085(.A (n_3768), .Y (n_4344));
INVX2 g15101(.A (n_3890), .Y (n_4125));
INVX2 g15134(.A (n_6474), .Y (n_6010));
INVX2 g15159(.A (n_3766), .Y (n_3977));
INVX2 g15167(.A (n_3766), .Y (n_3798));
INVX2 g15222(.A (n_6985), .Y (n_3764));
INVX1 g15241(.A (n_6469), .Y (n_3945));
INVX1 g15266(.A (n_4064), .Y (n_7680));
INVX2 g15272(.A (n_4064), .Y (n_4312));
NAND2X2 g15281(.A (n_3654), .B (n_3695), .Y (n_3786));
NAND2X1 g15290(.A (n_3754), .B (n_6609), .Y (n_3759));
NAND2X1 g15291(.A (n_3681), .B (n_2870), .Y (n_3758));
NAND2X1 g15296(.A (n_6700), .B (n_2776), .Y (n_3756));
OR2X1 g15300(.A (n_3754), .B (n_6609), .Y (n_3755));
NAND4X1 g15324(.A (n_3430), .B (n_3428), .C (n_2247), .D (n_3588), .Y(n_3863));
NAND4X1 g15352(.A (n_3420), .B (n_3074), .C (n_3310), .D (n_3587), .Y(n_3830));
NOR2X1 g15357(.A (n_3356), .B (n_3678), .Y (n_3752));
NAND4X1 g15396(.A (n_2987), .B (n_3166), .C (n_3164), .D (n_3589), .Y(n_3751));
NAND2X1 g14895(.A (n_6886), .B (desOut[33]), .Y (n_3748));
NAND2X1 g14903(.A (n_7406), .B (n_2790), .Y (n_3747));
NAND2X1 g14906(.A (n_3645), .B (desOut[1]), .Y (n_3746));
NAND2X1 g14909(.A (n_3639), .B (desOut[43]), .Y (n_3745));
NAND2X1 g14911(.A (n_3641), .B (desOut[35]), .Y (n_3744));
MX2X1 g15053(.A (desOut[45]), .B (n_2143), .S0 (n_3614), .Y (n_3771));
MX2X1 g15067(.A (desOut[37]), .B (n_2544), .S0 (n_7300), .Y (n_3742));
INVX1 g15086(.A (n_6382), .Y (n_3768));
CLKBUFX3 g15102(.A (n_6878), .Y (n_3890));
INVX2 g15168(.A (n_3704), .Y (n_3766));
INVX1 g15234(.A (n_6990), .Y (n_3738));
INVX1 g15265(.A (n_3824), .Y (n_3737));
INVX2 g15273(.A (n_3824), .Y (n_4064));
NAND2X1 g15292(.A (n_3680), .B (desOut[23]), .Y (n_3736));
NAND2X1 g15311(.A (n_3637), .B (desOut[53]), .Y (n_3734));
INVX1 g15326(.A (n_3732), .Y (n_3733));
INVX1 g15330(.A (n_3730), .Y (n_3731));
INVX1 g15374(.A (n_6700), .Y (n_3729));
INVX1 g15412(.A (n_3724), .Y (n_3725));
INVX1 g15427(.A (n_3720), .Y (n_3721));
NAND2X1 g14905(.A (n_6604), .B (n_2380), .Y (n_3712));
NAND2X1 g14907(.A (n_3710), .B (n_3709), .Y (n_3711));
NAND2X1 g14908(.A (n_3638), .B (n_2289), .Y (n_3708));
NAND2X1 g14910(.A (n_3640), .B (n_2294), .Y (n_3707));
MX2X1 g15169(.A (n_1897), .B (n_1896), .S0 (n_3576), .Y (n_3704));
INVX2 g15274(.A (n_3658), .Y (n_3824));
NAND2X1 g15307(.A (n_3596), .B (desOut[1]), .Y (n_3695));
NAND2X1 g15310(.A (n_6421), .B (n_2778), .Y (n_3693));
NAND2X1 g15312(.A (n_3613), .B (n_1480), .Y (n_3692));
NAND2X1 g15315(.A (n_3608), .B (desOut[41]), .Y (n_3691));
NAND4X1 g15327(.A (n_3478), .B (n_3229), .C (n_2973), .D (n_3544), .Y(n_3732));
NAND4X1 g15331(.A (n_5666), .B (n_3210), .C (n_3155), .D (n_5667), .Y(n_3730));
INVX1 g15338(.A (n_7406), .Y (n_3685));
NAND4X1 g15341(.A (n_5609), .B (n_3393), .C (n_5610), .D (n_3401), .Y(n_3683));
INVX1 g15353(.A (n_3680), .Y (n_3681));
NAND4X1 g15385(.A (n_3411), .B (n_3227), .C (n_3540), .D (n_3209), .Y(n_3754));
NAND3X1 g15402(.A (n_7520), .B (n_7521), .C (n_2970), .Y (n_3678));
OAI22X1 g15413(.A0 (n_3566), .A1 (n_3677), .B0 (n_3673), .B1 (n_74),.Y (n_3724));
AOI22X1 g15414(.A0 (n_3554), .A1 (n_1776), .B0 (n_3677), .B1(desIn[22]), .Y (n_5523));
INVX1 g15422(.A (n_7156), .Y (n_3675));
OAI22X1 g15428(.A0 (n_3560), .A1 (n_3677), .B0 (n_3673), .B1 (n_18),.Y (n_3720));
INVX1 g15439(.A (n_3669), .Y (n_3670));
INVX1 g15459(.A (n_3666), .Y (n_3667));
INVX1 g15461(.A (n_3664), .Y (n_3665));
MX2X1 g15275(.A (desOut[59]), .B (n_2287), .S0 (n_6435), .Y (n_3658));
NAND2X1 g15306(.A (n_6848), .B (n_2380), .Y (n_3654));
NAND2X1 g15313(.A (n_3612), .B (n_1478), .Y (n_3651));
NAND2X1 g15314(.A (n_6690), .B (n_2781), .Y (n_3650));
INVX1 g15332(.A (n_6604), .Y (n_3645));
INVX1 g15342(.A (n_3640), .Y (n_3641));
INVX1 g15344(.A (n_3638), .Y (n_3639));
NOR2X1 g15354(.A (n_3417), .B (n_7501), .Y (n_3680));
INVX1 g15379(.A (n_6421), .Y (n_3637));
INVX1 g15389(.A (n_3634), .Y (n_3635));
INVX1 g15420(.A (n_3629), .Y (n_3630));
OAI22X1 g15440(.A0 (n_3528), .A1 (n_3677), .B0 (n_1776), .B1 (n_24),.Y (n_3669));
NOR2X1 g15444(.A (n_3029), .B (n_3567), .Y (n_3624));
OAI22X1 g15460(.A0 (n_3526), .A1 (n_3677), .B0 (n_1776), .B1 (n_25),.Y (n_3666));
OAI22X1 g15462(.A0 (n_3524), .A1 (n_3677), .B0 (n_3673), .B1 (n_15),.Y (n_3664));
AOI22X1 g15511(.A0 (n_3549), .A1 (n_1776), .B0 (n_3677), .B1(desIn[54]), .Y (n_5526));
NAND2X1 g14897(.A (n_7092), .B (n_2294), .Y (n_3617));
NAND4X1 g15340(.A (n_5641), .B (n_2682), .C (n_5642), .D (n_2684), .Y(n_3710));
NAND4X1 g15343(.A (n_3346), .B (n_3192), .C (n_3498), .D (n_3006), .Y(n_3640));
NAND4X1 g15345(.A (n_3516), .B (n_3195), .C (n_3494), .D (n_2676), .Y(n_3638));
NOR2X1 g15348(.A (n_3426), .B (n_6229), .Y (n_3614));
INVX1 g15349(.A (n_3612), .Y (n_3613));
INVX1 g15364(.A (n_6690), .Y (n_3608));
INVX1 g15369(.A (n_3603), .Y (n_3604));
INVX1 g15372(.A (n_3601), .Y (n_3602));
NAND4X1 g15390(.A (n_7784), .B (n_2702), .C (n_7785), .D (n_2708), .Y(n_3634));
INVX1 g15393(.A (n_6848), .Y (n_3596));
NAND4X1 g15401(.A (n_3051), .B (n_2717), .C (n_3481), .D (n_3351), .Y(n_3593));
NAND4X1 g15403(.A (n_3199), .B (n_3314), .C (n_3472), .D (n_3473), .Y(n_3592));
OAI22X1 g15421(.A0 (n_3514), .A1 (n_3677), .B0 (n_3673), .B1 (n_90),.Y (n_3629));
NOR2X1 g15445(.A (n_3323), .B (n_3541), .Y (n_3589));
INVX1 g15452(.A (n_3571), .Y (n_3588));
INVX1 g15487(.A (n_3570), .Y (n_3587));
OR4X1 g15323(.A (n_3585), .B (n_7079), .C (n_7082), .D (n_7076), .Y(n_3586));
NOR2X1 g15350(.A (n_3284), .B (n_6576), .Y (n_3612));
NAND4X1 g15362(.A (n_5591), .B (n_3232), .C (n_5592), .D (n_3050), .Y(n_3578));
NAND4X1 g15370(.A (n_6083), .B (n_6084), .C (n_3444), .D (n_2736), .Y(n_3603));
NAND4X1 g15371(.A (n_3416), .B (n_3041), .C (n_3436), .D (n_3045), .Y(n_3576));
NAND4X1 g15373(.A (n_7790), .B (n_5596), .C (n_7791), .D (n_3039), .Y(n_3601));
NAND4X1 g15453(.A (n_3392), .B (n_3397), .C (n_3429), .D (n_3344), .Y(n_3571));
NAND4X1 g15488(.A (n_3186), .B (n_2766), .C (n_3398), .D (n_3248), .Y(n_3570));
INVX1 g15490(.A (n_6928), .Y (n_7520));
INVX1 g15497(.A (n_3537), .Y (n_3568));
NAND2X1 g15503(.A (n_3512), .B (n_3511), .Y (n_3567));
AOI22X1 g15519(.A0 (n_3468), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_36), .Y (n_3566));
AOI22X1 g15520(.A0 (n_3467), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_53), .Y (n_3565));
MX2X1 g15521(.A (FP_R_45), .B (n_3466), .S0 (n_1260), .Y (n_3564));
MX2X1 g15522(.A (FP_R_37), .B (n_3465), .S0 (n_1260), .Y (n_3563));
AOI22X1 g15527(.A0 (n_3507), .A1 (n_1260), .B0 (n_3550), .B1 (n_38),.Y (n_3561));
AOI22X1 g15528(.A0 (n_3510), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_49), .Y (n_3560));
AOI22X1 g15530(.A0 (n_3509), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_41), .Y (n_3558));
AOI22X1 g15533(.A0 (n_3506), .A1 (n_1260), .B0 (n_3550), .B1 (n_7),.Y (n_3557));
MX2X1 g15534(.A (FP_R_61), .B (n_3508), .S0 (n_1260), .Y (n_3554));
MX2X1 g15680(.A (FP_R_33), .B (n_3504), .S0 (n_1260), .Y (n_3553));
AOI22X1 g15683(.A0 (n_3503), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_40), .Y (n_3552));
MX2X1 g16074(.A (FP_R_57), .B (n_3442), .S0 (n_1268), .Y (n_3549));
MX2X1 g16076(.A (FP_R_63), .B (n_3440), .S0 (n_1260), .Y (n_3548));
NOR2X1 g15448(.A (n_3493), .B (n_3421), .Y (n_3544));
NOR2X1 g15449(.A (n_3410), .B (n_3492), .Y (n_5666));
NOR2X1 g15457(.A (n_3491), .B (n_3400), .Y (n_5609));
NAND2X1 g15483(.A (n_3471), .B (n_3403), .Y (n_3541));
NOR2X1 g15484(.A (n_3418), .B (n_3479), .Y (n_3540));
NAND3X1 g15498(.A (n_3480), .B (n_3234), .C (n_2977), .Y (n_3537));
MX2X1 g15517(.A (FP_R_32), .B (n_3460), .S0 (n_1260), .Y (n_3536));
OAI22X1 g15524(.A0 (n_3463), .A1 (n_3550), .B0 (n_1268), .B1(FP_R_46), .Y (n_3535));
MX2X1 g15525(.A (FP_R_38), .B (n_3462), .S0 (n_1260), .Y (n_3534));
MX2X1 g15529(.A (FP_R_39), .B (n_3459), .S0 (n_1260), .Y (n_3532));
MX2X1 g15531(.A (FP_R_58), .B (n_3458), .S0 (n_1260), .Y (n_3531));
AOI22X1 g15535(.A0 (n_3457), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_59), .Y (n_3530));
MX2X1 g15536(.A (FP_R_56), .B (n_3456), .S0 (n_1260), .Y (n_3529));
AOI22X1 g15537(.A0 (n_3455), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_51), .Y (n_3528));
MX2X1 g15538(.A (FP_R_43), .B (n_3454), .S0 (n_1260), .Y (n_3527));
AOI22X1 g15681(.A0 (n_3453), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_48), .Y (n_3526));
AOI22X1 g15682(.A0 (n_3451), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_42), .Y (n_3524));
AOI22X1 g16075(.A0 (n_3387), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_62), .Y (n_3522));
MX2X1 g16077(.A (FP_R_52), .B (n_3377), .S0 (n_1260), .Y (n_3521));
NOR2X1 g15474(.A (n_3399), .B (n_3196), .Y (n_3516));
AOI22X1 g15518(.A0 (n_3313), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_44), .Y (n_3515));
AOI22X1 g15523(.A0 (n_3391), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_54), .Y (n_3514));
MX2X1 g15532(.A (FP_R_50), .B (n_3390), .S0 (n_1260), .Y (n_3513));
NOR2X1 g15616(.A (n_3318), .B (n_3395), .Y (n_3512));
NOR2X1 g15619(.A (n_3394), .B (n_2969), .Y (n_3511));
MX2X1 g16061(.A (L_80), .B (FP_R_49), .S0 (n_7846), .Y (n_3510));
MX2X1 g16062(.A (L_72), .B (FP_R_41), .S0 (n_7846), .Y (n_3509));
MX2X1 g16065(.A (L_92), .B (FP_R_61), .S0 (n_7846), .Y (n_3508));
MX2X1 g16068(.A (L_78), .B (n_38), .S0 (n_7846), .Y (n_3507));
MX2X1 g16069(.A (L_65), .B (n_7), .S0 (n_7846), .Y (n_3506));
MX2X1 g16642(.A (L_64), .B (FP_R_33), .S0 (n_7846), .Y (n_3504));
MX2X1 g16645(.A (L_71), .B (FP_R_40), .S0 (n_7846), .Y (n_3503));
NAND4X1 g15405(.A (n_6101), .B (n_6102), .C (n_5684), .D (n_3080), .Y(n_3501));
NOR2X1 g15447(.A (n_3251), .B (n_3378), .Y (n_3498));
NOR2X1 g15451(.A (n_3084), .B (n_3382), .Y (n_5641));
NOR2X1 g15455(.A (n_2774), .B (n_3380), .Y (n_6081));
NOR2X1 g15456(.A (n_3381), .B (n_3252), .Y (n_3494));
NAND2X1 g15465(.A (n_7648), .B (n_7649), .Y (n_3493));
NAND2X1 g15469(.A (n_3355), .B (n_3354), .Y (n_3492));
NAND2X1 g15479(.A (n_3345), .B (n_3190), .Y (n_3491));
NOR2X1 g15501(.A (n_3267), .B (n_3361), .Y (n_3487));
NOR2X1 g15504(.A (n_3262), .B (n_3352), .Y (n_7784));
AOI22X1 g15515(.A0 (n_3151), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_35), .Y (n_3485));
AOI22X1 g15526(.A0 (n_3311), .A1 (n_1260), .B0 (n_3550), .B1(FP_R_55), .Y (n_3483));
NOR2X1 g15565(.A (n_3002), .B (n_3337), .Y (n_3481));
NOR2X1 g15567(.A (n_3319), .B (n_3235), .Y (n_3480));
NAND2X1 g15585(.A (n_3048), .B (n_3336), .Y (n_3479));
NOR2X1 g15587(.A (n_3178), .B (n_3338), .Y (n_3478));
AND2X1 g15617(.A (n_2991), .B (n_3329), .Y (n_5667));
NOR2X1 g15625(.A (n_3317), .B (n_3026), .Y (n_7785));
NOR2X1 g15643(.A (n_3316), .B (n_3325), .Y (n_3473));
NOR2X1 g15644(.A (n_3201), .B (n_3324), .Y (n_3472));
NOR2X1 g15647(.A (n_3315), .B (n_3322), .Y (n_3471));
MX2X1 g16053(.A (L_67), .B (FP_R_36), .S0 (n_7846), .Y (n_3468));
MX2X1 g16054(.A (L_84), .B (FP_R_53), .S0 (n_7846), .Y (n_3467));
MX2X1 g16055(.A (L_76), .B (FP_R_45), .S0 (n_7846), .Y (n_3466));
MX2X1 g16056(.A (L_68), .B (FP_R_37), .S0 (n_7846), .Y (n_3465));
AOI21X1 g16058(.A0 (n_99), .A1 (n_7846), .B0 (n_3309), .Y (n_3463));
MX2X1 g16059(.A (L_69), .B (FP_R_38), .S0 (n_7846), .Y (n_3462));
MX2X1 g16063(.A (L), .B (FP_R_32), .S0 (n_7846), .Y (n_3460));
MX2X1 g16064(.A (L_70), .B (FP_R_39), .S0 (n_7846), .Y (n_3459));
MX2X1 g16066(.A (L_89), .B (FP_R_58), .S0 (n_7846), .Y (n_3458));
MX2X1 g16070(.A (L_90), .B (FP_R_59), .S0 (n_7846), .Y (n_3457));
MX2X1 g16071(.A (L_87), .B (FP_R_56), .S0 (n_7846), .Y (n_3456));
MX2X1 g16072(.A (L_82), .B (FP_R_51), .S0 (n_7846), .Y (n_3455));
MX2X1 g16073(.A (L_74), .B (FP_R_43), .S0 (n_7846), .Y (n_3454));
MX2X1 g16643(.A (L_79), .B (FP_R_48), .S0 (n_7846), .Y (n_3453));
MX2X1 g16644(.A (L_73), .B (FP_R_42), .S0 (n_7846), .Y (n_3451));
NOR2X1 g15480(.A (n_3287), .B (n_3282), .Y (n_3446));
NOR2X1 g15481(.A (n_5898), .B (n_5897), .Y (n_3445));
NOR2X1 g15482(.A (n_3273), .B (n_3272), .Y (n_3444));
NOR2X1 g15489(.A (n_7675), .B (n_7674), .Y (n_5591));
MX2X1 g17140(.A (L_88), .B (FP_R_57), .S0 (n_7846), .Y (n_3442));
MX2X1 g17142(.A (L_94), .B (FP_R_63), .S0 (n_7846), .Y (n_3440));
NOR2X1 g15500(.A (n_3269), .B (n_3268), .Y (n_3436));
NOR2X1 g15502(.A (n_2782), .B (n_3266), .Y (n_7790));
NOR2X1 g15507(.A (n_3258), .B (n_3257), .Y (n_3432));
AND2X1 g15540(.A (n_3185), .B (n_3247), .Y (n_3430));
AND2X1 g15541(.A (n_3144), .B (n_3160), .Y (n_3429));
AOI21X1 g15542(.A0 (n_2369), .A1 (n_170), .B0 (n_3183), .Y (n_3428));
NAND3X1 g15548(.A (n_3070), .B (n_2642), .C (n_3133), .Y (n_3426));
NAND2X1 g15557(.A (n_3180), .B (n_3240), .Y (n_3425));
AND2X1 g15564(.A (n_3176), .B (n_3238), .Y (n_3423));
NOR2X1 g15569(.A (n_3011), .B (n_3233), .Y (n_3422));
NAND2X1 g15578(.A (n_7676), .B (n_7677), .Y (n_3421));
AND2X1 g15581(.A (n_3177), .B (n_2767), .Y (n_3420));
NAND3X1 g15582(.A (n_7891), .B (n_3149), .C (n_7892), .Y (n_3419));
NAND2X1 g15584(.A (n_3208), .B (n_2738), .Y (n_3418));
NAND2X1 g15590(.A (n_2998), .B (n_3226), .Y (n_3417));
NOR2X1 g15591(.A (n_3174), .B (n_3223), .Y (n_3416));
NOR2X1 g15599(.A (n_3173), .B (n_3221), .Y (n_3414));
AND2X1 g15612(.A (n_3057), .B (n_3228), .Y (n_3411));
NAND2X1 g15620(.A (n_3171), .B (n_3028), .Y (n_3410));
NAND3X1 g15635(.A (n_3203), .B (n_1798), .C (n_2582), .Y (n_3406));
NOR2X1 g15639(.A (n_3167), .B (n_2985), .Y (n_3405));
NAND2X1 g15642(.A (n_2988), .B (n_3202), .Y (n_3404));
NOR2X1 g15648(.A (n_3198), .B (n_3197), .Y (n_3403));
NOR2X1 g15669(.A (n_3162), .B (n_3191), .Y (n_5610));
AND2X1 g15670(.A (n_3161), .B (n_2833), .Y (n_3401));
NAND3X1 g15671(.A (n_3188), .B (n_2206), .C (n_2570), .Y (n_3400));
NAND2X1 g15675(.A (n_2644), .B (n_3158), .Y (n_3399));
AOI21X1 g15688(.A0 (n_2007), .A1 (n_2490), .B0 (n_3305), .Y (n_3398));
AND2X1 g15692(.A (n_3304), .B (n_2893), .Y (n_3397));
NAND2X1 g15838(.A (n_2841), .B (n_3303), .Y (n_3395));
NAND2X1 g15840(.A (n_2903), .B (n_3302), .Y (n_3394));
AND2X1 g15936(.A (n_3301), .B (n_2805), .Y (n_3393));
AND2X1 g15939(.A (n_1842), .B (n_3308), .Y (n_3392));
MX2X1 g16057(.A (L_85), .B (FP_R_54), .S0 (n_7846), .Y (n_3391));
MX2X1 g16067(.A (L_81), .B (FP_R_50), .S0 (n_7846), .Y (n_3390));
MX2X1 g17141(.A (L_93), .B (FP_R_62), .S0 (n_7846), .Y (n_3387));
NAND2X1 g15472(.A (n_2269), .B (n_3085), .Y (n_3383));
NAND3X1 g15473(.A (n_2291), .B (n_2892), .C (n_1705), .Y (n_3382));
NAND2X1 g15475(.A (n_3076), .B (n_2651), .Y (n_3381));
NAND3X1 g15476(.A (n_1860), .B (n_1888), .C (n_2764), .Y (n_3380));
NAND3X1 g15477(.A (n_3081), .B (n_2573), .C (n_2103), .Y (n_3379));
NAND2X1 g15478(.A (n_2770), .B (n_3078), .Y (n_3378));
MX2X1 g17139(.A (L_83), .B (FP_R_52), .S0 (n_7846), .Y (n_3377));
NAND3X1 g15554(.A (n_3065), .B (n_2223), .C (n_2595), .Y (n_3372));
NOR2X1 g15579(.A (n_3056), .B (n_3021), .Y (n_6084));
NOR2X1 g15589(.A (n_3060), .B (n_3061), .Y (n_5592));
NAND3X1 g15601(.A (n_2720), .B (n_2960), .C (n_2608), .Y (n_3361));
NOR2X1 g15602(.A (n_2994), .B (n_3040), .Y (n_5596));
NOR2X1 g15607(.A (n_2993), .B (n_3030), .Y (n_6082));
NAND2X1 g15608(.A (n_2716), .B (n_3036), .Y (n_3358));
NAND2X1 g15610(.A (n_2713), .B (n_3035), .Y (n_3357));
NAND2X1 g15613(.A (n_2992), .B (n_3033), .Y (n_3356));
AOI21X1 g15622(.A0 (n_1995), .A1 (n_2931), .B0 (n_2980), .Y (n_3355));
AOI21X1 g15623(.A0 (n_2792), .A1 (n_3159), .B0 (n_2979), .Y (n_3354));
AOI21X1 g15624(.A0 (n_2944), .A1 (n_177), .B0 (n_2982), .Y (n_7648));
NAND3X1 g15627(.A (n_2704), .B (n_2955), .C (n_2627), .Y (n_3352));
NOR2X1 g15628(.A (n_2989), .B (n_2670), .Y (n_3351));
NOR2X1 g15641(.A (n_2655), .B (n_3016), .Y (n_3349));
NOR2X1 g15663(.A (n_3008), .B (n_3007), .Y (n_3346));
AOI21X1 g15677(.A0 (n_7684), .A1 (n_2613), .B0 (n_3147), .Y (n_3345));
AND2X1 g15693(.A (n_2812), .B (n_3135), .Y (n_3344));
AOI21X1 g15730(.A0 (n_2801), .A1 (n_177), .B0 (n_2921), .Y (n_3342));
AOI21X1 g15734(.A0 (n_1979), .A1 (n_3194), .B0 (n_3142), .Y (n_3341));
NAND2X1 g15740(.A (n_3129), .B (n_3115), .Y (n_3340));
NAND2X1 g15744(.A (n_2925), .B (n_3143), .Y (n_3339));
NAND2X1 g15758(.A (n_2874), .B (n_3132), .Y (n_3338));
NAND2X1 g15767(.A (n_3140), .B (n_2455), .Y (n_3337));
AOI21X1 g15773(.A0 (n_2799), .A1 (n_7301), .B0 (n_2891), .Y (n_3336));
AOI21X1 g15833(.A0 (n_2798), .A1 (n_2842), .B0 (n_2417), .Y (n_7521));
AOI21X1 g15839(.A0 (n_1947), .A1 (n_170), .B0 (n_3120), .Y (n_3329));
NAND2X1 g15881(.A (n_2819), .B (n_3109), .Y (n_3325));
NAND2X1 g15885(.A (n_3107), .B (n_2818), .Y (n_3324));
OR2X1 g15891(.A (n_3105), .B (n_2310), .Y (n_3323));
OR2X1 g15892(.A (n_2390), .B (n_3101), .Y (n_3322));
AOI21X1 g15951(.A0 (n_1855), .A1 (n_3153), .B0 (n_3130), .Y (n_3321));
NAND2X1 g15955(.A (n_2234), .B (n_3116), .Y (n_3320));
NAND2X1 g15958(.A (n_1833), .B (n_3128), .Y (n_3319));
NAND2X1 g15977(.A (n_2959), .B (n_3122), .Y (n_3318));
NAND2X1 g15981(.A (n_6017), .B (n_6018), .Y (n_3317));
NAND2X1 g15992(.A (n_2578), .B (n_3110), .Y (n_3316));
NAND2X1 g15996(.A (n_2213), .B (n_3103), .Y (n_3315));
INVX1 g16046(.A (n_3152), .Y (n_3314));
MX2X1 g16052(.A (L_75), .B (FP_R_44), .S0 (n_7846), .Y (n_3313));
MX2X1 g16060(.A (L_86), .B (FP_R_55), .S0 (n_7846), .Y (n_3311));
AOI22X1 g16026(.A0 (n_2990), .A1 (n_3153), .B0 (n_3154), .B1(n_2624), .Y (n_3310));
NOR2X1 g16122(.A (L_77), .B (n_7846), .Y (n_3309));
INVX1 g16197(.A (n_3145), .Y (n_3308));
AOI21X1 g16340(.A0 (n_2340), .A1 (n_2034), .B0 (n_275), .Y (n_3305));
NAND2X1 g16344(.A (n_2802), .B (n_177), .Y (n_3304));
NAND2X1 g16514(.A (n_2788), .B (n_3189), .Y (n_3303));
NAND2X1 g16516(.A (n_2795), .B (n_2842), .Y (n_3302));
NAND2X1 g16525(.A (n_2797), .B (n_3134), .Y (n_3301));
CLKBUFX1 gbuf_d_65(.A(desOut[53]), .Y(d_out_65));
CLKBUFX1 gbuf_q_65(.A(q_in_65), .Y(L_80));
CLKBUFX1 gbuf_d_66(.A(desOut[51]), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(L_72));
CLKBUFX1 gbuf_d_67(.A(desOut[41]), .Y(d_out_67));
CLKBUFX1 gbuf_q_67(.A(q_in_67), .Y(L_65));
CLKBUFX1 gbuf_d_68(.A(desOut[19]), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(L_76));
CLKBUFX1 gbuf_d_69(.A(desOut[21]), .Y(d_out_69));
CLKBUFX1 gbuf_q_69(.A(q_in_69), .Y(L_84));
CLKBUFX1 gbuf_d_70(.A(desOut[17]), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(L_68));
CLKBUFX1 gbuf_d_71(.A(desOut[25]), .Y(d_out_71));
CLKBUFX1 gbuf_q_71(.A(q_in_71), .Y(L_67));
CLKBUFX1 gbuf_d_72(.A(desOut[3]), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(L_78));
CLKBUFX1 gbuf_d_73(.A(desOut[23]), .Y(d_out_73));
CLKBUFX1 gbuf_q_73(.A(q_in_73), .Y(L_92));
CLKBUFX1 gbuf_d_74(.A(desOut[59]), .Y(d_out_74));
CLKBUFX1 gbuf_q_74(.A(q_in_74), .Y(L_71));
CLKBUFX1 gbuf_d_75(.A(desOut[49]), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(L_64));
NAND2X1 g15543(.A (n_2263), .B (n_2761), .Y (n_3287));
NAND2X1 g15553(.A (n_2672), .B (n_2282), .Y (n_3285));
NAND3X1 g15555(.A (n_2759), .B (n_1822), .C (n_2196), .Y (n_3284));
NAND2X1 g15559(.A (n_2705), .B (n_2734), .Y (n_3282));
NAND3X1 g15562(.A (n_2711), .B (n_2636), .C (n_2403), .Y (n_3281));
NAND3X1 g15563(.A (n_2753), .B (n_2237), .C (n_1832), .Y (n_3280));
NAND2X1 g15575(.A (n_5668), .B (n_5669), .Y (n_5897));
NAND2X1 g15576(.A (n_2667), .B (n_1883), .Y (n_3276));
NAND3X1 g15577(.A (n_2742), .B (n_2612), .C (n_1824), .Y (n_3275));
NAND2X1 g15580(.A (n_2709), .B (n_2740), .Y (n_5898));
NAND2X1 g15583(.A (n_5694), .B (n_5695), .Y (n_3273));
NAND2X1 g15586(.A (n_6091), .B (n_6092), .Y (n_3272));
NAND2X1 g15594(.A (n_2665), .B (n_2729), .Y (n_3271));
NAND2X1 g15595(.A (n_2728), .B (n_2727), .Y (n_3270));
NAND3X1 g15597(.A (n_2723), .B (n_2610), .C (n_2437), .Y (n_3269));
NAND3X1 g15598(.A (n_2721), .B (n_2607), .C (n_2605), .Y (n_3268));
NAND2X1 g15600(.A (n_2664), .B (n_2725), .Y (n_3267));
NAND3X1 g15604(.A (n_5968), .B (n_5969), .C (n_1812), .Y (n_3266));
NAND2X1 g15618(.A (n_2737), .B (n_2765), .Y (n_7674));
NAND2X1 g15621(.A (n_7801), .B (n_7802), .Y (n_7675));
NAND2X1 g15626(.A (n_5970), .B (n_5971), .Y (n_3262));
NAND2X1 g15645(.A (n_2654), .B (n_2693), .Y (n_3258));
NAND3X1 g15646(.A (n_2689), .B (n_1794), .C (n_1792), .Y (n_3257));
NAND2X1 g15651(.A (n_2271), .B (n_2688), .Y (n_3255));
NOR2X1 g15653(.A (n_2256), .B (n_2685), .Y (n_5642));
NAND2X1 g15661(.A (n_2650), .B (n_2674), .Y (n_3252));
NAND2X1 g15666(.A (n_2283), .B (n_2673), .Y (n_3251));
AOI21X1 g15687(.A0 (n_2317), .A1 (n_3194), .B0 (n_2201), .Y (n_3248));
AOI21X1 g15690(.A0 (n_2004), .A1 (n_2744), .B0 (n_2896), .Y (n_3247));
AOI21X1 g15698(.A0 (n_1923), .A1 (n_2735), .B0 (n_2871), .Y (n_3245));
AOI21X1 g15700(.A0 (n_2318), .A1 (n_2686), .B0 (n_1754), .Y (n_3244));
NAND2X1 g15701(.A (n_2932), .B (n_2491), .Y (n_3243));
AOI21X1 g15721(.A0 (n_2306), .A1 (n_7341), .B0 (n_2383), .Y (n_3240));
AOI21X1 g15729(.A0 (n_1969), .A1 (n_2490), .B0 (n_2883), .Y (n_3238));
OR2X1 g15732(.A (n_2476), .B (n_2881), .Y (n_3235));
AND2X1 g15733(.A (n_2878), .B (n_2927), .Y (n_3234));
NAND2X1 g15745(.A (n_2876), .B (n_2469), .Y (n_3233));
AOI21X1 g15747(.A0 (n_1602), .A1 (n_3054), .B0 (n_2930), .Y (n_3232));
AOI21X1 g15760(.A0 (n_2355), .A1 (n_2931), .B0 (n_2834), .Y (n_7676));
AND2X1 g15764(.A (n_2829), .B (n_2843), .Y (n_3229));
AOI21X1 g15766(.A0 (n_2359), .A1 (n_3153), .B0 (n_2868), .Y (n_3228));
AND2X1 g15774(.A (n_2827), .B (n_2538), .Y (n_3227));
AOI21X1 g15781(.A0 (n_2322), .A1 (n_2744), .B0 (n_2095), .Y (n_3226));
NAND2X1 g15786(.A (n_2917), .B (n_2859), .Y (n_3223));
NAND2X1 g15793(.A (n_2914), .B (n_2857), .Y (n_3221));
AOI21X1 g15834(.A0 (n_2326), .A1 (n_2931), .B0 (n_2905), .Y (n_3211));
AND2X1 g15843(.A (n_2902), .B (n_2832), .Y (n_3210));
AND2X1 g15844(.A (n_2872), .B (n_2918), .Y (n_3209));
AOI21X1 g15846(.A0 (n_2344), .A1 (n_3044), .B0 (n_2936), .Y (n_3208));
NAND2X1 g15856(.A (n_2826), .B (n_2459), .Y (n_3207));
AOI21X1 g15868(.A0 (n_2316), .A1 (n_2402), .B0 (n_2377), .Y (n_3204));
AOI21X1 g15871(.A0 (n_2314), .A1 (n_7341), .B0 (n_2395), .Y (n_3203));
AOI21X1 g15880(.A0 (n_1954), .A1 (n_3121), .B0 (n_2822), .Y (n_3202));
NAND2X1 g15883(.A (n_2540), .B (n_2900), .Y (n_3201));
AOI21X1 g15884(.A0 (n_2312), .A1 (n_3106), .B0 (n_2040), .Y (n_3200));
AOI21X1 g15886(.A0 (n_1914), .A1 (n_170), .B0 (n_2809), .Y (n_3199));
OR2X1 g15893(.A (n_2388), .B (n_2815), .Y (n_3198));
OR2X1 g15894(.A (n_2158), .B (n_2899), .Y (n_3197));
NAND2X1 g15917(.A (n_2150), .B (n_2860), .Y (n_3196));
AOI21X1 g15921(.A0 (n_2305), .A1 (n_3194), .B0 (n_2014), .Y (n_3195));
AOI21X1 g15926(.A0 (n_2361), .A1 (n_2402), .B0 (n_2941), .Y (n_3193));
AOI21X1 g15932(.A0 (n_2261), .A1 (n_2624), .B0 (n_2013), .Y (n_3192));
OR2X1 g15933(.A (n_2898), .B (n_2375), .Y (n_3191));
AOI21X1 g15934(.A0 (n_2339), .A1 (n_3189), .B0 (n_2011), .Y (n_3190));
AOI21X1 g15935(.A0 (n_1482), .A1 (n_7341), .B0 (n_2807), .Y (n_3188));
AOI21X1 g15937(.A0 (n_2956), .A1 (n_2668), .B0 (n_2889), .Y (n_3186));
AOI21X1 g15938(.A0 (n_1786), .A1 (n_2624), .B0 (n_2897), .Y (n_3185));
AOI21X1 g15940(.A0 (n_2806), .A1 (n_3146), .B0 (n_2182), .Y (n_3183));
NAND2X1 g15942(.A (n_2965), .B (n_2828), .Y (n_3181));
AOI21X1 g15948(.A0 (n_2649), .A1 (n_3179), .B0 (n_2831), .Y (n_3180));
NAND2X1 g15956(.A (n_2615), .B (n_2923), .Y (n_3178));
AOI21X1 g15960(.A0 (n_3170), .A1 (n_2613), .B0 (n_2493), .Y (n_3177));
AOI21X1 g15962(.A0 (n_2639), .A1 (n_2668), .B0 (n_2867), .Y (n_3176));
NAND2X1 g15965(.A (n_2962), .B (n_2862), .Y (n_3174));
NAND2X1 g15969(.A (n_2609), .B (n_2915), .Y (n_3173));
AOI21X1 g15979(.A0 (n_3170), .A1 (n_2668), .B0 (n_2840), .Y (n_3171));
NAND2X1 g15983(.A (n_2953), .B (n_2399), .Y (n_3168));
NAND2X1 g15988(.A (n_2580), .B (n_2817), .Y (n_3167));
AOI21X1 g15995(.A0 (n_2238), .A1 (n_2613), .B0 (n_2886), .Y (n_3166));
AOI21X1 g15997(.A0 (n_2671), .A1 (n_3153), .B0 (n_2814), .Y (n_3164));
NAND2X1 g16009(.A (n_2242), .B (n_2810), .Y (n_3162));
INVX1 g16010(.A (n_2984), .Y (n_3161));
NAND2X1 g16012(.A (n_2966), .B (n_3159), .Y (n_3160));
CLKBUFX1 gbuf_d_76(.A(desOut[3]), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(FP_R_15));
NAND2X1 g16021(.A (n_2943), .B (n_7301), .Y (n_3158));
CLKBUFX1 gbuf_d_77(.A(desOut[23]), .Y(d_out_77));
CLKBUFX1 gbuf_q_77(.A(q_in_77), .Y(FP_R_29));
CLKBUFX1 gbuf_d_78(.A(desOut[59]), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(FP_R_8));
CLKBUFX1 gbuf_d_79(.A(desOut[51]), .Y(d_out_79));
CLKBUFX1 gbuf_q_79(.A(q_in_79), .Y(FP_R_9));
CLKBUFX1 gbuf_d_80(.A(desOut[41]), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(FP_R_2));
CLKBUFX1 gbuf_d_81(.A(desOut[53]), .Y(d_out_81));
CLKBUFX1 gbuf_q_81(.A(q_in_81), .Y(FP_R_17));
CLKBUFX1 gbuf_d_82(.A(desOut[25]), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(FP_R_4));
CLKBUFX1 gbuf_d_83(.A(desOut[17]), .Y(d_out_83));
CLKBUFX1 gbuf_q_83(.A(q_in_83), .Y(FP_R_5));
CLKBUFX1 gbuf_d_84(.A(desOut[21]), .Y(d_out_84));
CLKBUFX1 gbuf_q_84(.A(q_in_84), .Y(FP_R_21));
CLKBUFX1 gbuf_d_85(.A(desOut[19]), .Y(d_out_85));
CLKBUFX1 gbuf_q_85(.A(q_in_85), .Y(FP_R_13));
CLKBUFX1 gbuf_d_86(.A(desOut[49]), .Y(d_out_86));
CLKBUFX1 gbuf_q_86(.A(q_in_86), .Y(FP_R_1));
AOI21X1 g16043(.A0 (n_3154), .A1 (n_3153), .B0 (n_2957), .Y (n_3155));
NAND2X1 g16047(.A (n_2950), .B (n_2947), .Y (n_3152));
MX2X1 g16050(.A (L_66), .B (FP_R_35), .S0 (n_7846), .Y (n_3151));
CLKBUFX1 gbuf_d_87(.A(desOut[57]), .Y(d_out_87));
CLKBUFX1 gbuf_q_87(.A(q_in_87), .Y(FP_R));
NAND2X1 g16135(.A (n_7683), .B (n_2668), .Y (n_3149));
AOI21X1 g16025(.A0 (n_2838), .A1 (n_3146), .B0 (n_329), .Y (n_3147));
AOI21X1 g16198(.A0 (n_1942), .A1 (n_2039), .B0 (n_235), .Y (n_3145));
INVX1 g16200(.A (n_2939), .Y (n_3144));
NAND2X1 g16208(.A (n_2351), .B (n_2928), .Y (n_3143));
AOI21X1 g16225(.A0 (n_2396), .A1 (n_1619), .B0 (n_7437), .Y (n_3142));
NAND2X1 g16228(.A (n_2349), .B (n_189), .Y (n_3140));
NAND2X1 g16266(.A (n_2364), .B (n_2974), .Y (n_3139));
INVX1 g16279(.A (n_2908), .Y (n_3138));
NAND2X1 g16299(.A (n_2362), .B (n_2539), .Y (n_6017));
NAND2X1 g16347(.A (n_2371), .B (n_3134), .Y (n_3135));
NAND2X1 g16353(.A (n_2365), .B (n_170), .Y (n_3133));
NAND2X1 g16383(.A (n_2345), .B (n_3189), .Y (n_3132));
AOI21X1 g16387(.A0 (n_1312), .A1 (n_7442), .B0 (n_2440), .Y (n_3130));
NAND2X1 g16396(.A (n_2357), .B (n_3044), .Y (n_3129));
NAND2X1 g16422(.A (n_2348), .B (n_2842), .Y (n_3128));
NAND2X1 g16478(.A (n_2337), .B (n_2666), .Y (n_3126));
NAND2X1 g16479(.A (n_2315), .B (n_170), .Y (n_3125));
NAND2X1 g16493(.A (n_2331), .B (n_7301), .Y (n_3123));
NAND2X1 g16509(.A (n_2324), .B (n_3121), .Y (n_3122));
AOI21X1 g16515(.A0 (n_1942), .A1 (n_1616), .B0 (n_2488), .Y (n_3120));
AOI21X1 g16534(.A0 (n_2396), .A1 (n_3117), .B0 (n_297), .Y (n_3119));
NAND2X1 g16539(.A (n_2341), .B (n_2404), .Y (n_3116));
NAND2X1 g16549(.A (n_2353), .B (n_7301), .Y (n_3115));
NAND2X1 g16556(.A (n_2367), .B (n_177), .Y (n_3114));
NAND2X1 g16558(.A (n_2304), .B (n_2735), .Y (n_3112));
NAND2X1 g16575(.A (n_2313), .B (n_2686), .Y (n_3110));
NAND2X1 g16577(.A (n_2325), .B (n_7301), .Y (n_3109));
NAND2X1 g16578(.A (n_2354), .B (n_3106), .Y (n_3107));
AOI21X1 g16584(.A0 (n_2105), .A1 (n_3104), .B0 (n_2440), .Y (n_3105));
NAND2X1 g16586(.A (n_2278), .B (n_177), .Y (n_3103));
AND2X1 g16589(.A (n_2307), .B (n_3159), .Y (n_3101));
CLKBUFX1 gbuf_d_88(.A(desOut[63]), .Y(d_out_88));
CLKBUFX1 gbuf_q_88(.A(q_in_88), .Y(L_87));
CLKBUFX1 gbuf_d_89(.A(desOut[9]), .Y(d_out_89));
CLKBUFX1 gbuf_q_89(.A(q_in_89), .Y(L_69));
CLKBUFX1 gbuf_d_90(.A(desOut[57]), .Y(d_out_90));
CLKBUFX1 gbuf_q_90(.A(q_in_90), .Y(L));
CLKBUFX1 gbuf_d_91(.A(desOut[1]), .Y(d_out_91));
CLKBUFX1 gbuf_q_91(.A(q_in_91), .Y(L_70));
CLKBUFX1 gbuf_d_92(.A(desOut[37]), .Y(d_out_92));
CLKBUFX1 gbuf_q_92(.A(q_in_92), .Y(L_82));
CLKBUFX1 gbuf_d_93(.A(desOut[47]), .Y(d_out_93));
CLKBUFX1 gbuf_q_93(.A(q_in_93), .Y(L_89));
CLKBUFX1 gbuf_d_94(.A(desOut[39]), .Y(d_out_94));
CLKBUFX1 gbuf_q_94(.A(q_in_94), .Y(L_90));
CLKBUFX1 gbuf_d_95(.A(desOut[35]), .Y(d_out_95));
CLKBUFX1 gbuf_q_95(.A(q_in_95), .Y(L_74));
NAND3X1 g15468(.A (n_1876), .B (n_1878), .C (n_2072), .Y (n_3093));
CLKBUFX1 gbuf_d_96(.A(desOut[61]), .Y(d_out_96));
CLKBUFX1 gbuf_q_96(.A(q_in_96), .Y(L_79));
CLKBUFX1 gbuf_d_97(.A(desOut[43]), .Y(d_out_97));
CLKBUFX1 gbuf_q_97(.A(q_in_97), .Y(L_73));
NAND2X1 g15573(.A (n_2547), .B (n_1849), .Y (n_3090));
CLKBUFX1 gbuf_d_98(.A(desOut[7]), .Y(d_out_98));
CLKBUFX1 gbuf_q_98(.A(q_in_98), .Y(L_94));
CLKBUFX1 gbuf_d_99(.A(desOut[55]), .Y(d_out_99));
CLKBUFX1 gbuf_q_99(.A(q_in_99), .Y(L_88));
AOI21X1 g15652(.A0 (n_2211), .A1 (n_7344), .B0 (n_1398), .Y (n_3085));
NAND3X1 g15654(.A (n_7898), .B (n_7899), .C (n_1416), .Y (n_3084));
AOI21X1 g15662(.A0 (n_1732), .A1 (n_6805), .B0 (n_2252), .Y (n_3081));
NOR2X1 g15664(.A (n_2254), .B (n_2266), .Y (n_3080));
NOR2X1 g15665(.A (n_2265), .B (n_2264), .Y (n_6102));
NOR2X1 g15668(.A (n_1778), .B (n_2246), .Y (n_3078));
AOI21X1 g15672(.A0 (n_1133), .A1 (n_7341), .B0 (n_2249), .Y (n_5684));
AOI21X1 g15676(.A0 (n_2619), .A1 (n_2653), .B0 (n_2253), .Y (n_3076));
AOI21X1 g15689(.A0 (n_1941), .A1 (n_2842), .B0 (n_2568), .Y (n_3074));
AOI21X1 g15704(.A0 (n_1940), .A1 (n_2735), .B0 (n_2454), .Y (n_3071));
NOR2X1 g15706(.A (n_2198), .B (n_2489), .Y (n_3070));
NAND2X1 g15709(.A (n_2172), .B (n_2483), .Y (n_3068));
NAND2X1 g15711(.A (n_2482), .B (n_2565), .Y (n_3067));
NOR2X1 g15714(.A (n_2564), .B (n_2130), .Y (n_3065));
NAND2X1 g15739(.A (n_2460), .B (n_2411), .Y (n_3061));
NAND2X1 g15741(.A (n_2545), .B (n_2381), .Y (n_3060));
NAND2X1 g15749(.A (n_2110), .B (n_2552), .Y (n_3059));
NAND2X1 g15750(.A (n_2109), .B (n_2468), .Y (n_3058));
AOI21X1 g15752(.A0 (n_1939), .A1 (n_3121), .B0 (n_2461), .Y (n_3057));
NAND2X1 g15753(.A (n_7798), .B (n_7799), .Y (n_3056));
NAND2X1 g15759(.A (n_2135), .B (n_2484), .Y (n_3053));
AOI21X1 g15761(.A0 (n_1949), .A1 (n_2171), .B0 (n_1848), .Y (n_7677));
AOI21X1 g15768(.A0 (n_1579), .A1 (n_3054), .B0 (n_2457), .Y (n_3051));
AOI21X1 g15770(.A0 (n_1692), .A1 (n_3049), .B0 (n_2551), .Y (n_3050));
NOR2X1 g15772(.A (n_2049), .B (n_2406), .Y (n_3048));
NAND2X1 g15782(.A (n_2535), .B (n_2536), .Y (n_3047));
AOI21X1 g15789(.A0 (n_1929), .A1 (n_3044), .B0 (n_2531), .Y (n_3045));
NAND2X1 g15795(.A (n_2438), .B (n_2430), .Y (n_3043));
AOI21X1 g15800(.A0 (n_1977), .A1 (n_3049), .B0 (n_1734), .Y (n_3042));
AOI21X1 g15801(.A0 (n_1566), .A1 (n_7301), .B0 (n_2434), .Y (n_3041));
NAND2X1 g15802(.A (n_2530), .B (n_2433), .Y (n_3040));
AOI21X1 g15803(.A0 (n_1956), .A1 (n_2695), .B0 (n_2431), .Y (n_3039));
AOI21X1 g15806(.A0 (n_1955), .A1 (n_204), .B0 (n_2429), .Y (n_7791));
AOI21X1 g15816(.A0 (n_1952), .A1 (n_7301), .B0 (n_2175), .Y (n_3036));
AOI21X1 g15819(.A0 (n_1510), .A1 (n_2856), .B0 (n_2523), .Y (n_3035));
AOI21X1 g15827(.A0 (n_1497), .A1 (n_170), .B0 (n_2522), .Y (n_3033));
NAND2X1 g15835(.A (n_1769), .B (n_2405), .Y (n_3030));
OR2X1 g15836(.A (n_2409), .B (n_2407), .Y (n_3029));
AOI21X1 g15841(.A0 (n_1931), .A1 (n_7301), .B0 (n_2517), .Y (n_3028));
AOI21X1 g15842(.A0 (n_1975), .A1 (n_7301), .B0 (n_2225), .Y (n_3027));
NAND2X1 g15849(.A (n_2510), .B (n_2400), .Y (n_3026));
AOI21X1 g15854(.A0 (n_2001), .A1 (n_2863), .B0 (n_1710), .Y (n_7892));
NAND2X1 g15863(.A (n_2463), .B (n_2466), .Y (n_3021));
AOI21X1 g15864(.A0 (n_1429), .A1 (n_2719), .B0 (n_2397), .Y (n_7886));
NAND2X1 g15875(.A (n_2393), .B (n_2494), .Y (n_3019));
NAND2X1 g15882(.A (n_2502), .B (n_2501), .Y (n_3016));
AOI21X1 g15890(.A0 (n_1963), .A1 (n_177), .B0 (n_2032), .Y (n_3015));
NAND2X1 g15895(.A (n_2387), .B (n_2386), .Y (n_3014));
NAND2X1 g15896(.A (n_2385), .B (n_1763), .Y (n_3013));
NAND2X1 g15899(.A (n_2498), .B (n_2193), .Y (n_3011));
NAND2X1 g15901(.A (n_2465), .B (n_2549), .Y (n_3010));
NAND2X1 g15911(.A (n_2496), .B (n_2379), .Y (n_3009));
NAND2X1 g15922(.A (n_2514), .B (n_2057), .Y (n_3008));
NAND2X1 g15924(.A (n_2378), .B (n_2537), .Y (n_3007));
AOI21X1 g15925(.A0 (n_1685), .A1 (n_2744), .B0 (n_2475), .Y (n_3006));
NAND2X1 g15952(.A (n_2625), .B (n_2472), .Y (n_3002));
NAND2X1 g15954(.A (n_2623), .B (n_1729), .Y (n_3000));
NAND2X1 g15961(.A (n_2239), .B (n_2413), .Y (n_2999));
AOI21X1 g15963(.A0 (n_2257), .A1 (n_2624), .B0 (n_2534), .Y (n_2998));
NAND2X1 g15964(.A (n_2229), .B (n_2449), .Y (n_2997));
NAND2X1 g15968(.A (n_1816), .B (n_2439), .Y (n_2995));
NAND2X1 g15971(.A (n_2603), .B (n_2104), .Y (n_2994));
NAND2X1 g15973(.A (n_2601), .B (n_2520), .Y (n_2993));
AOI21X1 g15974(.A0 (n_2626), .A1 (n_3153), .B0 (n_2419), .Y (n_2992));
AOI21X1 g15978(.A0 (n_2990), .A1 (n_2624), .B0 (n_2063), .Y (n_2991));
NAND2X1 g15985(.A (n_2222), .B (n_2451), .Y (n_2989));
AOI21X1 g15991(.A0 (n_2660), .A1 (n_2624), .B0 (n_2504), .Y (n_2988));
AOI21X1 g15994(.A0 (n_2594), .A1 (n_2624), .B0 (n_2500), .Y (n_2987));
NAND2X1 g15999(.A (n_1828), .B (n_2555), .Y (n_2986));
NAND2X1 g16000(.A (n_2576), .B (n_2435), .Y (n_2985));
AOI21X1 g16011(.A0 (n_2981), .A1 (n_2830), .B0 (n_235), .Y (n_2984));
AOI21X1 g16014(.A0 (n_1753), .A1 (n_2981), .B0 (n_192), .Y (n_2983));
AOI21X1 g16015(.A0 (n_2935), .A1 (n_2981), .B0 (n_2042), .Y (n_2982));
AOI21X1 g16016(.A0 (n_3146), .A1 (n_2506), .B0 (n_2042), .Y (n_2980));
AOI21X1 g16017(.A0 (n_2981), .A1 (n_1310), .B0 (n_275), .Y (n_2979));
CLKBUFX1 gbuf_d_100(.A(desOut[9]), .Y(d_out_100));
CLKBUFX1 gbuf_q_100(.A(q_in_100), .Y(FP_R_6));
CLKBUFX1 gbuf_d_101(.A(desOut[43]), .Y(d_out_101));
CLKBUFX1 gbuf_q_101(.A(q_in_101), .Y(FP_R_10));
CLKBUFX1 gbuf_d_102(.A(desOut[35]), .Y(d_out_102));
CLKBUFX1 gbuf_q_102(.A(q_in_102), .Y(FP_R_11));
CLKBUFX1 gbuf_d_103(.A(desOut[63]), .Y(d_out_103));
CLKBUFX1 gbuf_q_103(.A(q_in_103), .Y(FP_R_24));
CLKBUFX1 gbuf_d_104(.A(desOut[47]), .Y(d_out_104));
CLKBUFX1 gbuf_q_104(.A(q_in_104), .Y(FP_R_26));
CLKBUFX1 gbuf_d_105(.A(desOut[39]), .Y(d_out_105));
CLKBUFX1 gbuf_q_105(.A(q_in_105), .Y(FP_R_27));
CLKBUFX1 gbuf_d_106(.A(desOut[37]), .Y(d_out_106));
CLKBUFX1 gbuf_q_106(.A(q_in_106), .Y(FP_R_19));
CLKBUFX1 gbuf_d_107(.A(desOut[1]), .Y(d_out_107));
CLKBUFX1 gbuf_q_107(.A(q_in_107), .Y(FP_R_7));
CLKBUFX1 gbuf_d_108(.A(desOut[61]), .Y(d_out_108));
CLKBUFX1 gbuf_q_108(.A(q_in_108), .Y(FP_R_16));
CLKBUFX1 gbuf_d_109(.A(desOut[7]), .Y(d_out_109));
CLKBUFX1 gbuf_q_109(.A(q_in_109), .Y(FP_R_31));
CLKBUFX1 gbuf_d_110(.A(desOut[55]), .Y(d_out_110));
CLKBUFX1 gbuf_q_110(.A(q_in_110), .Y(FP_R_25));
AND2X1 g16032(.A (n_1831), .B (n_2632), .Y (n_2977));
AND2X1 g16036(.A (n_1803), .B (n_2630), .Y (n_2973));
AOI22X1 g16041(.A0 (n_2588), .A1 (n_2613), .B0 (n_2954), .B1(n_2624), .Y (n_2970));
NAND2X1 g16042(.A (n_2593), .B (n_2591), .Y (n_2969));
INVX1 g16048(.A (n_2645), .Y (n_6101));
CLKBUFX1 gbuf_d_111(.A(desOut[29]), .Y(d_out_111));
CLKBUFX1 gbuf_q_111(.A(q_in_111), .Y(L_83));
NAND2X1 g16082(.A (n_2981), .B (n_2511), .Y (n_2966));
NAND2X1 g16085(.A (n_2949), .B (n_2668), .Y (n_2965));
NAND2X1 g16086(.A (n_2946), .B (n_2624), .Y (n_2964));
NAND2X1 g16124(.A (n_2958), .B (n_2668), .Y (n_2962));
NAND2X1 g16136(.A (n_2952), .B (n_2746), .Y (n_2960));
NAND2X1 g16150(.A (n_2958), .B (n_2613), .Y (n_2959));
AND2X1 g16154(.A (n_2956), .B (n_2613), .Y (n_2957));
NAND2X1 g16158(.A (n_2954), .B (n_2666), .Y (n_2955));
NAND2X1 g16159(.A (n_2952), .B (n_6600), .Y (n_2953));
NAND2X1 g16174(.A (n_2949), .B (n_2613), .Y (n_2950));
NAND2X1 g16175(.A (n_2946), .B (n_3153), .Y (n_2947));
NAND2X1 g16179(.A (n_1942), .B (n_2250), .Y (n_2944));
NAND2X1 g16189(.A (n_1435), .B (n_2981), .Y (n_2943));
AOI21X1 g16199(.A0 (n_1619), .A1 (n_2854), .B0 (n_7340), .Y (n_2941));
AOI21X1 g16201(.A0 (n_1767), .A1 (n_1616), .B0 (n_7437), .Y (n_2939));
AOI21X1 g16202(.A0 (n_2935), .A1 (n_2034), .B0 (n_7437), .Y (n_2936));
NAND2X1 g16204(.A (n_1957), .B (n_2931), .Y (n_2932));
AOI21X1 g16214(.A0 (n_2521), .A1 (n_2882), .B0 (n_253), .Y (n_2930));
NAND2X1 g16219(.A (n_1970), .B (n_2928), .Y (n_2929));
INVX1 g16223(.A (n_2559), .Y (n_2927));
AOI21X1 g16229(.A0 (n_1465), .A1 (n_1623), .B0 (n_1405), .Y (n_2926));
NAND2X1 g16231(.A (n_1989), .B (n_2171), .Y (n_2925));
NAND2X1 g16240(.A (n_1994), .B (n_7341), .Y (n_2923));
AOI21X1 g16243(.A0 (n_2794), .A1 (n_2105), .B0 (n_235), .Y (n_2921));
CLKBUFX1 gbuf_d_112(.A(desOut[27]), .Y(d_out_112));
CLKBUFX1 gbuf_q_112(.A(q_in_112), .Y(FP_R_12));
INVX1 g16246(.A (n_2543), .Y (n_2918));
NAND2X1 g16258(.A (n_1964), .B (n_2928), .Y (n_2917));
AOI21X1 g16262(.A0 (n_2347), .A1 (n_2137), .B0 (n_1405), .Y (n_2916));
NAND2X1 g16263(.A (n_1961), .B (n_2495), .Y (n_2915));
NAND2X1 g16264(.A (n_1959), .B (n_2913), .Y (n_2914));
NAND2X1 g16267(.A (n_1935), .B (n_7341), .Y (n_2912));
INVX1 g16269(.A (n_2528), .Y (n_2911));
AOI21X1 g16277(.A0 (n_2879), .A1 (n_7563), .B0 (n_7340), .Y (n_2909));
AOI21X1 g16280(.A0 (n_5732), .A1 (n_5921), .B0 (n_2907), .Y (n_2908));
AOI21X1 g16287(.A0 (n_6800), .A1 (n_2330), .B0 (n_235), .Y (n_2905));
NAND2X1 g16290(.A (n_1936), .B (n_7341), .Y (n_2903));
INVX1 g16295(.A (n_2512), .Y (n_2902));
CLKBUFX1 gbuf_d_113(.A(desOut[31]), .Y(d_out_113));
CLKBUFX1 gbuf_q_113(.A(q_in_113), .Y(FP_R_28));
NAND2X1 g16313(.A (n_1915), .B (n_2913), .Y (n_2900));
AOI21X1 g16317(.A0 (n_6058), .A1 (n_2882), .B0 (n_7437), .Y (n_2899));
AOI21X1 g16335(.A0 (n_2895), .A1 (n_2118), .B0 (n_7437), .Y (n_2898));
AOI21X1 g16341(.A0 (n_2935), .A1 (n_1846), .B0 (n_2813), .Y (n_2897));
AOI21X1 g16342(.A0 (n_2895), .A1 (n_1310), .B0 (n_6801), .Y (n_2896));
NAND2X1 g16345(.A (n_1976), .B (n_7301), .Y (n_2893));
NAND2X1 g16020(.A (n_2209), .B (n_2719), .Y (n_2892));
AOI21X1 g16362(.A0 (n_2888), .A1 (n_2456), .B0 (n_2042), .Y (n_2891));
AOI21X1 g16367(.A0 (n_2888), .A1 (n_2505), .B0 (n_440), .Y (n_2889));
CLKBUFX1 gbuf_d_114(.A(desOut[13]), .Y(d_out_114));
CLKBUFX1 gbuf_q_114(.A(q_in_114), .Y(FP_R_22));
AOI21X1 g16384(.A0 (n_1654), .A1 (n_7563), .B0 (n_6801), .Y (n_2886));
AOI21X1 g16386(.A0 (n_2408), .A1 (n_2882), .B0 (n_2050), .Y (n_2883));
AOI21X1 g16390(.A0 (n_6800), .A1 (n_2879), .B0 (n_2488), .Y (n_2881));
NAND2X1 g16391(.A (n_1991), .B (n_170), .Y (n_2878));
NAND2X1 g16403(.A (n_1974), .B (n_2666), .Y (n_2876));
NAND2X1 g16407(.A (n_2092), .B (n_170), .Y (n_2874));
NAND2X1 g16412(.A (n_2002), .B (n_2842), .Y (n_2872));
AOI21X1 g16424(.A0 (n_7559), .A1 (n_2550), .B0 (n_2488), .Y (n_2871));
INVX1 g17863(.A (desOut[23]), .Y (n_2870));
AOI21X1 g16429(.A0 (n_2839), .A1 (n_2836), .B0 (n_2067), .Y (n_2868));
AOI21X1 g16435(.A0 (n_1997), .A1 (n_7563), .B0 (n_440), .Y (n_2867));
NAND2X1 g16439(.A (n_1913), .B (n_2464), .Y (n_2865));
NAND2X1 g16442(.A (n_1968), .B (n_2863), .Y (n_2864));
NAND2X1 g16444(.A (n_1967), .B (n_2680), .Y (n_2862));
NAND2X1 g16445(.A (n_1944), .B (n_2680), .Y (n_2860));
NAND2X1 g16447(.A (n_1922), .B (n_177), .Y (n_2859));
NAND2X1 g16450(.A (n_1962), .B (n_7301), .Y (n_7891));
NAND2X1 g16456(.A (n_1958), .B (n_2856), .Y (n_2857));
AOI21X1 g16477(.A0 (n_2105), .A1 (n_2854), .B0 (n_2042), .Y (n_2855));
AOI21X1 g16484(.A0 (n_1528), .A1 (n_2557), .B0 (n_2067), .Y (n_2852));
INVX1 g17856(.A (n_7458), .Y (desOut[19]));
NAND2X1 g16494(.A (n_1919), .B (n_3194), .Y (n_2850));
NAND2X1 g16495(.A (n_1986), .B (n_2811), .Y (n_2848));
NAND2X1 g16497(.A (n_2157), .B (n_177), .Y (n_2847));
NAND2X1 g16504(.A (n_1930), .B (n_2735), .Y (n_2845));
NAND2X1 g16508(.A (n_1982), .B (n_2842), .Y (n_2843));
NAND2X1 g16511(.A (n_1926), .B (n_170), .Y (n_2841));
AOI21X1 g16518(.A0 (n_2839), .A1 (n_2838), .B0 (n_274), .Y (n_2840));
AOI21X1 g16520(.A0 (n_2366), .A1 (n_2836), .B0 (n_329), .Y (n_2837));
CLKBUFX1 gbuf_d_115(.A(desOut[15]), .Y(d_out_115));
CLKBUFX1 gbuf_q_115(.A(q_in_115), .Y(FP_R_30));
AOI21X1 g16522(.A0 (n_2839), .A1 (n_2806), .B0 (n_200), .Y (n_2834));
NAND2X1 g16526(.A (n_2098), .B (n_3159), .Y (n_2833));
NAND2X1 g16529(.A (n_1928), .B (n_2842), .Y (n_2832));
AOI21X1 g16532(.A0 (n_1578), .A1 (n_2830), .B0 (n_2440), .Y (n_2831));
NAND2X1 g16533(.A (n_1937), .B (n_3121), .Y (n_2829));
NAND2X1 g16535(.A (n_1924), .B (n_3044), .Y (n_2828));
NAND2X1 g16538(.A (n_1921), .B (n_170), .Y (n_2827));
NAND2X1 g16550(.A (n_2008), .B (n_3049), .Y (n_2826));
AOI21X1 g16552(.A0 (n_2374), .A1 (n_2830), .B0 (n_281), .Y (n_2825));
NAND2X1 g16566(.A (n_1917), .B (n_7301), .Y (n_2824));
AOI21X1 g16573(.A0 (n_6065), .A1 (n_1528), .B0 (n_6801), .Y (n_2822));
NAND2X1 g16576(.A (n_1993), .B (n_3044), .Y (n_2819));
NAND2X1 g16579(.A (n_1985), .B (n_2680), .Y (n_2818));
NAND2X1 g16580(.A (n_1996), .B (n_1882), .Y (n_2817));
AOI21X1 g16591(.A0 (n_7451), .A1 (n_1619), .B0 (n_2050), .Y (n_2815));
AOI21X1 g16592(.A0 (n_2131), .A1 (n_2879), .B0 (n_2813), .Y (n_2814));
NAND2X1 g16594(.A (n_2003), .B (n_2811), .Y (n_2812));
NAND2X1 g16608(.A (n_1912), .B (n_2811), .Y (n_2810));
AOI21X1 g16626(.A0 (n_1656), .A1 (n_2882), .B0 (n_2488), .Y (n_2809));
AOI21X1 g16640(.A0 (n_2806), .A1 (n_1616), .B0 (n_6801), .Y (n_2807));
NAND2X1 g16641(.A (n_1933), .B (n_177), .Y (n_2805));
CLKBUFX1 gbuf_d_116(.A(desOut[13]), .Y(d_out_116));
CLKBUFX1 gbuf_q_116(.A(q_in_116), .Y(L_85));
CLKBUFX1 gbuf_d_117(.A(desOut[27]), .Y(d_out_117));
CLKBUFX1 gbuf_q_117(.A(q_in_117), .Y(L_75));
CLKBUFX1 gbuf_d_118(.A(desOut[45]), .Y(d_out_118));
CLKBUFX1 gbuf_q_118(.A(q_in_118), .Y(L_81));
CLKBUFX1 gbuf_d_119(.A(desOut[11]), .Y(d_out_119));
CLKBUFX1 gbuf_qn_119(.A(qn_in_119), .Y(L_77));
NAND2X1 g16717(.A (n_2542), .B (n_1948), .Y (n_2802));
CLKBUFX1 gbuf_d_120(.A(desOut[11]), .Y(d_out_120));
CLKBUFX1 gbuf_q_120(.A(q_in_120), .Y(FP_R_14));
NAND2X1 g16856(.A (n_2526), .B (n_2793), .Y (n_2801));
NAND2X1 g16888(.A (n_2396), .B (n_2558), .Y (n_2800));
OR2X1 g16972(.A (n_1422), .B (n_1470), .Y (n_2799));
NAND2X1 g16978(.A (n_2363), .B (n_2389), .Y (n_2798));
NAND2X1 g17005(.A (n_1948), .B (n_2368), .Y (n_2797));
NAND2X1 g17010(.A (n_2794), .B (n_2793), .Y (n_2795));
OR2X1 g17022(.A (n_1437), .B (n_1885), .Y (n_2792));
NAND2X1 g17090(.A (n_2793), .B (n_2499), .Y (n_2789));
NAND2X1 g17110(.A (n_2396), .B (n_1454), .Y (n_2788));
MX2X1 g15516(.A (FP_R_60), .B (n_1241), .S0 (n_1260), .Y (n_2787));
NAND2X1 g15550(.A (n_1858), .B (n_1887), .Y (n_2786));
NAND3X1 g15561(.A (n_1886), .B (n_1835), .C (n_1809), .Y (n_2785));
NAND2X1 g15603(.A (n_1856), .B (n_1879), .Y (n_2782));
INVX1 g17814(.A (n_2781), .Y (desOut[41]));
INVX1 g17820(.A (n_2783), .Y (desOut[51]));
INVX1 g17834(.A (n_2790), .Y (desOut[17]));
NAND2X1 g15611(.A (n_7903), .B (n_7904), .Y (n_2777));
INVX1 g17817(.A (n_2778), .Y (desOut[53]));
INVX1 g17879(.A (n_2776), .Y (desOut[21]));
NAND2X1 g15640(.A (n_1853), .B (n_1862), .Y (n_2774));
CLKBUFX1 gbuf_d_121(.A(desOut[15]), .Y(d_out_121));
CLKBUFX1 gbuf_q_121(.A(q_in_121), .Y(L_93));
AOI21X1 g15667(.A0 (n_1255), .A1 (n_2134), .B0 (n_1850), .Y (n_2770));
INVX1 g17964(.A (n_2769), .Y (desOut[49]));
AOI21X1 g15685(.A0 (n_1633), .A1 (n_3121), .B0 (n_2147), .Y (n_2767));
AOI21X1 g15686(.A0 (n_1652), .A1 (n_7301), .B0 (n_2204), .Y (n_2766));
AOI21X1 g15694(.A0 (n_1537), .A1 (n_2692), .B0 (n_1375), .Y (n_2765));
NAND2X1 g15696(.A (n_2666), .B (n_2763), .Y (n_2764));
AOI21X1 g15703(.A0 (n_1713), .A1 (n_2752), .B0 (n_1755), .Y (n_2762));
AOI21X1 g15708(.A0 (n_1659), .A1 (n_2432), .B0 (n_2138), .Y (n_2761));
AOI21X1 g15716(.A0 (n_1475), .A1 (n_3189), .B0 (n_1749), .Y (n_2759));
NAND2X1 g15718(.A (n_2194), .B (n_1744), .Y (n_2757));
AOI21X1 g15728(.A0 (n_1604), .A1 (n_2752), .B0 (n_2119), .Y (n_2753));
AOI21X1 g15735(.A0 (n_1324), .A1 (n_3049), .B0 (n_2117), .Y (n_2751));
NAND2X1 g15737(.A (n_2114), .B (n_2113), .Y (n_2749));
NAND2X1 g15743(.A (n_2747), .B (n_2746), .Y (n_2748));
AOI21X1 g15751(.A0 (n_1594), .A1 (n_2842), .B0 (n_2107), .Y (n_2743));
AOI21X1 g15755(.A0 (n_1539), .A1 (n_2842), .B0 (n_2061), .Y (n_2742));
AOI21X1 g15756(.A0 (n_1605), .A1 (n_7301), .B0 (n_1390), .Y (n_5669));
AOI21X1 g15762(.A0 (n_1527), .A1 (n_1745), .B0 (n_1766), .Y (n_2740));
AOI21X1 g15763(.A0 (n_1679), .A1 (n_2746), .B0 (n_2188), .Y (n_7801));
AOI21X1 g15769(.A0 (n_1621), .A1 (n_204), .B0 (n_2166), .Y (n_2738));
AOI21X1 g15771(.A0 (n_1321), .A1 (n_2624), .B0 (n_2056), .Y (n_2737));
AOI21X1 g15775(.A0 (n_1690), .A1 (n_2735), .B0 (n_2028), .Y (n_2736));
AOI21X1 g15777(.A0 (n_1657), .A1 (n_2548), .B0 (n_2148), .Y (n_2734));
AOI21X1 g15779(.A0 (n_1608), .A1 (n_2666), .B0 (n_2179), .Y (n_6083));
AOI21X1 g15780(.A0 (n_1575), .A1 (n_7301), .B0 (n_2181), .Y (n_6091));
AOI21X1 g15788(.A0 (n_1506), .A1 (n_7301), .B0 (n_2090), .Y (n_2729));
AOI21X1 g15790(.A0 (n_1516), .A1 (n_3044), .B0 (n_2089), .Y (n_2728));
AOI21X1 g15791(.A0 (n_1577), .A1 (n_204), .B0 (n_2087), .Y (n_2727));
AOI21X1 g15794(.A0 (n_1689), .A1 (n_2863), .B0 (n_2084), .Y (n_2726));
AOI21X1 g15796(.A0 (n_1335), .A1 (n_7344), .B0 (n_2079), .Y (n_2725));
AOI21X1 g15797(.A0 (n_1570), .A1 (n_189), .B0 (n_2081), .Y (n_2723));
NOR2X1 g15798(.A (n_2075), .B (n_1735), .Y (n_2721));
AOI21X1 g15799(.A0 (n_1328), .A1 (n_2719), .B0 (n_2076), .Y (n_2720));
NOR2X1 g15805(.A (n_1379), .B (n_2073), .Y (n_5969));
NOR2X1 g15807(.A (n_2176), .B (n_1436), .Y (n_2717));
AOI21X1 g15815(.A0 (n_1561), .A1 (n_2410), .B0 (n_2071), .Y (n_2716));
NAND2X1 g18232(.A (n_3677), .B (desIn[32]), .Y (n_2715));
AOI21X1 g15817(.A0 (n_1560), .A1 (n_3049), .B0 (n_2173), .Y (n_2713));
NAND2X1 g18243(.A (n_3677), .B (desIn[20]), .Y (n_2712));
NOR2X1 g15845(.A (n_2066), .B (n_1409), .Y (n_2711));
AOI21X1 g15847(.A0 (n_1668), .A1 (n_2284), .B0 (n_2141), .Y (n_5694));
AOI21X1 g15848(.A0 (n_1601), .A1 (n_2467), .B0 (n_1779), .Y (n_2709));
NOR2X1 g15850(.A (n_1872), .B (n_2055), .Y (n_2708));
AOI21X1 g15851(.A0 (n_1521), .A1 (n_6805), .B0 (n_2169), .Y (n_5971));
AOI21X1 g15852(.A0 (n_1531), .A1 (n_7301), .B0 (n_2123), .Y (n_2705));
AOI21X1 g15853(.A0 (n_1509), .A1 (n_2719), .B0 (n_1725), .Y (n_2704));
AOI21X1 g15855(.A0 (n_1639), .A1 (n_2490), .B0 (n_2052), .Y (n_2702));
AOI21X1 g15858(.A0 (n_1486), .A1 (n_3194), .B0 (n_2096), .Y (n_2701));
AOI21X1 g15859(.A0 (n_1507), .A1 (n_2719), .B0 (n_2139), .Y (n_2700));
AOI21X1 g15861(.A0 (n_1137), .A1 (n_7341), .B0 (n_2047), .Y (n_2699));
CLKBUFX1 gbuf_d_122(.A(desOut[29]), .Y(d_out_122));
CLKBUFX1 gbuf_q_122(.A(q_in_122), .Y(FP_R_20));
AOI21X1 g15878(.A0 (n_1615), .A1 (n_2735), .B0 (n_1370), .Y (n_2694));
CLKBUFX1 gbuf_d_123(.A(desOut[31]), .Y(d_out_123));
CLKBUFX1 gbuf_q_123(.A(q_in_123), .Y(L_91));
AOI21X1 g15887(.A0 (n_1501), .A1 (n_2692), .B0 (n_2037), .Y (n_2693));
AOI21X1 g15889(.A0 (n_1498), .A1 (n_2752), .B0 (n_2035), .Y (n_2689));
AOI21X1 g15900(.A0 (n_1132), .A1 (n_2719), .B0 (n_2027), .Y (n_2688));
NAND2X1 g15904(.A (n_2155), .B (n_1706), .Y (n_2685));
AOI21X1 g15905(.A0 (n_1490), .A1 (n_2856), .B0 (n_2154), .Y (n_2684));
AOI21X1 g15908(.A0 (n_1545), .A1 (n_2863), .B0 (n_2025), .Y (n_2682));
AOI21X1 g15909(.A0 (n_1489), .A1 (n_2680), .B0 (n_1280), .Y (n_5620));
AOI21X1 g15915(.A0 (n_1161), .A1 (n_7341), .B0 (n_2022), .Y (n_2678));
AOI21X1 g15918(.A0 (n_1500), .A1 (n_177), .B0 (n_2149), .Y (n_2676));
AOI21X1 g15920(.A0 (n_1487), .A1 (n_2692), .B0 (n_2170), .Y (n_2674));
AOI21X1 g15928(.A0 (n_985), .A1 (n_2546), .B0 (n_2064), .Y (n_2673));
AOI21X1 g15945(.A0 (n_2671), .A1 (n_2624), .B0 (n_2145), .Y (n_2672));
NAND2X1 g15946(.A (n_2241), .B (n_1742), .Y (n_2670));
AOI21X1 g15957(.A0 (n_2236), .A1 (n_2668), .B0 (n_2097), .Y (n_7649));
AOI21X1 g15959(.A0 (n_2666), .A1 (n_2616), .B0 (n_2190), .Y (n_2667));
AOI21X1 g15967(.A0 (n_1419), .A1 (n_6600), .B0 (n_2177), .Y (n_2665));
AOI21X1 g15970(.A0 (n_2657), .A1 (n_2624), .B0 (n_1737), .Y (n_2664));
AOI21X1 g15976(.A0 (n_2604), .A1 (n_2668), .B0 (n_2065), .Y (n_2662));
AOI21X1 g15980(.A0 (n_2660), .A1 (n_2666), .B0 (n_2200), .Y (n_2661));
AOI21X1 g15982(.A0 (n_2598), .A1 (n_2746), .B0 (n_2053), .Y (n_5970));
AOI21X1 g15984(.A0 (n_2657), .A1 (n_2666), .B0 (n_1387), .Y (n_2658));
NAND2X1 g15987(.A (n_2218), .B (n_2045), .Y (n_2656));
NAND2X1 g15990(.A (n_2215), .B (n_2041), .Y (n_2655));
AOI21X1 g15993(.A0 (n_2572), .A1 (n_2653), .B0 (n_2159), .Y (n_2654));
NAND2X1 g16002(.A (n_2208), .B (n_1761), .Y (n_2652));
AOI21X1 g16005(.A0 (n_2633), .A1 (n_2746), .B0 (n_1730), .Y (n_2651));
AOI21X1 g16006(.A0 (n_2649), .A1 (n_2635), .B0 (n_2016), .Y (n_2650));
CLKBUFX1 gbuf_d_124(.A(desOut[45]), .Y(d_out_124));
CLKBUFX1 gbuf_q_124(.A(q_in_124), .Y(FP_R_18));
NAND2X1 g16049(.A (n_1807), .B (n_2230), .Y (n_2645));
NAND2X1 g16084(.A (n_2621), .B (n_2637), .Y (n_2644));
NAND2X1 g16087(.A (n_2577), .B (n_2974), .Y (n_2643));
NAND2X1 g16088(.A (n_2631), .B (n_2624), .Y (n_2642));
NAND2X1 g16090(.A (n_2639), .B (n_2746), .Y (n_2640));
NAND2X1 g16096(.A (n_2614), .B (n_2637), .Y (n_2638));
NAND2X1 g16098(.A (n_2629), .B (n_2635), .Y (n_2636));
NAND2X1 g16103(.A (n_2633), .B (n_2668), .Y (n_2634));
NAND2X1 g16104(.A (n_2631), .B (n_3153), .Y (n_2632));
NAND2X1 g16105(.A (n_2629), .B (n_3179), .Y (n_2630));
NAND2X1 g16106(.A (n_2581), .B (n_2637), .Y (n_2628));
NAND2X1 g16107(.A (n_2626), .B (n_2635), .Y (n_2627));
NAND2X1 g16108(.A (n_2569), .B (n_2624), .Y (n_2625));
NAND2X1 g16111(.A (n_2611), .B (n_6600), .Y (n_2623));
NAND2X1 g16113(.A (n_2621), .B (n_2974), .Y (n_2622));
NAND2X1 g16114(.A (n_2619), .B (n_2624), .Y (n_2620));
AND2X1 g16115(.A (n_2616), .B (n_2624), .Y (n_2617));
NAND2X1 g16116(.A (n_2614), .B (n_2613), .Y (n_2615));
NAND2X1 g16120(.A (n_2611), .B (n_2746), .Y (n_2612));
NAND2X1 g16132(.A (n_2590), .B (n_2666), .Y (n_2610));
NAND2X1 g16134(.A (n_2584), .B (n_2600), .Y (n_2609));
NAND2X1 g16137(.A (n_2586), .B (n_2666), .Y (n_2608));
NAND2X1 g16138(.A (n_2592), .B (n_2624), .Y (n_2607));
NAND2X1 g16139(.A (n_2604), .B (n_2974), .Y (n_2605));
NAND2X1 g16140(.A (n_2575), .B (n_2216), .Y (n_2603));
NAND2X1 g16141(.A (n_2579), .B (n_2666), .Y (n_5968));
NAND2X1 g16144(.A (n_2600), .B (n_2596), .Y (n_2601));
NAND2X1 g16146(.A (n_2598), .B (n_2668), .Y (n_2599));
AND2X1 g16147(.A (n_2596), .B (n_2746), .Y (n_2597));
NAND2X1 g16151(.A (n_2594), .B (n_2666), .Y (n_2595));
NAND2X1 g16152(.A (n_2592), .B (n_3179), .Y (n_2593));
NAND2X1 g16153(.A (n_2590), .B (n_2624), .Y (n_2591));
NAND2X1 g16157(.A (n_2588), .B (n_6600), .Y (n_6018));
NAND2X1 g16161(.A (n_2586), .B (n_2624), .Y (n_2587));
NAND2X1 g16162(.A (n_2584), .B (n_2746), .Y (n_2585));
CLKBUFX1 gbuf_d_125(.A(desOut[33]), .Y(d_out_125));
CLKBUFX1 gbuf_q_125(.A(q_in_125), .Y(FP_R_3));
NAND2X1 g16168(.A (n_2581), .B (n_2613), .Y (n_2582));
NAND2X1 g16171(.A (n_2579), .B (n_2624), .Y (n_2580));
NAND2X1 g16173(.A (n_2577), .B (n_2637), .Y (n_2578));
NAND2X1 g16180(.A (n_2575), .B (n_2974), .Y (n_2576));
CLKBUFX1 gbuf_d_126(.A(desOut[5]), .Y(d_out_126));
CLKBUFX1 gbuf_q_126(.A(q_in_126), .Y(FP_R_23));
NAND2X1 g16190(.A (n_2572), .B (n_2624), .Y (n_2573));
INVX2 g17892(.A (n_6379), .Y (desOut[3]));
NAND2X1 g16193(.A (n_2569), .B (n_3153), .Y (n_2570));
AOI21X1 g16196(.A0 (n_1578), .A1 (n_1988), .B0 (n_2182), .Y (n_2568));
AOI21X1 g16206(.A0 (n_7728), .A1 (n_1918), .B0 (n_235), .Y (n_2566));
NAND2X1 g16209(.A (n_1663), .B (n_2529), .Y (n_2565));
AOI21X1 g16210(.A0 (n_7445), .A1 (n_1404), .B0 (n_7340), .Y (n_2564));
NAND2X1 g16217(.A (n_1442), .B (n_2495), .Y (n_2562));
AOI21X1 g16222(.A0 (n_2029), .A1 (n_1330), .B0 (n_1405), .Y (n_2561));
AOI21X1 g16224(.A0 (n_2558), .A1 (n_2557), .B0 (n_2182), .Y (n_2559));
NAND2X1 g16226(.A (n_1642), .B (n_1760), .Y (n_2556));
NAND2X1 g16227(.A (n_1433), .B (n_7341), .Y (n_2555));
NAND2X1 g16232(.A (n_1638), .B (n_1760), .Y (n_2552));
AOI21X1 g16233(.A0 (n_2550), .A1 (n_2086), .B0 (n_198), .Y (n_2551));
NAND2X1 g16236(.A (n_1618), .B (n_2548), .Y (n_2549));
NAND2X1 g16238(.A (n_1549), .B (n_2546), .Y (n_2547));
NAND2X1 g16245(.A (n_1606), .B (n_204), .Y (n_2545));
AOI21X1 g16247(.A0 (n_2542), .A1 (n_2541), .B0 (n_191), .Y (n_2543));
NAND2X1 g16248(.A (n_1680), .B (n_2539), .Y (n_2540));
INVX1 g16249(.A (n_2185), .Y (n_2538));
NAND2X1 g16251(.A (n_1552), .B (n_2974), .Y (n_2537));
NAND2X1 g16252(.A (n_1589), .B (n_2913), .Y (n_2536));
NAND2X1 g16253(.A (n_1590), .B (n_2539), .Y (n_2535));
AOI21X1 g16254(.A0 (n_7732), .A1 (n_2347), .B0 (n_7340), .Y (n_2534));
AOI22X1 g17881(.A0 (n_1271), .A1 (n_1776), .B0 (n_2298), .B1(desIn[21]), .Y (n_2776));
NAND2X1 g16259(.A (n_1843), .B (n_7341), .Y (n_2532));
AOI21X1 g16261(.A0 (n_6022), .A1 (n_2422), .B0 (n_1405), .Y (n_2531));
NAND2X1 g16265(.A (n_1568), .B (n_2529), .Y (n_2530));
AOI21X1 g16270(.A0 (n_1656), .A1 (n_2526), .B0 (n_253), .Y (n_2528));
AOI21X1 g16275(.A0 (n_2396), .A1 (n_1312), .B0 (n_1405), .Y (n_2523));
AOI21X1 g16278(.A0 (n_2521), .A1 (n_1662), .B0 (n_2182), .Y (n_2522));
NAND2X1 g16281(.A (n_1544), .B (n_2171), .Y (n_2520));
AOI21X1 g16292(.A0 (n_2895), .A1 (n_1753), .B0 (n_235), .Y (n_2517));
NAND2X1 g16293(.A (n_1684), .B (n_1760), .Y (n_2516));
NAND2X1 g16294(.A (n_1768), .B (n_7341), .Y (n_2514));
AOI21X1 g16296(.A0 (n_1551), .A1 (n_2511), .B0 (n_2182), .Y (n_2512));
NAND2X1 g16300(.A (n_1669), .B (n_2928), .Y (n_2510));
AOI21X1 g16303(.A0 (n_2503), .A1 (n_6800), .B0 (n_198), .Y (n_2509));
AOI21X1 g16304(.A0 (n_2506), .A1 (n_2505), .B0 (n_2907), .Y (n_2507));
AOI21X1 g16310(.A0 (n_2329), .A1 (n_2503), .B0 (n_2182), .Y (n_2504));
NAND2X1 g16311(.A (n_1563), .B (n_2539), .Y (n_2502));
NAND2X1 g16312(.A (n_1502), .B (n_2913), .Y (n_2501));
AOI21X1 g16315(.A0 (n_2499), .A1 (n_5929), .B0 (n_2182), .Y (n_2500));
NAND2X1 g16318(.A (n_1530), .B (n_7341), .Y (n_2498));
NAND2X1 g16328(.A (n_1583), .B (n_2495), .Y (n_2496));
NAND2X1 g16333(.A (n_1782), .B (n_7436), .Y (n_2494));
AOI21X1 g16338(.A0 (n_2184), .A1 (n_2376), .B0 (n_2440), .Y (n_2493));
NAND2X1 g16346(.A (n_1613), .B (n_2863), .Y (n_2492));
NAND2X1 g16350(.A (n_1522), .B (n_2490), .Y (n_2491));
AOI21X1 g16354(.A0 (n_2363), .A1 (n_2422), .B0 (n_2488), .Y (n_2489));
NAND2X1 g16355(.A (n_1631), .B (n_1880), .Y (n_2487));
NAND2X1 g16357(.A (n_1646), .B (n_3044), .Y (n_2486));
NAND2X1 g16359(.A (n_1647), .B (n_2680), .Y (n_2484));
NAND2X1 g16360(.A (n_1532), .B (n_7301), .Y (n_2483));
NAND2X1 g16363(.A (n_1554), .B (n_3194), .Y (n_2482));
AOI21X1 g16364(.A0 (n_2453), .A1 (n_1152), .B0 (n_2122), .Y (n_2480));
NAND2X1 g16380(.A (n_1592), .B (n_2811), .Y (n_2479));
NAND2X1 g16381(.A (n_1678), .B (n_177), .Y (n_2477));
AOI21X1 g16389(.A0 (n_7732), .A1 (n_2054), .B0 (n_329), .Y (n_2476));
AOI21X1 g16392(.A0 (n_2542), .A1 (n_2456), .B0 (n_2440), .Y (n_2475));
NAND2X1 g16393(.A (n_1644), .B (n_2680), .Y (n_2474));
NAND2X1 g16394(.A (n_1643), .B (n_7301), .Y (n_2473));
NAND2X1 g16397(.A (n_1636), .B (n_2692), .Y (n_2472));
NAND2X1 g16400(.A (n_1518), .B (n_1882), .Y (n_2471));
NAND2X1 g16405(.A (n_1620), .B (n_170), .Y (n_2469));
NAND2X1 g16411(.A (n_1612), .B (n_2467), .Y (n_2468));
NAND2X1 g16416(.A (n_1534), .B (n_2752), .Y (n_2466));
NAND2X1 g16418(.A (n_1597), .B (n_2464), .Y (n_2465));
NAND2X1 g16425(.A (n_1617), .B (n_170), .Y (n_2463));
AOI21X1 g16427(.A0 (n_2895), .A1 (n_1651), .B0 (n_136), .Y (n_2461));
NAND2X1 g16428(.A (n_1526), .B (n_2464), .Y (n_2460));
OAI21X1 g17864(.A0 (n_1267), .A1 (n_2298), .B0 (n_919), .Y(desOut[23]));
NAND2X1 g16431(.A (n_1553), .B (n_7301), .Y (n_2459));
AOI21X1 g16432(.A0 (n_2356), .A1 (n_2456), .B0 (n_183), .Y (n_2457));
NAND2X1 g16433(.A (n_1587), .B (n_2402), .Y (n_2455));
AOI21X1 g16434(.A0 (n_2453), .A1 (n_5835), .B0 (n_6801), .Y (n_2454));
NAND2X1 g16436(.A (n_1585), .B (n_3189), .Y (n_2451));
NAND2X1 g16438(.A (n_1676), .B (n_3049), .Y (n_2449));
NAND2X1 g16440(.A (n_1586), .B (n_7301), .Y (n_2448));
NAND2X1 g16441(.A (n_1484), .B (n_2686), .Y (n_2447));
AOI21X1 g16443(.A0 (n_7446), .A1 (n_2557), .B0 (n_329), .Y (n_2446));
NAND2X1 g16446(.A (n_1582), .B (n_1882), .Y (n_2444));
NAND2X1 g16448(.A (n_1580), .B (n_2842), .Y (n_2443));
AOI21X1 g16453(.A0 (n_2558), .A1 (n_2499), .B0 (n_2440), .Y (n_2441));
NAND2X1 g16454(.A (n_1574), .B (n_6805), .Y (n_2439));
NAND2X1 g16455(.A (n_1571), .B (n_170), .Y (n_2438));
NAND2X1 g16458(.A (n_1584), .B (n_2436), .Y (n_2437));
NAND2X1 g16466(.A (n_1655), .B (n_3189), .Y (n_2435));
AOI21X1 g16467(.A0 (n_2124), .A1 (n_1656), .B0 (n_297), .Y (n_2434));
NAND2X1 g16468(.A (n_1567), .B (n_2432), .Y (n_2433));
AOI21X1 g16469(.A0 (n_1711), .A1 (n_2199), .B0 (n_2136), .Y (n_2431));
NAND2X1 g16472(.A (n_1564), .B (n_2719), .Y (n_2430));
AOI21X1 g16475(.A0 (n_7445), .A1 (n_5838), .B0 (n_127), .Y (n_2429));
AOI21X1 g16480(.A0 (n_7451), .A1 (n_2558), .B0 (n_274), .Y (n_2427));
AOI21X1 g16481(.A0 (n_2054), .A1 (n_2503), .B0 (n_275), .Y (n_2425));
AOI21X1 g16487(.A0 (n_2422), .A1 (n_6797), .B0 (n_2440), .Y (n_2423));
AOI21X1 g16490(.A0 (n_2131), .A1 (n_5908), .B0 (n_136), .Y (n_2420));
AOI21X1 g16491(.A0 (n_2174), .A1 (n_2309), .B0 (n_2813), .Y (n_2419));
AOI21X1 g16499(.A0 (n_2094), .A1 (n_2131), .B0 (n_2067), .Y (n_2417));
NAND2X1 g16501(.A (n_1672), .B (n_7301), .Y (n_2415));
NAND2X1 g16503(.A (n_1664), .B (n_2412), .Y (n_2413));
NAND2X1 g16505(.A (n_1525), .B (n_2410), .Y (n_2411));
AOI21X1 g16506(.A0 (n_2408), .A1 (n_2557), .B0 (n_2042), .Y (n_2409));
AOI21X1 g16507(.A0 (n_2526), .A1 (n_2558), .B0 (n_281), .Y (n_2407));
AND2X1 g16512(.A (n_1427), .B (n_177), .Y (n_2406));
NAND2X1 g16524(.A (n_1728), .B (n_2404), .Y (n_2405));
NAND2X1 g16536(.A (n_1519), .B (n_2402), .Y (n_2403));
NAND2X1 g16537(.A (n_1624), .B (n_2635), .Y (n_7799));
NAND2X1 g16540(.A (n_1515), .B (n_2686), .Y (n_2400));
NAND2X1 g16548(.A (n_1512), .B (n_2410), .Y (n_2399));
NAND2X1 g16555(.A (n_1576), .B (n_3134), .Y (n_2398));
AOI21X1 g16557(.A0 (n_2396), .A1 (n_6052), .B0 (n_2248), .Y (n_2397));
AOI21X1 g16562(.A0 (n_1948), .A1 (n_2311), .B0 (n_2440), .Y (n_2395));
NAND2X1 g16563(.A (n_1773), .B (n_2842), .Y (n_2394));
NAND2X1 g16565(.A (n_1488), .B (n_2464), .Y (n_2393));
AOI21X1 g16571(.A0 (n_2422), .A1 (n_1733), .B0 (n_127), .Y (n_2392));
AOI21X1 g16588(.A0 (n_2389), .A1 (n_2068), .B0 (n_274), .Y (n_2390));
AOI21X1 g16590(.A0 (n_2503), .A1 (n_2422), .B0 (n_297), .Y (n_2388));
NAND2X1 g16597(.A (n_1665), .B (n_2464), .Y (n_2387));
NAND2X1 g16598(.A (n_1635), .B (n_2695), .Y (n_2386));
NAND2X1 g16599(.A (n_1688), .B (n_2410), .Y (n_2385));
AOI21X1 g16602(.A0 (n_2836), .A1 (n_2505), .B0 (n_2050), .Y (n_2384));
AOI21X1 g16605(.A0 (n_2029), .A1 (n_2838), .B0 (n_2488), .Y (n_2383));
NAND2X1 g16606(.A (n_1599), .B (n_172), .Y (n_2381));
NAND2X1 g16616(.A (n_1673), .B (n_2412), .Y (n_2379));
NAND2X1 g16629(.A (n_1536), .B (n_2735), .Y (n_2378));
AOI21X1 g16632(.A0 (n_2376), .A1 (n_1551), .B0 (n_2488), .Y (n_2377));
AOI21X1 g16638(.A0 (n_2374), .A1 (n_2511), .B0 (n_2050), .Y (n_2375));
CLKBUFX1 gbuf_d_127(.A(desOut[33]), .Y(d_out_127));
CLKBUFX1 gbuf_q_127(.A(q_in_127), .Y(L_66));
CLKBUFX1 gbuf_d_128(.A(desOut[5]), .Y(d_out_128));
CLKBUFX1 gbuf_q_128(.A(q_in_128), .Y(L_86));
NAND2X1 g16696(.A (n_6065), .B (n_1619), .Y (n_2373));
NAND2X1 g16721(.A (n_2010), .B (n_1551), .Y (n_2371));
NAND2X1 g16723(.A (n_2839), .B (n_2368), .Y (n_2369));
NAND2X1 g16727(.A (n_2366), .B (n_2368), .Y (n_2367));
NAND2X1 g16751(.A (n_5835), .B (n_1528), .Y (n_2365));
NAND2X1 g16752(.A (n_2363), .B (n_7563), .Y (n_2364));
NAND2X1 g16767(.A (n_2046), .B (n_1619), .Y (n_2362));
NAND2X1 g16783(.A (n_5921), .B (n_2054), .Y (n_2361));
NAND2X1 g16787(.A (n_2010), .B (n_1627), .Y (n_2359));
NAND2X1 g16800(.A (n_2356), .B (n_1616), .Y (n_2357));
NAND2X1 g16804(.A (n_2888), .B (n_2039), .Y (n_2355));
NAND2X1 g16805(.A (n_1619), .B (n_2499), .Y (n_2354));
NAND2X1 g16806(.A (n_2118), .B (n_2034), .Y (n_2353));
NAND2X1 g16814(.A (n_2340), .B (n_1562), .Y (n_2351));
NAND2X1 g16822(.A (n_2376), .B (n_2034), .Y (n_2350));
NAND2X1 g16824(.A (n_2180), .B (n_7682), .Y (n_2349));
NAND2X1 g16840(.A (n_2330), .B (n_2347), .Y (n_2348));
OR2X1 g16857(.A (n_6799), .B (n_1256), .Y (n_2346));
NAND2X1 g16862(.A (n_2319), .B (n_1310), .Y (n_2345));
OR2X1 g16867(.A (n_1902), .B (n_1065), .Y (n_2344));
NAND2X1 g16908(.A (n_1670), .B (n_5921), .Y (n_2343));
NAND2X1 g16922(.A (n_2340), .B (n_1337), .Y (n_2341));
NAND2X1 g16927(.A (n_2542), .B (n_1821), .Y (n_2339));
NAND2X1 g16943(.A (n_5835), .B (n_1619), .Y (n_2337));
NAND2X1 g16951(.A (n_2882), .B (n_5929), .Y (n_2334));
OR2X1 g16963(.A (n_1854), .B (n_932), .Y (n_2332));
NAND2X1 g16966(.A (n_2330), .B (n_2329), .Y (n_2331));
NAND2X1 g16993(.A (n_2069), .B (n_2879), .Y (n_2326));
NAND2X1 g16996(.A (n_2422), .B (n_2137), .Y (n_2325));
NAND2X1 g16998(.A (n_2453), .B (n_2882), .Y (n_2324));
NAND2X1 g17013(.A (n_1767), .B (n_2366), .Y (n_3170));
OR2X1 g17023(.A (n_1005), .B (n_1911), .Y (n_2322));
AOI22X1 g17836(.A0 (n_1269), .A1 (n_1776), .B0 (n_2298), .B1(desIn[17]), .Y (n_2790));
NAND2X1 g17029(.A (n_2319), .B (n_2118), .Y (n_3154));
NAND2X1 g17030(.A (n_1562), .B (n_2118), .Y (n_2318));
NAND2X1 g17041(.A (n_2356), .B (n_7686), .Y (n_2317));
NAND2X1 g17075(.A (n_1846), .B (n_2118), .Y (n_2316));
NAND2X1 g17081(.A (n_7446), .B (n_2882), .Y (n_2315));
NAND2X1 g17082(.A (n_1616), .B (n_2838), .Y (n_2314));
NAND2X1 g17086(.A (n_5921), .B (n_7559), .Y (n_2313));
NAND2X1 g17089(.A (n_1821), .B (n_2311), .Y (n_2312));
AOI21X1 g16585(.A0 (n_2054), .A1 (n_2309), .B0 (n_2067), .Y (n_2310));
NAND2X1 g17100(.A (n_5921), .B (n_2329), .Y (n_2307));
OR2X1 g17106(.A (n_1481), .B (n_1541), .Y (n_2306));
NAND2X1 g17107(.A (n_2542), .B (n_2839), .Y (n_2305));
NAND2X1 g17124(.A (n_2203), .B (n_1310), .Y (n_2304));
CLKBUFX1 g17831(.A (n_6635), .Y (desOut[9]));
AOI21X1 g17966(.A0 (n_3677), .A1 (desIn[49]), .B0 (n_1445), .Y(n_2769));
AOI22X1 g17822(.A0 (n_1294), .A1 (n_879), .B0 (n_2298), .B1(desIn[51]), .Y (n_2783));
AOI22X1 g17819(.A0 (n_1290), .A1 (n_1776), .B0 (n_755), .B1(desIn[53]), .Y (n_2778));
INVX1 g17869(.A (n_2293), .Y (desOut[47]));
AOI22X1 g17816(.A0 (n_1276), .A1 (n_879), .B0 (n_701), .B1(desIn[41]), .Y (n_2781));
AOI21X1 g15655(.A0 (n_1414), .A1 (n_2281), .B0 (n_1363), .Y (n_2291));
INVX1 g17975(.A (desOut[59]), .Y (n_3829));
INVX1 g17976(.A (desOut[59]), .Y (n_2287));
INVX1 g17967(.A (n_2289), .Y (desOut[43]));
INVX1 g17997(.A (n_6978), .Y (desOut[55]));
AOI21X1 g15695(.A0 (n_1259), .A1 (n_2284), .B0 (n_1408), .Y (n_5668));
AOI21X1 g15699(.A0 (n_1139), .A1 (n_2284), .B0 (n_1697), .Y (n_2283));
AOI21X1 g15713(.A0 (n_1352), .A1 (n_2281), .B0 (n_1751), .Y (n_2282));
NAND2X1 g15719(.A (n_1783), .B (n_1743), .Y (n_2280));
AOI21X1 g15765(.A0 (n_920), .A1 (n_1719), .B0 (n_1762), .Y (n_5695));
NAND2X1 g17109(.A (n_2854), .B (n_1528), .Y (n_2278));
AOI21X1 g15776(.A0 (n_1350), .A1 (n_2666), .B0 (n_1722), .Y (n_7802));
NAND2X1 g15837(.A (n_1709), .B (n_1726), .Y (n_2276));
NAND2X1 g15869(.A (n_1720), .B (n_1716), .Y (n_2275));
NAND2X1 g15870(.A (n_1715), .B (n_1443), .Y (n_2273));
AOI21X1 g15898(.A0 (n_1281), .A1 (n_2842), .B0 (n_1393), .Y (n_2271));
AOI21X1 g15902(.A0 (n_1320), .A1 (n_2624), .B0 (n_1367), .Y (n_2269));
NAND2X1 g15914(.A (n_1701), .B (n_1759), .Y (n_2267));
NAND2X1 g15923(.A (n_1699), .B (n_1698), .Y (n_2266));
NAND2X1 g15927(.A (n_1695), .B (n_1694), .Y (n_2265));
NAND2X1 g15930(.A (n_1757), .B (n_1758), .Y (n_2264));
AOI21X1 g15941(.A0 (n_1811), .A1 (n_2600), .B0 (n_1708), .Y (n_2263));
NAND2X1 g17098(.A (n_2029), .B (n_1686), .Y (n_2261));
AOI21X1 g15989(.A0 (n_2257), .A1 (n_2666), .B0 (n_1219), .Y (n_2258));
NAND2X1 g16001(.A (n_1791), .B (n_1707), .Y (n_2256));
NAND2X1 g16007(.A (n_1785), .B (n_1700), .Y (n_2254));
AOI21X1 g16022(.A0 (n_1767), .A1 (n_2250), .B0 (n_2036), .Y (n_2253));
AOI21X1 g16018(.A0 (n_1572), .A1 (n_1361), .B0 (n_2144), .Y (n_2252));
AOI21X1 g16024(.A0 (n_1538), .A1 (n_2245), .B0 (n_2248), .Y (n_2249));
AOI22X1 g16027(.A0 (n_1851), .A1 (n_3153), .B0 (n_2207), .B1(n_2613), .Y (n_2247));
AOI21X1 g16023(.A0 (n_2180), .A1 (n_2245), .B0 (n_240), .Y (n_2246));
NAND2X1 g16079(.A (n_2245), .B (n_1279), .Y (n_2747));
NAND2X1 g16081(.A (n_2221), .B (n_2668), .Y (n_2242));
NAND2X1 g16083(.A (n_1134), .B (n_2245), .Y (n_2763));
NAND2X1 g16089(.A (n_2205), .B (n_2666), .Y (n_2241));
NAND2X1 g16092(.A (n_2238), .B (n_2600), .Y (n_2239));
NAND2X1 g16099(.A (n_2236), .B (n_2746), .Y (n_2237));
NAND2X1 g16118(.A (n_2233), .B (n_6600), .Y (n_2234));
NAND2X1 g16119(.A (n_2228), .B (n_2746), .Y (n_2232));
INVX1 g18525(.A (n_3625), .Y (n_3631));
NAND2X1 g16125(.A (n_2214), .B (n_2746), .Y (n_2230));
NAND2X1 g16126(.A (n_2228), .B (n_6600), .Y (n_2229));
NAND2X1 g16127(.A (n_2217), .B (n_2974), .Y (n_2227));
NAND2X1 g16131(.A (n_2219), .B (n_2624), .Y (n_2226));
AOI21X1 g16519(.A0 (n_6797), .A1 (n_2347), .B0 (n_275), .Y (n_2225));
NAND2X1 g16148(.A (n_2212), .B (n_2746), .Y (n_2223));
NAND2X1 g16160(.A (n_2221), .B (n_2746), .Y (n_2222));
NAND2X1 g16163(.A (n_2219), .B (n_2653), .Y (n_7887));
NAND2X1 g16169(.A (n_2217), .B (n_2216), .Y (n_2218));
NAND2X1 g16172(.A (n_2214), .B (n_2637), .Y (n_2215));
NAND2X1 g16178(.A (n_2212), .B (n_2668), .Y (n_2213));
NAND2X1 g16181(.A (n_1215), .B (n_2245), .Y (n_2211));
NAND2X1 g16186(.A (n_863), .B (n_2245), .Y (n_2209));
NAND2X1 g16191(.A (n_2207), .B (n_2216), .Y (n_2208));
NAND2X1 g16194(.A (n_2205), .B (n_2624), .Y (n_2206));
AOI21X1 g16195(.A0 (n_1847), .A1 (n_2203), .B0 (n_7437), .Y (n_2204));
AOI21X1 g16203(.A0 (n_2183), .A1 (n_1627), .B0 (n_235), .Y (n_2201));
AOI21X1 g16205(.A0 (n_2199), .A1 (n_2094), .B0 (n_2182), .Y (n_2200));
AOI21X1 g16207(.A0 (n_2124), .A1 (n_6060), .B0 (n_2182), .Y (n_2198));
NAND2X1 g16212(.A (n_1336), .B (n_189), .Y (n_2196));
AOI21X1 g16213(.A0 (n_2178), .A1 (n_1499), .B0 (n_1405), .Y (n_2195));
NAND2X1 g16215(.A (n_1347), .B (n_7436), .Y (n_2194));
NAND2X1 g16234(.A (n_1317), .B (n_2746), .Y (n_2193));
AOI21X1 g16237(.A0 (n_2146), .A1 (n_2165), .B0 (n_2907), .Y (n_2191));
AOI21X1 g16239(.A0 (n_1623), .A1 (n_2029), .B0 (n_7340), .Y (n_2190));
NAND2X1 g16242(.A (n_1356), .B (n_7341), .Y (n_7798));
AOI21X1 g16244(.A0 (n_6567), .A1 (n_1550), .B0 (n_7340), .Y (n_2188));
AOI21X1 g16250(.A0 (n_2184), .A1 (n_2183), .B0 (n_2182), .Y (n_2185));
AOI21X1 g16255(.A0 (n_2180), .A1 (n_1543), .B0 (n_1777), .Y (n_2181));
INVX1 g17883(.A (desOut[37]), .Y (n_2544));
AOI21X1 g16257(.A0 (n_2101), .A1 (n_2178), .B0 (n_191), .Y (n_2179));
AOI21X1 g16260(.A0 (n_2046), .A1 (n_953), .B0 (n_2151), .Y (n_2177));
AOI21X1 g16268(.A0 (n_1770), .A1 (n_2034), .B0 (n_235), .Y (n_2176));
AOI21X1 g16271(.A0 (n_2174), .A1 (n_2137), .B0 (n_1777), .Y (n_2175));
AOI21X1 g16274(.A0 (n_2083), .A1 (n_2105), .B0 (n_198), .Y (n_2173));
NAND2X1 g16289(.A (n_1311), .B (n_2171), .Y (n_2172));
AOI21X1 g16291(.A0 (n_1649), .A1 (n_1634), .B0 (n_7340), .Y (n_2170));
AOI21X1 g16301(.A0 (n_1312), .A1 (n_1972), .B0 (n_7340), .Y (n_2169));
AOI21X1 g16302(.A0 (n_1943), .A1 (n_2165), .B0 (n_253), .Y (n_2166));
NAND2X1 g16305(.A (n_1334), .B (n_189), .Y (n_2163));
AOI21X1 g16306(.A0 (n_921), .A1 (n_2078), .B0 (n_198), .Y (n_2162));
AOI21X1 g16314(.A0 (n_2118), .A1 (n_1667), .B0 (n_7340), .Y (n_2159));
AOI21X1 g16316(.A0 (n_1656), .A1 (n_6065), .B0 (n_2907), .Y (n_2158));
NAND2X1 g16971(.A (n_2124), .B (n_1351), .Y (n_2157));
NAND2X1 g16322(.A (n_1319), .B (n_2529), .Y (n_2155));
AOI21X1 g16323(.A0 (n_1686), .A1 (n_1727), .B0 (n_1405), .Y (n_2154));
AOI21X1 g16326(.A0 (n_1573), .A1 (n_1703), .B0 (n_2151), .Y (n_2152));
NAND2X1 g16330(.A (n_1327), .B (n_2539), .Y (n_2150));
AOI21X1 g16331(.A0 (n_2184), .A1 (n_2178), .B0 (n_7437), .Y (n_2149));
AOI21X1 g16336(.A0 (n_1528), .A1 (n_1972), .B0 (n_1405), .Y (n_2148));
AOI21X1 g16339(.A0 (n_2146), .A1 (n_2311), .B0 (n_2067), .Y (n_2147));
AOI21X1 g16343(.A0 (n_2074), .A1 (n_5912), .B0 (n_2144), .Y (n_2145));
INVX1 g17873(.A (desOut[45]), .Y (n_2143));
AOI21X1 g16348(.A0 (n_863), .A1 (n_2020), .B0 (n_207), .Y (n_2141));
AOI21X1 g16349(.A0 (n_7728), .A1 (n_7559), .B0 (n_2248), .Y (n_2139));
AOI21X1 g16356(.A0 (n_1388), .A1 (n_2137), .B0 (n_2136), .Y (n_2138));
NAND2X1 g16358(.A (n_1359), .B (n_2134), .Y (n_2135));
AOI21X1 g16361(.A0 (n_6022), .A1 (n_2131), .B0 (n_6801), .Y (n_2133));
AOI21X1 g16366(.A0 (n_1645), .A1 (n_7733), .B0 (n_6801), .Y (n_2130));
AOI21X1 g16368(.A0 (n_1578), .A1 (n_1279), .B0 (n_234), .Y (n_2129));
AOI22X1 g17871(.A0 (n_1026), .A1 (n_879), .B0 (n_701), .B1(desIn[47]), .Y (n_2293));
NAND2X1 g16372(.A (n_1323), .B (n_1719), .Y (n_2126));
AOI21X1 g16376(.A0 (n_2124), .A1 (n_1163), .B0 (n_2036), .Y (n_2125));
AOI21X1 g16377(.A0 (n_6070), .A1 (n_5924), .B0 (n_2122), .Y (n_2123));
AOI21X1 g16378(.A0 (n_5722), .A1 (n_2137), .B0 (n_127), .Y (n_2121));
NAND2X1 g16964(.A (n_2091), .B (n_1330), .Y (n_2956));
AOI21X1 g16382(.A0 (n_6070), .A1 (n_1312), .B0 (n_2136), .Y (n_2120));
AOI21X1 g16385(.A0 (n_1578), .A1 (n_2118), .B0 (n_329), .Y (n_2119));
AOI21X1 g16395(.A0 (n_1649), .A1 (n_2100), .B0 (n_274), .Y (n_2117));
NAND2X1 g16398(.A (n_1344), .B (n_2281), .Y (n_2114));
NAND2X1 g16399(.A (n_1338), .B (n_2719), .Y (n_2113));
AOI21X1 g16404(.A0 (n_2010), .A1 (n_1562), .B0 (n_1750), .Y (n_2112));
NAND2X1 g16406(.A (n_1348), .B (n_3044), .Y (n_2110));
NAND2X1 g16410(.A (n_1362), .B (n_2134), .Y (n_2109));
AOI21X1 g16413(.A0 (n_1943), .A1 (n_2023), .B0 (n_2440), .Y (n_2108));
AOI21X1 g16414(.A0 (n_1662), .A1 (n_2105), .B0 (n_136), .Y (n_2107));
NAND2X1 g16415(.A (n_1373), .B (n_3044), .Y (n_2104));
NAND2X1 g16419(.A (n_1322), .B (n_2436), .Y (n_2103));
AOI21X1 g16421(.A0 (n_2101), .A1 (n_2100), .B0 (n_2042), .Y (n_2102));
NAND2X1 g17136(.A (n_2039), .B (n_2506), .Y (n_2098));
AOI21X1 g16426(.A0 (n_2010), .A1 (n_1649), .B0 (n_183), .Y (n_2097));
AOI21X1 g16430(.A0 (n_2165), .A1 (n_2024), .B0 (n_274), .Y (n_2096));
AOI21X1 g16437(.A0 (n_2094), .A1 (n_5732), .B0 (n_2440), .Y (n_2095));
NAND2X1 g17027(.A (n_2091), .B (n_2506), .Y (n_2092));
AOI21X1 g16449(.A0 (n_914), .A1 (n_7559), .B0 (n_2042), .Y (n_2090));
AOI21X1 g16451(.A0 (n_1619), .A1 (n_1972), .B0 (n_127), .Y (n_2089));
AOI21X1 g16452(.A0 (n_2086), .A1 (n_2137), .B0 (n_183), .Y (n_2087));
AOI21X1 g16457(.A0 (n_1528), .A1 (n_2083), .B0 (n_274), .Y (n_2084));
AOI21X1 g16459(.A0 (n_1351), .A1 (n_1640), .B0 (n_2144), .Y (n_2081));
AOI21X1 g16461(.A0 (n_1351), .A1 (n_2078), .B0 (n_6801), .Y (n_2079));
AOI21X1 g16462(.A0 (n_1645), .A1 (n_1258), .B0 (n_2440), .Y (n_2076));
AOI21X1 g16463(.A0 (n_2074), .A1 (n_6567), .B0 (n_2440), .Y (n_2075));
INVX1 g17849(.A (desOut[1]), .Y (n_2380));
AOI21X1 g16474(.A0 (n_1660), .A1 (n_2074), .B0 (n_6801), .Y (n_2073));
NAND2X1 g16476(.A (n_1326), .B (n_1719), .Y (n_2072));
AOI21X1 g16483(.A0 (n_2094), .A1 (n_2086), .B0 (n_274), .Y (n_2071));
AOI21X1 g16485(.A0 (n_2069), .A1 (n_2068), .B0 (n_2067), .Y (n_2070));
AOI21X1 g16486(.A0 (n_2018), .A1 (n_981), .B0 (n_2248), .Y (n_2066));
AOI21X1 g16500(.A0 (n_7446), .A1 (n_6065), .B0 (n_440), .Y (n_2065));
AOI21X1 g16502(.A0 (n_2060), .A1 (n_1573), .B0 (n_127), .Y (n_2064));
AOI21X1 g16510(.A0 (n_1943), .A1 (n_2368), .B0 (n_2813), .Y (n_2063));
AOI21X1 g16513(.A0 (n_2060), .A1 (n_7702), .B0 (n_2440), .Y (n_2061));
AOI21X1 g16527(.A0 (n_7664), .A1 (n_2183), .B0 (n_234), .Y (n_2058));
NAND2X1 g16528(.A (n_1332), .B (n_2842), .Y (n_2057));
AOI21X1 g16531(.A0 (n_1675), .A1 (n_2137), .B0 (n_2440), .Y (n_2056));
AOI21X1 g16542(.A0 (n_2054), .A1 (n_6796), .B0 (n_2042), .Y (n_2055));
AOI21X1 g16543(.A0 (n_7559), .A1 (n_5912), .B0 (n_231), .Y (n_2053));
AOI21X1 g16545(.A0 (n_2558), .A1 (n_6065), .B0 (n_2050), .Y (n_2052));
AOI21X1 g16546(.A0 (n_2146), .A1 (n_2000), .B0 (n_281), .Y (n_2049));
AOI21X1 g16554(.A0 (n_2046), .A1 (n_1227), .B0 (n_6801), .Y (n_2047));
NAND2X1 g16564(.A (n_1341), .B (n_2680), .Y (n_2045));
AOI21X1 g16567(.A0 (n_1629), .A1 (n_1528), .B0 (n_2136), .Y (n_2044));
AOI21X1 g16572(.A0 (n_7704), .A1 (n_2021), .B0 (n_2042), .Y (n_2043));
NAND2X1 g16574(.A (n_1331), .B (n_3049), .Y (n_2041));
AOI21X1 g16581(.A0 (n_2012), .A1 (n_2039), .B0 (n_274), .Y (n_2040));
AOI21X1 g16582(.A0 (n_998), .A1 (n_1495), .B0 (n_2036), .Y (n_2037));
AOI21X1 g16583(.A0 (n_1625), .A1 (n_2034), .B0 (n_2440), .Y (n_2035));
AOI21X1 g16587(.A0 (n_1627), .A1 (n_1591), .B0 (n_200), .Y (n_2032));
AOI21X1 g16595(.A0 (n_2015), .A1 (n_2029), .B0 (n_200), .Y (n_2030));
AOI21X1 g16603(.A0 (n_1279), .A1 (n_1603), .B0 (n_6801), .Y (n_2028));
AOI21X1 g16604(.A0 (n_1573), .A1 (n_1418), .B0 (n_1750), .Y (n_2027));
NAND2X1 g16612(.A (n_1413), .B (n_2666), .Y (n_7899));
AOI21X1 g16614(.A0 (n_2024), .A1 (n_2023), .B0 (n_2050), .Y (n_2025));
AOI21X1 g16621(.A0 (n_2021), .A1 (n_2020), .B0 (n_6801), .Y (n_2022));
AOI21X1 g16625(.A0 (n_1696), .A1 (n_2018), .B0 (n_127), .Y (n_2019));
AOI21X1 g16627(.A0 (n_2015), .A1 (n_1948), .B0 (n_2067), .Y (n_2016));
AOI21X1 g16628(.A0 (n_2146), .A1 (n_1607), .B0 (n_440), .Y (n_2014));
AOI21X1 g16637(.A0 (n_2024), .A1 (n_2012), .B0 (n_390), .Y (n_2013));
AOI21X1 g16639(.A0 (n_2010), .A1 (n_1987), .B0 (n_2440), .Y (n_2011));
NAND2X1 g16699(.A (n_1372), .B (n_1593), .Y (n_2009));
NAND2X1 g16701(.A (n_1312), .B (n_1514), .Y (n_2008));
NAND2X1 g16702(.A (n_2029), .B (n_2836), .Y (n_2007));
INVX1 g16704(.A (n_1360), .Y (n_3146));
NAND2X1 g16711(.A (n_1499), .B (n_1753), .Y (n_2004));
NAND2X1 g16719(.A (n_1435), .B (n_2374), .Y (n_2003));
NAND2X1 g16720(.A (n_2091), .B (n_2356), .Y (n_2002));
NAND2X1 g16728(.A (n_3117), .B (n_2854), .Y (n_2958));
NAND2X1 g16729(.A (n_2029), .B (n_2000), .Y (n_2001));
NAND2X1 g16733(.A (n_1372), .B (n_1670), .Y (n_2946));
INVX4 g16739(.A (n_1999), .Y (n_2981));
NAND2X1 g16746(.A (n_1997), .B (n_2174), .Y (n_1998));
NAND2X1 g16775(.A (n_2068), .B (n_2422), .Y (n_1996));
OR2X1 g16784(.A (n_1316), .B (n_1466), .Y (n_1995));
NAND2X1 g16791(.A (n_2124), .B (n_1141), .Y (n_2949));
NAND2X1 g16792(.A (n_2542), .B (n_1943), .Y (n_1994));
NAND2X1 g16795(.A (n_1312), .B (n_1629), .Y (n_1993));
NAND2X1 g16799(.A (n_2453), .B (n_6065), .Y (n_1991));
NAND2X1 g16810(.A (n_1988), .B (n_1987), .Y (n_1989));
NAND2X1 g16820(.A (n_2069), .B (n_1654), .Y (n_1986));
NAND2X1 g16823(.A (n_2854), .B (n_5924), .Y (n_1985));
OR2X1 g16826(.A (n_1065), .B (n_1286), .Y (n_1984));
NAND2X1 g16832(.A (n_1499), .B (n_2511), .Y (n_1982));
INVX1 g17843(.A (desOut[39]), .Y (n_1980));
NAND2X1 g16835(.A (n_5732), .B (n_5908), .Y (n_1979));
NAND2X1 g16844(.A (n_2521), .B (n_2124), .Y (n_1977));
NAND2X1 g16845(.A (n_1943), .B (n_2506), .Y (n_1976));
NAND2X1 g16852(.A (n_7732), .B (n_5732), .Y (n_1975));
NAND2X1 g16863(.A (n_1351), .B (n_1972), .Y (n_1974));
NAND2X1 g16866(.A (n_2456), .B (n_2012), .Y (n_1971));
NAND2X1 g16872(.A (n_2456), .B (n_2023), .Y (n_1970));
NAND2X1 g16878(.A (n_1670), .B (n_6797), .Y (n_1969));
NAND2X1 g16885(.A (n_2453), .B (n_2046), .Y (n_1968));
NAND2X1 g16889(.A (n_6058), .B (n_1629), .Y (n_1967));
NAND2X1 g16890(.A (n_2363), .B (n_1870), .Y (n_1964));
NAND2X1 g16902(.A (n_2376), .B (n_1987), .Y (n_1963));
NAND2X1 g16907(.A (n_2184), .B (n_1988), .Y (n_1962));
NAND2X1 g16913(.A (n_1711), .B (n_1598), .Y (n_1961));
NAND2X1 g16914(.A (n_5838), .B (n_6058), .Y (n_1960));
NAND2X1 g16915(.A (n_2094), .B (n_1550), .Y (n_1959));
NAND2X1 g16916(.A (n_6025), .B (n_2389), .Y (n_1958));
NAND2X1 g16917(.A (n_1358), .B (n_5908), .Y (n_1957));
NAND2X1 g16924(.A (n_2396), .B (n_5924), .Y (n_2952));
NAND2X1 g16933(.A (n_2396), .B (n_1351), .Y (n_1956));
NAND2X1 g16936(.A (n_2453), .B (n_1662), .Y (n_1955));
OR2X1 g16940(.A (n_7443), .B (n_1455), .Y (n_1954));
NAND2X1 g16946(.A (n_1997), .B (n_5732), .Y (n_1953));
NAND2X1 g16948(.A (n_2453), .B (n_999), .Y (n_1952));
NAND2X1 g16952(.A (n_3117), .B (n_6065), .Y (n_1951));
NAND2X1 g16953(.A (n_2309), .B (n_2347), .Y (n_1950));
NAND2X1 g16962(.A (n_1767), .B (n_1948), .Y (n_1949));
NAND2X1 g16965(.A (n_2935), .B (n_2374), .Y (n_1947));
NAND2X1 g16973(.A (n_2396), .B (n_953), .Y (n_2954));
NAND2X1 g16977(.A (n_1942), .B (n_2456), .Y (n_1946));
NAND2X1 g16980(.A (n_1943), .B (n_1942), .Y (n_1944));
NAND2X1 g16981(.A (n_2456), .B (n_2165), .Y (n_1941));
NAND2X1 g16983(.A (n_1381), .B (n_1351), .Y (n_1940));
NAND2X1 g16990(.A (n_1767), .B (n_2029), .Y (n_1939));
NAND2X1 g16999(.A (n_1435), .B (n_1987), .Y (n_2990));
NAND2X1 g17007(.A (n_1435), .B (n_1551), .Y (n_1937));
NAND2X1 g17009(.A (n_1670), .B (n_5908), .Y (n_1936));
NAND2X1 g16944(.A (n_2046), .B (n_1724), .Y (n_1935));
NAND2X1 g17012(.A (n_1551), .B (n_1753), .Y (n_1933));
OR2X1 g17018(.A (n_1043), .B (n_1076), .Y (n_1931));
NAND2X1 g17021(.A (n_2199), .B (n_1372), .Y (n_1930));
NAND2X1 g17026(.A (n_5838), .B (n_5924), .Y (n_1929));
NAND2X1 g17032(.A (n_2542), .B (n_2039), .Y (n_1928));
NAND2X1 g17034(.A (n_1997), .B (n_2054), .Y (n_1926));
NAND2X1 g17048(.A (n_2521), .B (n_2526), .Y (n_1924));
NAND2X1 g17063(.A (n_2389), .B (n_1658), .Y (n_1923));
NAND2X1 g17065(.A (n_2550), .B (n_2131), .Y (n_1922));
NAND2X1 g17066(.A (n_1499), .B (n_1988), .Y (n_1921));
NAND2X1 g17068(.A (n_2453), .B (n_2854), .Y (n_1920));
NAND2X1 g17071(.A (n_2550), .B (n_1918), .Y (n_1919));
NAND2X1 g17080(.A (n_1330), .B (n_2039), .Y (n_1917));
NAND2X1 g17088(.A (n_5722), .B (n_1184), .Y (n_1915));
OR2X1 g17131(.A (n_1449), .B (n_1314), .Y (n_1914));
NAND2X1 g17133(.A (n_1163), .B (n_1972), .Y (n_1913));
NAND2X1 g17135(.A (n_1943), .B (n_1330), .Y (n_1912));
INVX1 g17280(.A (n_1911), .Y (n_2793));
INVX1 g17825(.A (n_6579), .Y (desOut[63]));
CLKBUFX1 g17845(.A (n_1897), .Y (desOut[13]));
INVX1 g17846(.A (n_1897), .Y (n_1896));
INVX1 g17972(.A (desOut[61]), .Y (n_1893));
INVX2 g17866(.A (desOut[35]), .Y (n_2294));
AOI22X1 g17969(.A0 (n_1024), .A1 (n_1776), .B0 (n_3677), .B1(desIn[43]), .Y (n_2289));
NAND2X1 g17977(.A (n_743), .B (n_1277), .Y (desOut[59]));
INVX1 g17987(.A (desOut[7]), .Y (n_2286));
INVX1 g17993(.A (n_3891), .Y (desOut[29]));
NAND2X1 g15684(.A (n_1877), .B (n_2746), .Y (n_1888));
AOI21X1 g15724(.A0 (n_1142), .A1 (n_171), .B0 (n_1391), .Y (n_1887));
AOI21X1 g15725(.A0 (n_1049), .A1 (n_1861), .B0 (n_1389), .Y (n_1886));
NAND2X1 g15742(.A (n_1868), .B (n_2666), .Y (n_1884));
AOI21X1 g15754(.A0 (n_1151), .A1 (n_1882), .B0 (n_1385), .Y (n_1883));
AOI21X1 g15778(.A0 (n_1146), .A1 (n_1880), .B0 (n_1406), .Y (n_6092));
AOI21X1 g15804(.A0 (n_1153), .A1 (n_7341), .B0 (n_1382), .Y (n_1879));
NAND2X1 g15808(.A (n_6600), .B (n_1877), .Y (n_1878));
AOI21X1 g15822(.A0 (n_1150), .A1 (n_2284), .B0 (n_1402), .Y (n_1876));
AOI21X1 g15823(.A0 (n_1147), .A1 (n_7436), .B0 (n_1377), .Y (n_7903));
AOI21X1 g15824(.A0 (n_1209), .A1 (n_7301), .B0 (n_1376), .Y (n_7904));
AOI21X1 g16541(.A0 (n_7728), .A1 (n_1870), .B0 (n_274), .Y (n_1872));
NAND2X1 g15866(.A (n_1868), .B (n_2624), .Y (n_1869));
INVX1 g18506(.A (n_3677), .Y (n_3628));
INVX1 g18512(.A (n_3677), .Y (n_3673));
AOI21X1 g15877(.A0 (n_1166), .A1 (n_1861), .B0 (n_1371), .Y (n_1865));
AOI21X1 g15906(.A0 (n_1127), .A1 (n_1837), .B0 (n_1396), .Y (n_7898));
AOI21X1 g15913(.A0 (n_1068), .A1 (n_171), .B0 (n_1364), .Y (n_1863));
AOI21X1 g15929(.A0 (n_1194), .A1 (n_1861), .B0 (n_1198), .Y (n_1862));
AOI21X1 g15931(.A0 (n_1136), .A1 (n_7341), .B0 (n_1395), .Y (n_1860));
AOI21X1 g15944(.A0 (n_1838), .A1 (n_2666), .B0 (n_1411), .Y (n_1858));
AOI21X1 g15972(.A0 (n_1855), .A1 (n_2624), .B0 (n_1384), .Y (n_1856));
INVX1 g17716(.A (n_1854), .Y (n_3104));
AOI21X1 g15998(.A0 (n_2624), .A1 (n_1815), .B0 (n_1368), .Y (n_1853));
AOI21X1 g16003(.A0 (n_1851), .A1 (n_2624), .B0 (n_1365), .Y (n_1852));
AOI21X1 g16008(.A0 (n_1623), .A1 (n_1424), .B0 (n_2151), .Y (n_1850));
NAND2X1 g16013(.A (n_1423), .B (n_7301), .Y (n_1849));
AOI21X1 g16523(.A0 (n_1847), .A1 (n_1846), .B0 (n_440), .Y (n_1848));
NAND2X1 g16896(.A (n_6070), .B (n_2105), .Y (n_1843));
NAND2X1 g16080(.A (n_1788), .B (n_2668), .Y (n_1842));
NAND2X1 g16091(.A (n_1830), .B (n_2666), .Y (n_1841));
NAND2X1 g16093(.A (n_1834), .B (n_6600), .Y (n_1840));
NAND2X1 g16094(.A (n_1838), .B (n_1837), .Y (n_1839));
NAND2X1 g16095(.A (n_1805), .B (n_2746), .Y (n_1836));
NAND2X1 g16097(.A (n_1834), .B (n_2746), .Y (n_1835));
NAND2X1 g16100(.A (n_1825), .B (n_2613), .Y (n_1833));
NAND2X1 g16101(.A (n_1802), .B (n_2666), .Y (n_1832));
NAND2X1 g16102(.A (n_1830), .B (n_2624), .Y (n_1831));
NAND2X1 g16109(.A (n_1797), .B (n_2624), .Y (n_1828));
NAND2X1 g16110(.A (n_1823), .B (n_2666), .Y (n_1827));
INVX1 g18526(.A (n_3677), .Y (n_3625));
NAND2X1 g16117(.A (n_1825), .B (n_2668), .Y (n_1826));
NAND2X1 g16121(.A (n_1823), .B (n_2624), .Y (n_1824));
NAND2X1 g16123(.A (n_1808), .B (n_2666), .Y (n_1822));
INVX1 g17670(.A (n_1056), .Y (n_1821));
NAND2X1 g16128(.A (n_1795), .B (n_2666), .Y (n_1820));
NAND2X1 g16129(.A (n_1799), .B (n_2666), .Y (n_1819));
NAND2X1 g16130(.A (n_1817), .B (n_2974), .Y (n_1818));
NAND2X1 g16133(.A (n_2666), .B (n_1815), .Y (n_1816));
NAND2X1 g17039(.A (n_1691), .B (n_1724), .Y (n_1814));
CLKBUFX1 g18520(.A (n_3677), .Y (n_3668));
NAND2X1 g16142(.A (n_1811), .B (n_2746), .Y (n_1812));
NAND2X1 g16143(.A (n_1790), .B (n_2746), .Y (n_1810));
NAND2X1 g16145(.A (n_1808), .B (n_2624), .Y (n_1809));
NAND2X1 g16149(.A (n_1793), .B (n_2666), .Y (n_1807));
NAND2X1 g16155(.A (n_1805), .B (n_2668), .Y (n_1806));
NAND2X1 g16156(.A (n_1802), .B (n_2624), .Y (n_1803));
NAND2X1 g17042(.A (n_1517), .B (n_1595), .Y (n_2569));
NAND2X1 g16166(.A (n_1799), .B (n_2624), .Y (n_1800));
NAND2X1 g16167(.A (n_1797), .B (n_3179), .Y (n_1798));
NAND2X1 g16170(.A (n_1795), .B (n_2624), .Y (n_1796));
NAND2X1 g16176(.A (n_1793), .B (n_2624), .Y (n_1794));
NAND2X1 g16177(.A (n_1784), .B (n_2746), .Y (n_1792));
NAND2X1 g16182(.A (n_1790), .B (n_2216), .Y (n_1791));
NAND2X1 g16187(.A (n_1788), .B (n_2746), .Y (n_1789));
NAND2X1 g16188(.A (n_1786), .B (n_2666), .Y (n_1787));
NAND2X1 g16192(.A (n_1784), .B (n_6600), .Y (n_1785));
NAND2X1 g16216(.A (n_1169), .B (n_139), .Y (n_1783));
NAND2X1 g17079(.A (n_6025), .B (n_7559), .Y (n_1782));
AOI21X1 g16220(.A0 (n_6023), .A1 (n_2086), .B0 (n_1777), .Y (n_1779));
AOI21X1 g16235(.A0 (n_1337), .A1 (n_1052), .B0 (n_1777), .Y (n_1778));
NAND2X2 g17885(.A (n_752), .B (n_1038), .Y (desOut[37]));
NAND2X1 g17076(.A (n_1358), .B (n_2094), .Y (n_1773));
INVX1 g17877(.A (n_3709), .Y (desOut[27]));
AOI21X1 g16286(.A0 (n_1770), .A1 (n_7663), .B0 (n_7340), .Y (n_1771));
NAND2X1 g16288(.A (n_1140), .B (n_2548), .Y (n_1769));
NAND2X1 g17035(.A (n_1767), .B (n_2091), .Y (n_1768));
AOI21X1 g16298(.A0 (n_6060), .A1 (n_1374), .B0 (n_1405), .Y (n_1766));
NAND2X1 g17033(.A (n_1943), .B (n_2012), .Y (n_1764));
NAND2X1 g16319(.A (n_1004), .B (n_2548), .Y (n_1763));
AOI21X1 g16321(.A0 (n_956), .A1 (n_1681), .B0 (n_7437), .Y (n_1762));
NAND2X1 g16327(.A (n_1143), .B (n_1760), .Y (n_1761));
NAND2X1 g16329(.A (n_1051), .B (n_189), .Y (n_1759));
NAND2X1 g16332(.A (n_1053), .B (n_7436), .Y (n_1758));
NAND2X1 g16334(.A (n_1216), .B (n_2495), .Y (n_1757));
AOI21X1 g16351(.A0 (n_6025), .A1 (n_1682), .B0 (n_2440), .Y (n_1755));
AOI21X1 g16352(.A0 (n_1753), .A1 (n_2203), .B0 (n_2050), .Y (n_1754));
AOI21X1 g16365(.A0 (n_1711), .A1 (n_1682), .B0 (n_1750), .Y (n_1751));
AOI21X1 g16369(.A0 (n_1666), .A1 (n_1184), .B0 (n_2440), .Y (n_1749));
NAND2X1 g16371(.A (n_1178), .B (n_2284), .Y (n_1747));
NAND2X1 g16373(.A (n_1157), .B (n_1745), .Y (n_1746));
NAND2X1 g16374(.A (n_1167), .B (n_1880), .Y (n_1744));
NAND2X1 g16375(.A (n_1174), .B (n_7301), .Y (n_1743));
NAND2X1 g16388(.A (n_1177), .B (n_170), .Y (n_1742));
NAND2X1 g16997(.A (n_2010), .B (n_2034), .Y (n_2581));
NAND2X1 g16401(.A (n_1172), .B (n_2842), .Y (n_1740));
NAND2X1 g16994(.A (n_2091), .B (n_1572), .Y (n_1739));
AOI21X1 g16423(.A0 (n_6052), .A1 (n_1152), .B0 (n_1750), .Y (n_1738));
AOI21X1 g16460(.A0 (n_5836), .A1 (n_1600), .B0 (n_1750), .Y (n_1737));
AOI21X1 g16464(.A0 (n_1380), .A1 (n_7442), .B0 (n_2036), .Y (n_1735));
AOI21X1 g16465(.A0 (n_1918), .A1 (n_1733), .B0 (n_2050), .Y (n_1734));
NAND2X1 g16992(.A (n_1687), .B (n_2015), .Y (n_1732));
AOI21X1 g16488(.A0 (n_1770), .A1 (n_1611), .B0 (n_2440), .Y (n_1730));
INVX2 g17306(.A (n_1470), .Y (n_2340));
NAND2X1 g16517(.A (n_1145), .B (n_2284), .Y (n_1729));
NAND2X1 g17024(.A (n_998), .B (n_1727), .Y (n_1728));
NAND2X1 g16530(.A (n_1130), .B (n_2842), .Y (n_1726));
AOI21X1 g16544(.A0 (n_1374), .A1 (n_1724), .B0 (n_2440), .Y (n_1725));
NAND2X1 g16547(.A (n_1135), .B (n_171), .Y (n_1723));
AOI21X1 g16551(.A0 (n_6060), .A1 (n_6070), .B0 (n_2144), .Y (n_1722));
NAND2X1 g16553(.A (n_1212), .B (n_1719), .Y (n_1720));
NAND2X1 g16559(.A (n_1138), .B (n_7301), .Y (n_1716));
NAND2X1 g16560(.A (n_1176), .B (n_1745), .Y (n_1715));
NAND2X1 g17125(.A (n_7445), .B (n_829), .Y (n_1714));
NAND2X1 g16989(.A (n_1662), .B (n_1724), .Y (n_1713));
NAND2X2 g17851(.A (n_744), .B (n_1002), .Y (desOut[1]));
AOI21X1 g16568(.A0 (n_1711), .A1 (n_2074), .B0 (n_183), .Y (n_1712));
AOI21X1 g16596(.A0 (n_1767), .A1 (n_2541), .B0 (n_274), .Y (n_1710));
NAND2X1 g16600(.A (n_1228), .B (n_1861), .Y (n_1709));
NAND2X2 g17844(.A (n_750), .B (n_1036), .Y (desOut[39]));
INVX4 g17298(.A (n_1472), .Y (n_2882));
AOI21X1 g16609(.A0 (n_1598), .A1 (n_6796), .B0 (n_440), .Y (n_1708));
NAND2X1 g16610(.A (n_1190), .B (n_2412), .Y (n_1707));
NAND2X1 g16611(.A (n_1218), .B (n_2432), .Y (n_1706));
NAND2X1 g16613(.A (n_1129), .B (n_2842), .Y (n_1705));
AOI21X1 g16617(.A0 (n_2029), .A1 (n_1703), .B0 (n_127), .Y (n_1704));
NAND2X1 g16618(.A (n_1201), .B (n_2666), .Y (n_1702));
NAND2X1 g16622(.A (n_1034), .B (n_170), .Y (n_1701));
NAND2X1 g16630(.A (n_1148), .B (n_1719), .Y (n_1700));
NAND2X1 g16631(.A (n_1183), .B (n_1745), .Y (n_1699));
NAND2X1 g16633(.A (n_1155), .B (n_1880), .Y (n_1698));
AOI21X1 g16634(.A0 (n_1343), .A1 (n_1696), .B0 (n_200), .Y (n_1697));
NAND2X1 g16635(.A (n_1128), .B (n_2284), .Y (n_1695));
NAND2X1 g16636(.A (n_1192), .B (n_7301), .Y (n_1694));
OAI21X1 g17847(.A0 (n_934), .A1 (n_755), .B0 (n_809), .Y (n_1897));
NAND2X1 g16868(.A (n_1691), .B (n_1528), .Y (n_1692));
NAND2X1 g16836(.A (n_2034), .B (n_1591), .Y (n_1690));
NAND2X1 g16918(.A (n_6060), .B (n_1662), .Y (n_1689));
NAND2X1 g16695(.A (n_1687), .B (n_1686), .Y (n_1688));
NAND2X1 g16697(.A (n_2010), .B (n_2101), .Y (n_1685));
NAND2X1 g16714(.A (n_6567), .B (n_1682), .Y (n_1684));
NAND2X1 g16715(.A (n_1050), .B (n_1681), .Y (n_2633));
NAND2X1 g16716(.A (n_2094), .B (n_7559), .Y (n_2590));
NAND2X1 g16718(.A (n_1654), .B (n_2054), .Y (n_1680));
NAND2X1 g16724(.A (n_1662), .B (n_1312), .Y (n_1679));
NAND2X1 g16732(.A (n_7686), .B (n_1677), .Y (n_1678));
INVX2 g16740(.A (n_2245), .Y (n_1999));
NAND2X1 g16744(.A (n_2794), .B (n_1724), .Y (n_1676));
NAND2X1 g16749(.A (n_1675), .B (n_6796), .Y (n_2660));
NAND2X1 g16750(.A (n_1340), .B (n_2118), .Y (n_1673));
NAND2X1 g16776(.A (n_6796), .B (n_7559), .Y (n_1672));
NAND2X1 g16753(.A (n_1670), .B (n_2068), .Y (n_1671));
NAND2X1 g16755(.A (n_2794), .B (n_5924), .Y (n_1669));
NAND2X1 g16757(.A (n_1126), .B (n_1667), .Y (n_1668));
NAND2X1 g16758(.A (n_1666), .B (n_1508), .Y (n_2639));
NAND2X1 g16759(.A (n_2091), .B (n_1681), .Y (n_1665));
NAND2X1 g16760(.A (n_6025), .B (n_1520), .Y (n_1664));
NAND2X1 g16761(.A (n_1662), .B (n_1141), .Y (n_1663));
NAND2X1 g16762(.A (n_2199), .B (n_1660), .Y (n_1661));
NAND2X1 g16764(.A (n_2000), .B (n_1622), .Y (n_2621));
NAND2X1 g16772(.A (n_1658), .B (n_7559), .Y (n_1659));
NAND2X1 g16774(.A (n_1656), .B (n_999), .Y (n_1657));
NAND2X1 g16778(.A (n_1654), .B (n_5722), .Y (n_1655));
NAND2X1 g16779(.A (n_2101), .B (n_1651), .Y (n_1652));
NAND2X1 g16781(.A (n_1649), .B (n_1052), .Y (n_1650));
NAND2X1 g16785(.A (n_1372), .B (n_1675), .Y (n_1647));
NAND2X1 g16788(.A (n_1645), .B (n_6567), .Y (n_1646));
NAND2X1 g16789(.A (n_2311), .B (n_2541), .Y (n_1644));
NAND2X1 g16790(.A (n_1767), .B (n_2456), .Y (n_1643));
NAND2X1 g16793(.A (n_1163), .B (n_1640), .Y (n_1642));
NAND2X1 g16794(.A (n_5732), .B (n_2068), .Y (n_1639));
NAND2X1 g16802(.A (n_1343), .B (n_981), .Y (n_1638));
NAND2X1 g16803(.A (n_2015), .B (n_7685), .Y (n_1636));
NAND2X1 g16809(.A (n_1634), .B (n_1611), .Y (n_1635));
NAND2X1 g16811(.A (n_2000), .B (n_2541), .Y (n_1633));
NAND2X1 g16812(.A (n_1227), .B (n_1972), .Y (n_1632));
NAND2X1 g16813(.A (n_1380), .B (n_1629), .Y (n_1631));
NAND2X1 g16815(.A (n_1651), .B (n_1627), .Y (n_1628));
NAND2X1 g16817(.A (n_1651), .B (n_2203), .Y (n_1626));
NAND2X1 g16819(.A (n_1171), .B (n_1625), .Y (n_2619));
NAND2X1 g16821(.A (n_1623), .B (n_1622), .Y (n_1624));
OR2X1 g16825(.A (n_1292), .B (n_939), .Y (n_1621));
NAND2X1 g16827(.A (n_2124), .B (n_1619), .Y (n_1620));
NAND2X1 g16828(.A (n_2091), .B (n_1677), .Y (n_1618));
NAND2X1 g16829(.A (n_1616), .B (n_1491), .Y (n_1617));
NAND2X1 g16831(.A (n_1014), .B (n_5927), .Y (n_1615));
NAND2X1 g16833(.A (n_2165), .B (n_1355), .Y (n_1613));
NAND2X1 g16834(.A (n_964), .B (n_1622), .Y (n_1612));
NAND2X1 g16838(.A (n_2021), .B (n_1611), .Y (n_2572));
NAND2X1 g16839(.A (n_1649), .B (n_1188), .Y (n_1610));
NAND2X1 g16842(.A (n_2083), .B (n_5929), .Y (n_2631));
NAND2X1 g16843(.A (n_2456), .B (n_1607), .Y (n_1608));
NAND2X1 g16849(.A (n_1733), .B (n_7559), .Y (n_1606));
NAND2X1 g16855(.A (n_1629), .B (n_5927), .Y (n_1605));
NAND2X1 g16860(.A (n_2021), .B (n_1603), .Y (n_1604));
NAND2X1 g16861(.A (n_1258), .B (n_1870), .Y (n_1602));
NAND2X1 g16722(.A (n_1600), .B (n_1640), .Y (n_1601));
NAND2X1 g16864(.A (n_1658), .B (n_1598), .Y (n_1599));
NAND2X1 g16871(.A (n_7664), .B (n_1595), .Y (n_1597));
NAND2X1 g16875(.A (n_1593), .B (n_1733), .Y (n_1594));
NAND2X1 g16877(.A (n_2101), .B (n_1591), .Y (n_1592));
NAND2X1 g16879(.A (n_1666), .B (n_6796), .Y (n_1590));
NAND2X1 g16881(.A (n_2174), .B (n_914), .Y (n_1589));
NAND2X1 g16882(.A (n_1696), .B (n_1160), .Y (n_1587));
NAND2X1 g16883(.A (n_1660), .B (n_1670), .Y (n_1586));
NAND2X1 g16891(.A (n_1182), .B (n_1703), .Y (n_1585));
NAND2X1 g16892(.A (n_1662), .B (n_1528), .Y (n_1584));
NAND2X1 g16893(.A (n_2456), .B (n_1677), .Y (n_1583));
NAND2X1 g16897(.A (n_1870), .B (n_6796), .Y (n_1582));
NAND2X1 g16899(.A (n_5732), .B (n_1658), .Y (n_1580));
NAND2X1 g16900(.A (n_1578), .B (n_2183), .Y (n_1579));
NAND2X1 g16904(.A (n_999), .B (n_5924), .Y (n_1577));
NAND2X1 g16909(.A (n_1753), .B (n_1987), .Y (n_1576));
NAND2X1 g16910(.A (n_1703), .B (n_981), .Y (n_1575));
NAND2X1 g16911(.A (n_1573), .B (n_1572), .Y (n_1574));
NAND2X1 g16912(.A (n_7581), .B (n_7445), .Y (n_2584));
NAND2X1 g16919(.A (n_7637), .B (n_2021), .Y (n_1571));
NAND2X1 g16920(.A (n_6567), .B (n_1666), .Y (n_2657));
NAND2X1 g16921(.A (n_1675), .B (n_1184), .Y (n_1570));
NAND2X1 g16925(.A (n_1660), .B (n_1388), .Y (n_2586));
NAND2X1 g16926(.A (n_2174), .B (n_1658), .Y (n_2592));
NAND2X1 g16929(.A (n_2124), .B (n_1724), .Y (n_1568));
NAND2X1 g16930(.A (n_1152), .B (n_1619), .Y (n_2604));
NAND2X1 g16931(.A (n_1168), .B (n_1645), .Y (n_1567));
NAND2X1 g16932(.A (n_1358), .B (n_1654), .Y (n_1566));
NAND2X1 g16935(.A (n_1687), .B (n_2018), .Y (n_1564));
NAND2X1 g16938(.A (n_1651), .B (n_1562), .Y (n_1563));
NAND2X1 g16947(.A (n_1670), .B (n_7732), .Y (n_1561));
NAND2X1 g16950(.A (n_5912), .B (n_1682), .Y (n_1560));
NAND2X1 g16954(.A (n_964), .B (n_7685), .Y (n_2596));
NAND2X1 g16957(.A (n_2000), .B (n_7686), .Y (n_1556));
NAND2X1 g16958(.A (n_6963), .B (n_2094), .Y (n_1554));
NAND2X1 g16959(.A (n_2086), .B (n_5908), .Y (n_1553));
NAND2X1 g16960(.A (n_1551), .B (n_1533), .Y (n_1552));
NAND2X1 g16967(.A (n_1660), .B (n_1550), .Y (n_2598));
NAND2X1 g16969(.A (n_1325), .B (n_1064), .Y (n_1549));
NAND2X1 g16970(.A (n_1358), .B (n_6022), .Y (n_1548));
NAND2X1 g16974(.A (n_6963), .B (n_6567), .Y (n_2588));
NAND2X1 g16975(.A (n_1562), .B (n_1310), .Y (n_1545));
NAND2X1 g16979(.A (n_1543), .B (n_1595), .Y (n_1544));
OR2X1 g16985(.A (n_1284), .B (n_1541), .Y (n_1542));
NAND2X1 g16986(.A (n_2074), .B (n_1258), .Y (n_1540));
NAND2X1 g16991(.A (n_1538), .B (n_1041), .Y (n_1539));
NAND2X1 g17000(.A (n_1619), .B (n_1629), .Y (n_1537));
NAND2X1 g17004(.A (n_1649), .B (n_2183), .Y (n_1536));
NAND2X1 g17014(.A (n_937), .B (n_1533), .Y (n_1534));
NAND2X1 g17015(.A (n_1662), .B (n_1600), .Y (n_1532));
NAND2X1 g17017(.A (n_1227), .B (n_1691), .Y (n_1531));
NAND2X1 g17019(.A (n_7442), .B (n_1528), .Y (n_1530));
NAND2X1 g17031(.A (n_6567), .B (n_1346), .Y (n_1527));
NAND2X1 g17040(.A (n_2124), .B (n_2105), .Y (n_1526));
NAND2X1 g17043(.A (n_922), .B (n_1485), .Y (n_2616));
NAND2X1 g17044(.A (n_7442), .B (n_5929), .Y (n_1525));
NAND2X1 g17047(.A (n_2100), .B (n_2034), .Y (n_1523));
NAND2X1 g17049(.A (n_7446), .B (n_2083), .Y (n_1522));
NAND2X1 g17050(.A (n_2137), .B (n_1520), .Y (n_1521));
NAND2X1 g17051(.A (n_1667), .B (n_1134), .Y (n_1519));
NAND2X1 g17052(.A (n_1517), .B (n_2180), .Y (n_1518));
NAND2X1 g17053(.A (n_1572), .B (n_1064), .Y (n_2629));
NAND2X1 g17056(.A (n_2183), .B (n_1562), .Y (n_2614));
NAND2X1 g17057(.A (n_5912), .B (n_1550), .Y (n_1516));
NAND2X1 g17058(.A (n_2105), .B (n_1514), .Y (n_1515));
NAND2X1 g17059(.A (n_1675), .B (n_5921), .Y (n_1513));
NAND2X1 g17060(.A (n_1141), .B (n_1972), .Y (n_1512));
NAND2X1 g17061(.A (n_1381), .B (n_1141), .Y (n_1510));
NAND2X1 g17062(.A (n_1508), .B (n_1682), .Y (n_1509));
NAND2X1 g17064(.A (n_1381), .B (n_1619), .Y (n_1507));
NAND2X1 g17067(.A (n_1374), .B (n_1312), .Y (n_1506));
NAND2X1 g17073(.A (n_829), .B (n_789), .Y (n_2594));
NAND2X1 g17083(.A (n_2078), .B (n_1141), .Y (n_2579));
NAND2X1 g17087(.A (n_1543), .B (n_2100), .Y (n_1502));
NAND2X1 g17092(.A (n_1703), .B (n_1064), .Y (n_1501));
NAND2X1 g17094(.A (n_6058), .B (n_1514), .Y (n_2577));
NAND2X1 g17095(.A (n_1215), .B (n_1499), .Y (n_1500));
NAND2X1 g17096(.A (n_7686), .B (n_1681), .Y (n_1498));
NAND2X1 g17097(.A (n_2083), .B (n_1656), .Y (n_1497));
NAND2X1 g17103(.A (n_1623), .B (n_1495), .Y (n_1496));
NAND2X1 g17111(.A (n_1517), .B (n_1233), .Y (n_2611));
NAND2X1 g17114(.A (n_1428), .B (n_5912), .Y (n_2575));
NAND2X1 g17116(.A (n_921), .B (n_1640), .Y (n_2626));
NAND2X1 g17118(.A (n_2091), .B (n_1491), .Y (n_1493));
NAND2X1 g17119(.A (n_1616), .B (n_1418), .Y (n_1490));
NAND2X1 g17120(.A (n_7682), .B (n_1538), .Y (n_1489));
NAND2X1 g17122(.A (n_1662), .B (n_1619), .Y (n_1488));
NAND2X1 g17126(.A (n_2091), .B (n_1686), .Y (n_1487));
NAND2X1 g17127(.A (n_1616), .B (n_1485), .Y (n_1486));
NAND2X1 g17134(.A (n_6800), .B (n_5908), .Y (n_1484));
NAND2X1 g17138(.A (n_1846), .B (n_2178), .Y (n_1482));
INVX1 g17156(.A (n_2376), .Y (n_1481));
CLKBUFX1 g17994(.A (n_1480), .Y (n_3891));
INVX1 g17282(.A (n_1312), .Y (n_1911));
INVX1 g17995(.A (n_1480), .Y (n_1478));
NAND2X1 g16846(.A (n_7445), .B (n_1629), .Y (n_1475));
INVX1 g17419(.A (n_1466), .Y (n_2830));
INVX1 g17484(.A (n_1464), .Y (n_1465));
INVX2 g17485(.A (n_1464), .Y (n_2839));
INVX1 g17516(.A (n_1459), .Y (n_2888));
INVX1 g17601(.A (n_1070), .Y (n_2879));
INVX1 g17651(.A (n_1455), .Y (n_1454));
INVX1 g17671(.A (n_1056), .Y (n_2366));
INVX1 g17717(.A (n_1629), .Y (n_1854));
AOI21X1 g17980(.A0 (n_826), .A1 (n_925), .B0 (n_3677), .Y (n_1445));
NAND2X1 g16561(.A (n_1164), .B (n_1880), .Y (n_1443));
NAND2X1 g16869(.A (n_1520), .B (n_1508), .Y (n_1442));
OAI21X1 g17874(.A0 (n_942), .A1 (n_3677), .B0 (n_898), .Y(desOut[45]));
INVX1 g17812(.A (n_3585), .Y (desOut[31]));
INVX1 g17794(.A (n_1948), .Y (n_1885));
INVX2 g17498(.A (n_1437), .Y (n_2806));
INVX1 g17730(.A (n_1942), .Y (n_1902));
AOI21X1 g16297(.A0 (n_1435), .A1 (n_1627), .B0 (n_198), .Y (n_1436));
NAND2X1 g17104(.A (n_1696), .B (n_1035), .Y (n_1433));
NAND2X1 g17008(.A (n_1660), .B (n_1428), .Y (n_1429));
INVX1 g17722(.A (n_1449), .Y (n_2330));
NAND2X1 g17046(.A (n_1847), .B (n_2101), .Y (n_1427));
NAND2X1 g16078(.A (n_1424), .B (n_1160), .Y (n_1877));
NAND2X1 g16112(.A (n_1424), .B (n_1681), .Y (n_1423));
INVX1 g17392(.A (n_1422), .Y (n_2319));
NAND2X1 g16164(.A (n_1703), .B (n_1424), .Y (n_1868));
NAND2X1 g16165(.A (n_1419), .B (n_2746), .Y (n_1420));
NAND2X1 g17085(.A (n_963), .B (n_1418), .Y (n_2214));
INVX1 g17652(.A (n_2105), .Y (n_1455));
NAND2X1 g16184(.A (n_1415), .B (n_2746), .Y (n_1416));
NAND2X1 g16185(.A (n_1485), .B (n_1424), .Y (n_1414));
NAND2X1 g17084(.A (n_1343), .B (n_7702), .Y (n_1413));
AOI21X1 g16218(.A0 (n_914), .A1 (n_1339), .B0 (n_7340), .Y (n_1411));
AOI21X1 g16221(.A0 (n_1703), .A1 (n_1495), .B0 (n_7340), .Y (n_1409));
AOI21X1 g16241(.A0 (n_1380), .A1 (n_6070), .B0 (n_7437), .Y (n_1408));
AOI21X1 g16256(.A0 (n_7685), .A1 (n_1397), .B0 (n_1405), .Y (n_1406));
INVX2 g17368(.A (n_1403), .Y (n_2396));
INVX1 g17364(.A (n_1403), .Y (n_1404));
AOI21X1 g16276(.A0 (n_1171), .A1 (n_1154), .B0 (n_1405), .Y (n_1402));
INVX1 g17360(.A (n_1399), .Y (n_2526));
AOI21X1 g16320(.A0 (n_1696), .A1 (n_1397), .B0 (n_191), .Y (n_1398));
AOI21X1 g16324(.A0 (n_1622), .A1 (n_1681), .B0 (n_7340), .Y (n_1396));
AOI21X1 g16337(.A0 (n_1622), .A1 (n_1200), .B0 (n_1750), .Y (n_1395));
AOI21X1 g16370(.A0 (n_7704), .A1 (n_1188), .B0 (n_316), .Y (n_1393));
AOI21X1 g16379(.A0 (n_7354), .A1 (n_999), .B0 (n_6801), .Y (n_1391));
AOI21X1 g16408(.A0 (n_7700), .A1 (n_1181), .B0 (n_274), .Y (n_1390));
AOI21X1 g16409(.A0 (n_1388), .A1 (n_5912), .B0 (n_2440), .Y (n_1389));
AOI21X1 g16417(.A0 (n_6070), .A1 (n_1724), .B0 (n_1750), .Y (n_1387));
AOI21X1 g16420(.A0 (n_7634), .A1 (n_2020), .B0 (n_2144), .Y (n_1385));
CLKBUFX3 g17321(.A (n_1491), .Y (n_2836));
AOI21X1 g16470(.A0 (n_7733), .A1 (n_7700), .B0 (n_2144), .Y (n_1384));
AOI21X1 g16471(.A0 (n_1381), .A1 (n_1380), .B0 (n_2248), .Y (n_1382));
AOI21X1 g16473(.A0 (n_6963), .A1 (n_6759), .B0 (n_1750), .Y (n_1379));
AOI21X1 g16489(.A0 (n_1366), .A1 (n_7704), .B0 (n_127), .Y (n_1377));
AOI21X1 g16492(.A0 (n_1696), .A1 (n_1170), .B0 (n_207), .Y (n_1376));
AOI21X1 g16521(.A0 (n_1600), .A1 (n_1374), .B0 (n_6801), .Y (n_1375));
NAND2X1 g16928(.A (n_1372), .B (n_1682), .Y (n_1373));
AOI21X1 g16569(.A0 (n_7700), .A1 (n_979), .B0 (n_2248), .Y (n_1371));
AOI21X1 g16570(.A0 (n_6060), .A1 (n_972), .B0 (n_6801), .Y (n_1370));
NAND2X1 g16593(.A (n_970), .B (n_2624), .Y (n_1369));
AOI21X1 g16601(.A0 (n_2020), .A1 (n_1144), .B0 (n_2440), .Y (n_1368));
AOI21X1 g16607(.A0 (n_1366), .A1 (n_1543), .B0 (n_2440), .Y (n_1367));
AOI21X1 g16619(.A0 (n_1572), .A1 (n_1355), .B0 (n_2248), .Y (n_1365));
AOI21X1 g16620(.A0 (n_1538), .A1 (n_1667), .B0 (n_2144), .Y (n_1364));
AOI21X1 g16623(.A0 (n_1052), .A1 (n_1603), .B0 (n_1750), .Y (n_1363));
NAND2X1 g16984(.A (n_1543), .B (n_1052), .Y (n_1362));
INVX1 g16707(.A (n_1360), .Y (n_2250));
INVX1 g16708(.A (n_1360), .Y (n_1361));
NAND2X1 g16780(.A (n_1358), .B (n_1184), .Y (n_1359));
NAND2X1 g16725(.A (n_1770), .B (n_1603), .Y (n_2207));
NAND2X1 g16731(.A (n_1677), .B (n_1355), .Y (n_1356));
INVX4 g16741(.A (n_1353), .Y (n_2245));
NAND2X1 g16745(.A (n_1351), .B (n_1158), .Y (n_1352));
NAND2X1 g16747(.A (n_6027), .B (n_5732), .Y (n_1350));
NAND2X1 g16748(.A (n_5836), .B (n_967), .Y (n_2228));
NAND2X1 g16763(.A (n_951), .B (n_1603), .Y (n_1348));
NAND2X1 g16771(.A (n_988), .B (n_1346), .Y (n_1347));
OAI21X1 g18083(.A0 (n_880), .A1 (n_733), .B0 (n_878), .Y (n_1345));
NAND2X1 g16801(.A (n_1343), .B (n_2029), .Y (n_1344));
NAND2X1 g16807(.A (n_1343), .B (n_1355), .Y (n_2221));
NAND2X1 g16886(.A (n_1351), .B (n_6070), .Y (n_2217));
NAND2X1 g16818(.A (n_980), .B (n_1329), .Y (n_1341));
NAND2X1 g16858(.A (n_1340), .B (n_1625), .Y (n_2236));
NAND2X1 g16837(.A (n_794), .B (n_1339), .Y (n_2257));
NAND2X1 g16848(.A (n_1366), .B (n_1667), .Y (n_2233));
NAND2X1 g16851(.A (n_951), .B (n_1337), .Y (n_1338));
NAND2X1 g16859(.A (n_6027), .B (n_2074), .Y (n_1336));
NAND2X1 g16865(.A (n_951), .B (n_1667), .Y (n_2205));
NAND2X1 g16884(.A (n_7700), .B (n_1372), .Y (n_1335));
NAND2X1 g16768(.A (n_5835), .B (n_1351), .Y (n_1334));
NAND2X1 g17128(.A (n_1340), .B (n_1634), .Y (n_1332));
NAND2X1 g16903(.A (n_1330), .B (n_1355), .Y (n_1331));
NAND2X1 g16906(.A (n_1329), .B (n_1724), .Y (n_2219));
NAND2X1 g16923(.A (n_1163), .B (n_971), .Y (n_1328));
NAND2X1 g16982(.A (n_7664), .B (n_1052), .Y (n_1327));
NAND2X1 g16942(.A (n_1325), .B (n_963), .Y (n_1326));
NAND2X1 g16987(.A (n_1770), .B (n_1340), .Y (n_1324));
NAND2X1 g17003(.A (n_1099), .B (n_1156), .Y (n_1323));
NAND2X1 g17069(.A (n_1358), .B (n_6796), .Y (n_2238));
NAND2X1 g17072(.A (n_1325), .B (n_1696), .Y (n_1322));
NAND2X1 g17101(.A (n_7701), .B (n_914), .Y (n_1321));
NAND2X1 g17115(.A (n_1770), .B (n_937), .Y (n_1320));
NAND2X1 g17117(.A (n_1325), .B (n_1355), .Y (n_1319));
NAND2X1 g16796(.A (n_2074), .B (n_2068), .Y (n_1317));
CLKBUFX3 g17157(.A (n_1595), .Y (n_2376));
CLKBUFX3 g17214(.A (n_2023), .Y (n_2838));
AOI21X1 g17996(.A0 (n_753), .A1 (n_1469), .B0 (n_927), .Y (n_1480));
CLKBUFX1 g17247(.A (n_1593), .Y (n_2329));
NAND2X1 g16756(.A (n_1351), .B (n_1329), .Y (n_1311));
INVX2 g17299(.A (n_1972), .Y (n_1472));
INVX2 g17308(.A (n_2180), .Y (n_1470));
INVX2 g17335(.A (n_1305), .Y (n_2542));
INVX1 g17387(.A (n_1302), .Y (n_2309));
CLKBUFX3 g17413(.A (n_1514), .Y (n_2557));
INVX1 g17429(.A (n_1300), .Y (n_3117));
CLKBUFX1 g17439(.A (n_1649), .Y (n_2895));
CLKBUFX1 g17446(.A (n_1623), .Y (n_2356));
INVX2 g17499(.A (n_1686), .Y (n_1437));
CLKBUFX1 g17543(.A (n_1562), .Y (n_2374));
INVX2 g17589(.A (n_1378), .Y (n_2453));
CLKBUFX3 g17595(.A (n_1607), .Y (n_2506));
CLKBUFX3 g17614(.A (n_1691), .Y (n_2499));
NAND3X1 g17985(.A (n_923), .B (n_810), .C (n_758), .Y (n_1294));
INVX2 g17534(.A (n_1291), .Y (n_2854));
NAND3X1 g17984(.A (n_825), .B (n_720), .C (n_821), .Y (n_1290));
CLKBUFX1 g17697(.A (n_1660), .Y (n_1997));
CLKBUFX3 g17711(.A (n_1508), .Y (n_2503));
INVX4 g17731(.A (n_1251), .Y (n_1942));
INVX1 g17753(.A (n_1284), .Y (n_2511));
CLKBUFX3 g17758(.A (n_1428), .Y (n_2389));
INVX2 g17783(.A (n_1264), .Y (n_2550));
INVX1 g17805(.A (n_1272), .Y (n_2521));
INVX1 g17829(.A (n_7021), .Y (desOut[33]));
NAND2X1 g17054(.A (n_1372), .B (n_1349), .Y (n_2212));
NOR2X1 g17878(.A (n_725), .B (n_931), .Y (n_3709));
NAND2X1 g17112(.A (n_1343), .B (n_1193), .Y (n_1281));
INVX1 g17518(.A (n_2060), .Y (n_1459));
AOI21X1 g16615(.A0 (n_1517), .A1 (n_1279), .B0 (n_440), .Y (n_1280));
NAND2X1 g17979(.A (n_973), .B (n_879), .Y (n_1277));
NAND3X1 g17981(.A (n_822), .B (n_721), .C (n_908), .Y (n_1276));
AOI22X1 g17813(.A0 (n_909), .A1 (n_559), .B0 (n_701), .B1(desIn[31]), .Y (n_3585));
MX2X1 g18055(.A (FP_R_21), .B (n_812), .S0 (n_1268), .Y (n_1271));
CLKBUFX3 g17800(.A (n_1533), .Y (n_1988));
INVX1 g17508(.A (n_932), .Y (n_2408));
MX2X1 g18068(.A (FP_R_5), .B (n_874), .S0 (n_1268), .Y (n_1269));
AOI22X1 g18069(.A0 (n_811), .A1 (n_733), .B0 (n_3550), .B1 (FP_R_29),.Y (n_1267));
INVX2 g17486(.A (n_1573), .Y (n_1464));
NAND2X1 g17028(.A (n_1258), .B (n_1550), .Y (n_1259));
NAND2X1 g16976(.A (n_1770), .B (n_1517), .Y (n_1255));
INVX2 g17746(.A (n_1253), .Y (n_2422));
INVX2 g17456(.A (n_1256), .Y (n_2363));
INVX1 g17724(.A (n_2068), .Y (n_1449));
INVX1 g17420(.A (n_1591), .Y (n_1466));
MX2X1 g16051(.A (L_91), .B (FP_R_60), .S0 (n_7846), .Y (n_1241));
INVX2 g16742(.A (n_962), .Y (n_1353));
INVX4 g17406(.A (n_1237), .Y (n_1662));
INVX2 g17678(.A (n_1221), .Y (n_7682));
INVX1 g17172(.A (n_1499), .Y (n_1316));
INVX1 g17397(.A (n_1232), .Y (n_1233));
INVX4 g17653(.A (n_1229), .Y (n_2105));
INVX2 g17640(.A (n_1061), .Y (n_2794));
NAND2X1 g17036(.A (n_1366), .B (n_1041), .Y (n_1228));
INVX2 g17648(.A (n_1229), .Y (n_1227));
INVX2 g17643(.A (n_1225), .Y (n_2165));
INVX2 g17634(.A (n_1063), .Y (n_1616));
INVX2 g17679(.A (n_1221), .Y (n_2101));
CLKBUFX3 g17353(.A (n_1634), .Y (n_2935));
AOI21X1 g16309(.A0 (n_1180), .A1 (n_1346), .B0 (n_7340), .Y (n_1219));
NAND2X1 g17077(.A (n_1543), .B (n_1625), .Y (n_1218));
INVX4 g17300(.A (n_1103), .Y (n_1972));
NAND2X1 g17132(.A (n_1215), .B (n_7705), .Y (n_1216));
INVX1 g17618(.A (n_1213), .Y (n_7581));
NAND2X1 g17074(.A (n_6963), .B (n_1184), .Y (n_1212));
INVX1 g17336(.A (n_1325), .Y (n_1305));
NAND2X1 g16968(.A (n_1517), .B (n_1538), .Y (n_1209));
INVX1 g17591(.A (n_921), .Y (n_1378));
INVX1 g17322(.A (n_1206), .Y (n_1491));
INVX2 g17596(.A (n_1071), .Y (n_1607));
NAND2X1 g17978(.A (n_827), .B (n_879), .Y (n_1208));
INVX1 g17320(.A (n_1206), .Y (n_2012));
INVX2 g17158(.A (n_1125), .Y (n_1595));
INVX2 g17584(.A (n_1204), .Y (n_1654));
CLKBUFX1 g17424(.A (n_1340), .Y (n_2184));
INVX2 g17303(.A (n_1102), .Y (n_2021));
NAND2X1 g17020(.A (n_1538), .B (n_1543), .Y (n_2649));
NAND2X1 g16988(.A (n_1687), .B (n_1200), .Y (n_1201));
INVX1 g17167(.A (n_1195), .Y (n_2558));
AOI21X1 g16624(.A0 (n_1681), .A1 (n_1355), .B0 (n_6801), .Y (n_1198));
INVX1 g17389(.A (n_1184), .Y (n_1302));
NAND2X1 g16734(.A (n_7702), .B (n_1418), .Y (n_1194));
NAND2X1 g16765(.A (n_966), .B (n_1193), .Y (n_1784));
INVX4 g17312(.A (n_1100), .Y (n_1645));
NAND2X1 g16700(.A (n_7636), .B (n_7634), .Y (n_1192));
NAND2X1 g16703(.A (n_1215), .B (n_1667), .Y (n_1190));
INVX2 g16709(.A (n_1424), .Y (n_1360));
NAND2X1 g16712(.A (n_1182), .B (n_1397), .Y (n_1786));
NAND2X1 g16713(.A (n_7663), .B (n_1188), .Y (n_1788));
NAND2X1 g16726(.A (n_1149), .B (n_981), .Y (n_1851));
NAND2X1 g16730(.A (n_947), .B (n_1184), .Y (n_1811));
NAND2X1 g16735(.A (n_7632), .B (n_1182), .Y (n_1183));
NAND2X1 g16887(.A (n_2074), .B (n_1181), .Y (n_1795));
NAND2X1 g16766(.A (n_6963), .B (n_1180), .Y (n_1838));
NAND2X1 g16769(.A (n_7733), .B (n_1550), .Y (n_1808));
NAND2X1 g16770(.A (n_889), .B (n_1162), .Y (n_1178));
NAND2X1 g16777(.A (n_7663), .B (n_1279), .Y (n_1177));
NAND2X1 g16773(.A (n_1381), .B (n_953), .Y (n_1805));
NAND2X1 g16782(.A (n_6759), .B (n_1173), .Y (n_1176));
NAND2X1 g16797(.A (n_926), .B (n_1173), .Y (n_1174));
NAND2X1 g16798(.A (n_1366), .B (n_1171), .Y (n_1172));
NAND2X1 g16808(.A (n_1170), .B (n_1355), .Y (n_1823));
NAND2X1 g16816(.A (n_918), .B (n_1168), .Y (n_1169));
NAND2X1 g16830(.A (n_1168), .B (n_1388), .Y (n_1825));
NAND2X1 g16841(.A (n_7701), .B (n_794), .Y (n_1167));
NAND2X1 g16847(.A (n_1380), .B (n_1374), .Y (n_1166));
NAND2X1 g16853(.A (n_1163), .B (n_1162), .Y (n_1164));
NAND2X1 g16854(.A (n_7685), .B (n_1160), .Y (n_1161));
NAND2X1 g16873(.A (n_6053), .B (n_1158), .Y (n_1855));
NAND2X1 g16874(.A (n_5836), .B (n_1380), .Y (n_1157));
NAND2X1 g16895(.A (n_1381), .B (n_1156), .Y (n_1799));
NAND2X1 g16905(.A (n_7733), .B (n_1346), .Y (n_1817));
NAND2X1 g17129(.A (n_7663), .B (n_1154), .Y (n_1155));
NAND2X1 g16934(.A (n_1163), .B (n_1152), .Y (n_1153));
NAND2X1 g16949(.A (n_7705), .B (n_1279), .Y (n_1151));
NAND2X1 g16955(.A (n_1149), .B (n_1182), .Y (n_1150));
NAND2X1 g16956(.A (n_1050), .B (n_964), .Y (n_1148));
NAND2X1 g16961(.A (n_1215), .B (n_1337), .Y (n_1147));
NAND2X1 g16880(.A (n_1485), .B (n_7702), .Y (n_1146));
NAND2X1 g16876(.A (n_1611), .B (n_1144), .Y (n_1145));
NAND2X1 g16995(.A (n_1696), .B (n_1485), .Y (n_1143));
NAND2X1 g17001(.A (n_1141), .B (n_1374), .Y (n_1142));
NAND2X1 g17002(.A (n_1611), .B (n_1279), .Y (n_1140));
NAND2X1 g17006(.A (n_1366), .B (n_7664), .Y (n_1139));
NAND2X1 g17011(.A (n_1380), .B (n_1152), .Y (n_1138));
NAND2X1 g17016(.A (n_5732), .B (n_6796), .Y (n_1137));
NAND2X1 g17025(.A (n_1188), .B (n_1603), .Y (n_1136));
NAND2X1 g17037(.A (n_921), .B (n_7440), .Y (n_1834));
NAND2X1 g17038(.A (n_7445), .B (n_1374), .Y (n_1830));
INVX2 g17568(.A (n_1075), .Y (n_2183));
NAND2X1 g17055(.A (n_7664), .B (n_1134), .Y (n_1135));
NAND2X1 g17078(.A (n_1325), .B (n_7686), .Y (n_1797));
NAND2X1 g17099(.A (n_1337), .B (n_1144), .Y (n_1793));
NAND2X1 g16850(.A (n_1696), .B (n_1681), .Y (n_1802));
NAND2X1 g17105(.A (n_1366), .B (n_1517), .Y (n_1133));
NAND2X1 g17113(.A (n_1170), .B (n_1622), .Y (n_1132));
NAND2X1 g17121(.A (n_7636), .B (n_7655), .Y (n_1790));
NAND2X1 g17123(.A (n_7634), .B (n_1337), .Y (n_1130));
NAND2X1 g16941(.A (n_1611), .B (n_1188), .Y (n_1129));
NAND2X1 g17130(.A (n_1170), .B (n_922), .Y (n_1128));
NAND2X1 g17137(.A (n_1687), .B (n_1200), .Y (n_1127));
INVX1 g17159(.A (n_1125), .Y (n_1126));
CLKBUFX3 g17162(.A (n_1677), .Y (n_2311));
INVX2 g17215(.A (n_1116), .Y (n_2023));
INVX4 g17284(.A (n_1115), .Y (n_1312));
INVX1 g17246(.A (n_1113), .Y (n_1870));
INVX2 g17292(.A (n_1104), .Y (n_1310));
CLKBUFX3 g17263(.A (n_2086), .Y (n_2054));
INVX2 g17277(.A (n_1093), .Y (n_1670));
INVX2 g17544(.A (n_1106), .Y (n_1562));
INVX1 g17293(.A (n_1104), .Y (n_2178));
INVX2 g17309(.A (n_1102), .Y (n_2180));
INVX1 g17361(.A (n_2046), .Y (n_1399));
INVX1 g17369(.A (n_1099), .Y (n_1403));
CLKBUFX1 g17376(.A (n_1770), .Y (n_1847));
INVX1 g17393(.A (n_7664), .Y (n_1422));
INVX2 g17401(.A (n_1232), .Y (n_2118));
INVX2 g17414(.A (n_1094), .Y (n_1514));
INVX1 g17275(.A (n_1093), .Y (n_1520));
INVX2 g17421(.A (n_983), .Y (n_1591));
INVX4 g17243(.A (n_1013), .Y (n_2124));
INVX4 g17462(.A (n_1088), .Y (n_2094));
INVX4 g17487(.A (n_1085), .Y (n_1573));
INVX1 g17504(.A (n_1082), .Y (n_2347));
INVX2 g17514(.A (n_1081), .Y (n_2015));
INVX2 g17519(.A (n_1081), .Y (n_2060));
INVX1 g17535(.A (n_1374), .Y (n_1291));
INVX2 g17559(.A (n_1076), .Y (n_1846));
INVX4 g17603(.A (n_1070), .Y (n_2137));
NAND2X1 g16894(.A (n_1171), .B (n_7655), .Y (n_1068));
INVX1 g17615(.A (n_1213), .Y (n_1691));
INVX2 g17617(.A (n_1213), .Y (n_1640));
INVX1 g17628(.A (n_1063), .Y (n_1064));
INVX1 g17657(.A (n_1435), .Y (n_1292));
INVX2 g17673(.A (n_1056), .Y (n_1727));
INVX4 g17685(.A (n_1054), .Y (n_2034));
NAND2X1 g16698(.A (n_1171), .B (n_1052), .Y (n_1053));
INVX1 g17701(.A (n_990), .Y (n_2069));
NAND2X1 g17091(.A (n_1050), .B (n_1572), .Y (n_1051));
INVX1 g17710(.A (n_996), .Y (n_1658));
INVX2 g17719(.A (n_993), .Y (n_1629));
INVX2 g17733(.A (n_1343), .Y (n_1251));
NAND2X1 g16694(.A (n_1158), .B (n_5927), .Y (n_1049));
INVX1 g17749(.A (n_1550), .Y (n_1253));
INVX2 g17764(.A (n_1047), .Y (n_2000));
INVX4 g17272(.A (n_1107), .Y (n_1528));
INVX4 g17771(.A (n_1046), .Y (n_2091));
INVX2 g17787(.A (n_1372), .Y (n_1264));
INVX1 g17792(.A (n_1028), .Y (n_2024));
INVX1 g17801(.A (n_1033), .Y (n_1533));
INVX1 g17807(.A (n_1380), .Y (n_1272));
NAND2X1 g17108(.A (n_1052), .B (n_1041), .Y (n_1815));
INVX2 g17314(.A (n_1100), .Y (n_2174));
NAND2X1 g17924(.A (n_838), .B (n_559), .Y (n_1038));
NAND2X1 g17931(.A (n_837), .B (n_559), .Y (n_1036));
INVX1 g17515(.A (n_1081), .Y (n_1035));
INVX4 g17776(.A (n_1043), .Y (n_2010));
NAND2X1 g16786(.A (n_1170), .B (n_7686), .Y (n_1034));
INVX1 g17254(.A (n_1109), .Y (n_1651));
INVX1 g17799(.A (n_1033), .Y (n_2100));
INVX2 g17500(.A (n_1031), .Y (n_1686));
MX2X1 g18059(.A (n_736), .B (FP_R_13), .S0 (n_3550), .Y (n_1030));
INVX2 g17796(.A (n_1028), .Y (n_1948));
AOI22X1 g18053(.A0 (n_728), .A1 (n_733), .B0 (n_610), .B1 (FP_R_6),.Y (n_1027));
MX2X1 g18066(.A (FP_R_26), .B (n_737), .S0 (n_714), .Y (n_1026));
OAI21X1 g18085(.A0 (n_772), .A1 (n_714), .B0 (n_751), .Y (n_1025));
OR2X1 g18089(.A (n_796), .B (n_765), .Y (n_1024));
INVX1 g17248(.A (n_1113), .Y (n_1593));
NAND2X1 g17941(.A (n_834), .B (n_559), .Y (n_1018));
INVX1 g17754(.A (n_1052), .Y (n_1284));
INVX2 g17480(.A (n_1015), .Y (n_1551));
INVX1 g17241(.A (n_1013), .Y (n_1014));
INVX2 g17759(.A (n_1007), .Y (n_1428));
INVX2 g17757(.A (n_1007), .Y (n_1675));
INVX2 g17468(.A (n_1005), .Y (n_2083));
NAND2X1 g16937(.A (n_7664), .B (n_1625), .Y (n_1004));
NAND2X1 g17927(.A (n_801), .B (n_559), .Y (n_1003));
NAND2X1 g17926(.A (n_833), .B (n_559), .Y (n_1002));
NAND2X1 g17102(.A (n_1380), .B (n_999), .Y (n_2671));
INVX2 g17457(.A (n_1711), .Y (n_1256));
INVX2 g17216(.A (n_1116), .Y (n_998));
INVX2 g17447(.A (n_1089), .Y (n_1623));
INVX1 g17448(.A (n_1089), .Y (n_2018));
INVX2 g17712(.A (n_996), .Y (n_1508));
INVX4 g17440(.A (n_995), .Y (n_1649));
INVX1 g17210(.A (n_2131), .Y (n_1314));
INVX1 g17715(.A (n_993), .Y (n_2078));
INVX4 g17434(.A (n_992), .Y (n_2456));
INVX1 g17430(.A (n_1163), .Y (n_1300));
INVX1 g17707(.A (n_1330), .Y (n_1286));
INVX4 g17186(.A (n_997), .Y (n_1619));
INVX4 g18378(.A (n_3550), .Y (n_1260));
CLKBUFX3 g17698(.A (n_988), .Y (n_1660));
NAND2X1 g17093(.A (n_1687), .B (n_1572), .Y (n_985));
INVX4 g17330(.A (n_968), .Y (n_1351));
INVX2 g17408(.A (n_1162), .Y (n_1237));
INVX2 g17402(.A (n_863), .Y (n_1232));
INVX2 g17674(.A (n_981), .Y (n_1056));
INVX1 g17662(.A (n_965), .Y (n_980));
INVX1 g17168(.A (n_1141), .Y (n_1195));
CLKBUFX1 g17658(.A (n_1366), .Y (n_1435));
INVX1 g17160(.A (n_7656), .Y (n_1125));
INVX2 g17606(.A (n_1181), .Y (n_1070));
CLKBUFX3 g17362(.A (n_1158), .Y (n_2046));
INVX1 g17713(.A (n_979), .Y (n_996));
INVX2 g17692(.A (n_939), .Y (n_1578));
NAND2X1 g17370(.A (n_912), .B (n_852), .Y (n_1099));
AOI22X1 g18062(.A0 (n_716), .A1 (n_835), .B0 (n_941), .B1 (FP_R_14),.Y (n_977));
NAND2X1 g18090(.A (n_731), .B (n_775), .Y (n_973));
INVX2 g17619(.A (n_972), .Y (n_1213));
INVX1 g17343(.A (n_7441), .Y (n_971));
INVX1 g17612(.A (n_7686), .Y (n_1065));
INVX2 g17310(.A (n_891), .Y (n_1102));
CLKBUFX3 g17340(.A (n_7701), .Y (n_1358));
NAND2X1 g17070(.A (n_7632), .B (n_1495), .Y (n_970));
INVX2 g17654(.A (n_967), .Y (n_1229));
INVX1 g17450(.A (n_966), .Y (n_1089));
CLKBUFX3 g17425(.A (n_7705), .Y (n_1340));
INVX2 g17437(.A (n_1050), .Y (n_992));
INVX2 g17661(.A (n_965), .Y (n_1656));
INVX1 g17501(.A (n_964), .Y (n_1031));
INVX1 g17560(.A (n_1543), .Y (n_1076));
INVX1 g17570(.A (n_1538), .Y (n_1075));
INVX2 g17221(.A (n_955), .Y (n_963));
INVX2 g17287(.A (n_789), .Y (n_1115));
NAND2X1 g16743(.A (n_958), .B (n_864), .Y (n_962));
CLKBUFX1 g17236(.A (n_1495), .Y (n_2541));
INVX1 g17294(.A (n_1144), .Y (n_1104));
NAND2X1 g16901(.A (n_1180), .B (n_1682), .Y (n_1419));
CLKBUFX3 g17163(.A (n_1200), .Y (n_1677));
CLKBUFX1 g17173(.A (n_1517), .Y (n_1499));
NAND2X2 g16710(.A (n_958), .B (n_883), .Y (n_1424));
INVX2 g17207(.A (n_957), .Y (n_1598));
INVX2 g17211(.A (n_957), .Y (n_2131));
INVX1 g17220(.A (n_955), .Y (n_956));
INVX4 g17227(.A (n_955), .Y (n_2029));
CLKBUFX1 g17230(.A (n_1696), .Y (n_2146));
INVX1 g17232(.A (n_954), .Y (n_2203));
NAND2X1 g16754(.A (n_1154), .B (n_2020), .Y (n_1415));
CLKBUFX3 g17264(.A (n_1339), .Y (n_2086));
INVX2 g17273(.A (n_953), .Y (n_1107));
INVX2 g17301(.A (n_6838), .Y (n_1103));
INVX2 g17315(.A (n_1173), .Y (n_1100));
INVX2 g17342(.A (n_7441), .Y (n_1329));
INVX2 g17350(.A (n_950), .Y (n_951));
INVX1 g17371(.A (n_948), .Y (n_1918));
CLKBUFX3 g17377(.A (n_7635), .Y (n_1770));
CLKBUFX3 g17386(.A (n_1184), .Y (n_1733));
INVX1 g17278(.A (n_947), .Y (n_1093));
INVX2 g17465(.A (n_1168), .Y (n_1088));
INVX2 g17471(.A (n_1152), .Y (n_1005));
INVX1 g17505(.A (n_1682), .Y (n_1082));
INVX1 g17539(.A (n_943), .Y (n_2505));
AOI21X1 g18067(.A0 (n_941), .A1 (FP_R_18), .B0 (n_760), .Y (n_942));
INVX2 g17585(.A (n_1258), .Y (n_1204));
INVX1 g17597(.A (n_1418), .Y (n_1071));
INVX1 g17635(.A (n_905), .Y (n_1063));
INVX1 g17641(.A (n_1381), .Y (n_1061));
INVX1 g17645(.A (n_1703), .Y (n_1225));
INVX2 g17687(.A (n_1041), .Y (n_1054));
CLKBUFX3 g17700(.A (n_1666), .Y (n_2199));
INVX1 g17767(.A (n_1572), .Y (n_1047));
CLKBUFX1 g17790(.A (n_1603), .Y (n_1987));
INVX1 g17797(.A (n_1193), .Y (n_1028));
INVX1 g17803(.A (n_1134), .Y (n_1033));
INVX1 g17547(.A (n_937), .Y (n_1106));
CLKBUFX3 g17260(.A (n_1622), .Y (n_2039));
INVX2 g17520(.A (n_1149), .Y (n_1081));
OR2X1 g17983(.A (n_754), .B (n_759), .Y (n_935));
INVX2 g17680(.A (n_1171), .Y (n_1221));
AOI22X1 g18057(.A0 (n_722), .A1 (n_835), .B0 (n_941), .B1 (FP_R_22),.Y (n_934));
INVX2 g17244(.A (n_829), .Y (n_1013));
INVX1 g17250(.A (n_1388), .Y (n_1113));
INVX1 g17255(.A (n_1279), .Y (n_1109));
AND2X1 g17962(.A (n_761), .B (n_559), .Y (n_931));
MX2X1 g18054(.A (n_726), .B (FP_R_4), .S0 (n_610), .Y (n_929));
OAI21X1 g18084(.A0 (n_724), .A1 (n_733), .B0 (n_719), .Y (n_928));
OAI21X1 g18086(.A0 (n_732), .A1 (n_614), .B0 (n_702), .Y (n_927));
CLKBUFX3 g17788(.A (n_926), .Y (n_1372));
NAND2X1 g18092(.A (R_95), .B (n_764), .Y (n_925));
NAND2X1 g18231(.A (n_2298), .B (desIn[9]), .Y (n_924));
NAND3X1 g18127(.A (n_733), .B (FP_R_9), .C (n_7824), .Y (n_923));
INVX2 g17491(.A (n_922), .Y (n_1085));
INVX2 g17354(.A (n_950), .Y (n_1634));
INVX2 g17781(.A (n_1215), .Y (n_1043));
INVX2 g17218(.A (n_1397), .Y (n_1116));
INVX2 g17772(.A (n_1182), .Y (n_1046));
INVX1 g17482(.A (n_1611), .Y (n_1015));
NAND2X1 g16870(.A (n_1337), .B (n_1625), .Y (n_920));
CLKBUFX3 g17477(.A (n_1170), .Y (n_1767));
CLKBUFX3 g17474(.A (n_1687), .Y (n_1943));
NAND2X1 g18224(.A (n_2298), .B (desIn[23]), .Y (n_919));
INVX2 g17760(.A (n_918), .Y (n_1007));
INVX4 g17734(.A (n_938), .Y (n_1343));
INVX4 g17458(.A (n_915), .Y (n_1711));
INVX1 g17324(.A (n_1160), .Y (n_1206));
INVX2 g17443(.A (n_7637), .Y (n_995));
INVX1 g17720(.A (n_854), .Y (n_993));
INVX2 g17415(.A (n_999), .Y (n_1094));
INVX1 g17703(.A (n_1666), .Y (n_990));
INVX1 g17196(.A (n_1627), .Y (n_1541));
CLKBUFX1 g17708(.A (n_1485), .Y (n_1330));
INVX1 g17422(.A (n_1188), .Y (n_983));
NAND2X1 g17699(.A (n_912), .B (n_6874), .Y (n_988));
INVX2 g17187(.A (n_7354), .Y (n_997));
NAND2X2 g17688(.A (n_888), .B (n_881), .Y (n_1041));
NAND2X2 g17809(.A (n_869), .B (n_448), .Y (n_1380));
NAND2X2 g17789(.A (n_6758), .B (n_828), .Y (n_926));
NAND3X1 g17982(.A (n_729), .B (n_680), .C (n_700), .Y (n_909));
NAND2X2 g17174(.A (n_7662), .B (n_784), .Y (n_1517));
NAND2X2 g17791(.A (n_7805), .B (n_902), .Y (n_1603));
NAND3X1 g18133(.A (n_714), .B (R_96), .C (n_7859), .Y (n_908));
CLKBUFX3 g17664(.A (n_1156), .Y (n_1600));
NAND2X2 g17773(.A (n_865), .B (n_884), .Y (n_1182));
NAND2X2 g17164(.A (n_881), .B (n_877), .Y (n_1200));
NAND2X2 g17385(.A (n_849), .B (n_7806), .Y (n_6053));
NAND2X2 g17646(.A (n_840), .B (n_7349), .Y (n_1703));
NAND2X2 g17155(.A (n_886), .B (n_860), .Y (n_5927));
NAND2X2 g17642(.A (n_858), .B (n_901), .Y (n_1381));
NAND2X1 g17636(.A (n_876), .B (n_815), .Y (n_905));
NAND2X1 g17655(.A (n_885), .B (n_870), .Y (n_967));
NAND2X2 g17607(.A (n_872), .B (n_881), .Y (n_1181));
NAND2X2 g17620(.A (n_6560), .B (n_6837), .Y (n_972));
NAND2X2 g17593(.A (n_7805), .B (n_6962), .Y (n_921));
NAND2X2 g17338(.A (n_814), .B (n_7349), .Y (n_1325));
NAND2X2 g17316(.A (n_6794), .B (n_786), .Y (n_1173));
NAND2X2 g17675(.A (n_902), .B (n_901), .Y (n_981));
NAND2X2 g17598(.A (n_873), .B (n_855), .Y (n_1418));
NAND2X2 g17521(.A (n_766), .B (n_899), .Y (n_1149));
NAND2X1 g18226(.A (n_3677), .B (desIn[45]), .Y (n_898));
NAND2X2 g17475(.A (n_793), .B (n_815), .Y (n_1687));
CLKBUFX3 g17586(.A (n_1180), .Y (n_1258));
NAND2X1 g17311(.A (n_861), .B (n_6564), .Y (n_891));
NAND2X2 g17727(.A (n_6831), .B (n_881), .Y (n_914));
INVX1 g17373(.A (n_2074), .Y (n_948));
INVX2 g17212(.A (n_1346), .Y (n_957));
INVX2 g17331(.A (n_889), .Y (n_968));
NAND2X2 g17274(.A (n_798), .B (n_790), .Y (n_953));
NAND2X2 g17251(.A (n_871), .B (n_886), .Y (n_1388));
NAND2X2 g17265(.A (n_884), .B (n_885), .Y (n_1339));
NAND2X2 g17231(.A (n_785), .B (n_883), .Y (n_1696));
NAND2X2 g17193(.A (n_788), .B (n_866), .Y (n_1349));
NAND2X2 g17180(.A (n_868), .B (n_881), .Y (n_5912));
NAND2X1 g18253(.A (n_879), .B (FP_R_25), .Y (n_880));
NAND2X1 g18245(.A (n_755), .B (desIn[55]), .Y (n_878));
NAND2X2 g17169(.A (n_867), .B (n_870), .Y (n_1141));
NAND2X1 g17548(.A (n_876), .B (n_6795), .Y (n_937));
CLKBUFX3 g17197(.A (n_2020), .Y (n_1627));
CLKBUFX1 g17205(.A (n_1625), .Y (n_1753));
MX2X1 g18206(.A (R_99), .B (FP_R_5), .S0 (n_7824), .Y (n_874));
NAND2X2 g17295(.A (n_783), .B (n_873), .Y (n_1144));
NAND2X2 g17319(.A (n_871), .B (n_872), .Y (n_6070));
NAND2X2 g17325(.A (n_843), .B (n_870), .Y (n_1160));
INVX2 g17355(.A (n_1154), .Y (n_950));
NAND2X2 g17363(.A (n_868), .B (n_901), .Y (n_1158));
NAND2X2 g17391(.A (n_853), .B (n_548), .Y (n_1184));
NAND2X2 g17279(.A (n_866), .B (n_867), .Y (n_947));
NAND2X2 g17403(.A (n_856), .B (n_883), .Y (n_863));
NAND2X2 g17409(.A (n_6753), .B (n_777), .Y (n_1162));
NAND2X1 g17451(.A (n_861), .B (n_860), .Y (n_966));
NAND2X2 g17483(.A (n_839), .B (n_870), .Y (n_1611));
NAND2X1 g17531(.A (n_815), .B (n_7353), .Y (n_859));
NAND2X2 g17537(.A (n_791), .B (n_852), .Y (n_1374));
INVX1 g17541(.A (n_1355), .Y (n_943));
NAND2X2 g17555(.A (n_858), .B (n_7805), .Y (n_7733));
NAND2X2 g17561(.A (n_846), .B (n_6795), .Y (n_1543));
NAND2X2 g17571(.A (n_7335), .B (n_887), .Y (n_1538));
NAND2X2 g17659(.A (n_803), .B (n_884), .Y (n_1366));
INVX1 g17663(.A (n_1156), .Y (n_965));
NAND2X2 g17709(.A (n_856), .B (n_855), .Y (n_1485));
NAND2X1 g17721(.A (n_853), .B (n_852), .Y (n_854));
INVX2 g17737(.A (n_7633), .Y (n_938));
NAND2X2 g17756(.A (n_831), .B (n_887), .Y (n_1052));
NAND2X2 g17761(.A (n_849), .B (n_6648), .Y (n_918));
MX2X1 g18060(.A (n_684), .B (FP_R), .S0 (n_610), .Y (n_848));
NAND2X2 g17261(.A (n_846), .B (n_842), .Y (n_1622));
NAND2X2 g17681(.A (n_792), .B (n_7806), .Y (n_1171));
NAND2X2 g17804(.A (n_843), .B (n_842), .Y (n_1134));
NAND2X2 g17256(.A (n_866), .B (n_840), .Y (n_1279));
INVX1 g17512(.A (n_1724), .Y (n_932));
NAND2X2 g17798(.A (n_839), .B (n_884), .Y (n_1193));
OAI22X1 g18061(.A0 (n_696), .A1 (n_836), .B0 (n_835), .B1 (n_695), .Y(n_838));
OAI22X1 g18064(.A0 (n_711), .A1 (n_836), .B0 (n_835), .B1 (n_710), .Y(n_837));
OAI22X1 g18065(.A0 (n_693), .A1 (n_836), .B0 (n_835), .B1 (n_692), .Y(n_834));
OAI22X1 g18070(.A0 (n_698), .A1 (n_836), .B0 (n_835), .B1 (n_697), .Y(n_833));
NAND2X2 g17502(.A (n_831), .B (n_790), .Y (n_964));
NAND2X2 g17245(.A (n_828), .B (n_883), .Y (n_829));
OAI22X1 g18088(.A0 (n_66), .A1 (n_730), .B0 (n_764), .B1 (n_41), .Y(n_827));
NAND2X1 g18094(.A (FP_R_1), .B (n_730), .Y (n_826));
NAND3X1 g18106(.A (n_714), .B (FP_R_17), .C (n_7813), .Y (n_825));
NAND3X1 g18116(.A (n_714), .B (FP_R_2), .C (n_7813), .Y (n_822));
NAND3X1 g18124(.A (n_714), .B (R_111), .C (n_7812), .Y (n_821));
MX2X1 g18144(.A (R_119), .B (FP_R_25), .S0 (n_7813), .Y (n_820));
MX2X1 g18145(.A (R_124), .B (FP_R_30), .S0 (n_7858), .Y (n_818));
NAND2X1 g18229(.A (n_3677), .B (desIn[61]), .Y (n_817));
NAND2X2 g17492(.A (n_7661), .B (n_815), .Y (n_922));
NAND2X2 g17782(.A (n_814), .B (n_6837), .Y (n_1215));
MX2X1 g18202(.A (R_115), .B (FP_R_21), .S0 (n_7813), .Y (n_812));
MX2X1 g18213(.A (R_123), .B (FP_R_29), .S0 (n_7824), .Y (n_811));
NAND2X1 g18216(.A (n_610), .B (FP_R_9), .Y (n_810));
NAND2X1 g18225(.A (n_755), .B (desIn[13]), .Y (n_809));
NAND2X1 g18248(.A (n_755), .B (desIn[11]), .Y (n_808));
NAND2X2 g17768(.A (n_7335), .B (n_766), .Y (n_1572));
NAND2X2 g17478(.A (n_803), .B (n_6758), .Y (n_1170));
INVX1 g17234(.A (n_1667), .Y (n_954));
CLKBUFX1 g17762(.A (n_1681), .Y (n_2368));
OAI21X1 g18063(.A0 (n_709), .A1 (n_836), .B0 (n_690), .Y (n_801));
NAND2X2 g17472(.A (n_797), .B (n_6648), .Y (n_1152));
NAND2X2 g17219(.A (n_781), .B (n_870), .Y (n_1397));
NAND2X2 g17751(.A (n_798), .B (n_852), .Y (n_1550));
INVX2 g17228(.A (n_773), .Y (n_955));
NAND2X2 g17466(.A (n_797), .B (n_790), .Y (n_1168));
AND2X1 g18100(.A (FP_R_10), .B (n_730), .Y (n_796));
INVX2 g17460(.A (n_794), .Y (n_915));
INVX1 g18392(.A (n_3550), .Y (n_1268));
INVX8 g18530(.A (n_1776), .Y (n_3677));
NAND2X2 g17438(.A (n_792), .B (n_6837), .Y (n_1050));
NAND2X2 g17714(.A (n_791), .B (n_790), .Y (n_979));
NAND2X2 g17288(.A (n_788), .B (n_766), .Y (n_789));
NAND2X2 g17432(.A (n_786), .B (n_881), .Y (n_1163));
NAND2X2 g17704(.A (n_779), .B (n_783), .Y (n_1666));
NAND2X2 g17416(.A (n_6790), .B (n_871), .Y (n_999));
NAND2X2 g17423(.A (n_781), .B (n_6837), .Y (n_1188));
INVX2 g17695(.A (n_1337), .Y (n_939));
NAND4X1 g17170(.A (n_497), .B (n_321), .C (n_553), .D (n_239), .Y(n_958));
NAND2X2 g17542(.A (n_746), .B (n_6837), .Y (n_1355));
NAND2X2 g17332(.A (n_778), .B (n_7806), .Y (n_889));
NAND2X2 g17374(.A (n_778), .B (n_777), .Y (n_2074));
NAND2X2 g17627(.A (n_770), .B (n_815), .Y (n_5836));
NAND2X2 g17507(.A (n_768), .B (n_777), .Y (n_1682));
NAND2X1 g18093(.A (R_102), .B (n_764), .Y (n_775));
NAND2X2 g17665(.A (n_774), .B (n_7806), .Y (n_1156));
NAND2X2 g17213(.A (n_774), .B (n_887), .Y (n_1346));
NAND2X1 g17229(.A (n_741), .B (n_475), .Y (n_773));
NAND2X1 g18257(.A (n_1776), .B (FP_R_30), .Y (n_772));
NAND2X2 g17356(.A (n_887), .B (n_742), .Y (n_1154));
NAND2X2 g17461(.A (n_770), .B (n_7806), .Y (n_794));
NAND2X2 g17513(.A (n_768), .B (n_855), .Y (n_1724));
NAND2X2 g17587(.A (n_767), .B (n_766), .Y (n_1180));
AND2X1 g18091(.A (R_104), .B (n_764), .Y (n_765));
NAND2X2 g17763(.A (n_739), .B (n_7806), .Y (n_1681));
INVX8 g18531(.A (n_755), .Y (n_1776));
NAND2X1 g18056(.A (n_685), .B (n_707), .Y (n_763));
MX2X1 g18071(.A (FP_R_12), .B (n_602), .S0 (n_714), .Y (n_761));
AOI21X1 g18072(.A0 (n_544), .A1 (n_613), .B0 (n_941), .Y (n_760));
MX2X1 g18087(.A (FP_R_24), .B (n_568), .S0 (n_658), .Y (n_759));
NAND3X1 g18110(.A (n_835), .B (R_103), .C (n_7812), .Y (n_758));
NAND2X1 g18234(.A (n_755), .B (desIn[35]), .Y (n_756));
INVX1 g18140(.A (n_715), .Y (n_754));
MX2X1 g18143(.A (R_114), .B (FP_R_20), .S0 (n_7819), .Y (n_753));
NAND2X1 g18230(.A (n_755), .B (desIn[37]), .Y (n_752));
NAND4X1 g17946(.A (n_5992), .B (n_432), .C (n_5993), .D (n_233), .Y(n_912));
NAND2X1 g18228(.A (n_755), .B (desIn[15]), .Y (n_751));
NAND2X1 g18244(.A (n_701), .B (desIn[39]), .Y (n_750));
NAND2X1 g18247(.A (n_701), .B (desIn[3]), .Y (n_748));
NAND2X2 g17235(.A (n_7805), .B (n_746), .Y (n_1667));
INVX4 g18393(.A (n_714), .Y (n_3550));
NAND2X1 g18223(.A (n_701), .B (desIn[1]), .Y (n_744));
NAND2X1 g18222(.A (n_755), .B (desIn[59]), .Y (n_743));
NAND2X2 g17696(.A (n_741), .B (n_784), .Y (n_1337));
NAND2X2 g17206(.A (n_739), .B (n_842), .Y (n_1625));
INVX1 g18539(.A (n_879), .Y (n_2298));
NAND2X2 g17198(.A (n_6643), .B (n_7805), .Y (n_2020));
MX2X1 g18210(.A (R_120), .B (FP_R_26), .S0 (n_7858), .Y (n_737));
NAND2X2 g17904(.A (n_676), .B (n_626), .Y (n_843));
NAND2X2 g17905(.A (n_527), .B (n_633), .Y (n_840));
MX2X1 g18198(.A (R_107), .B (FP_R_13), .S0 (n_7819), .Y (n_736));
NAND2X2 g17920(.A (n_5612), .B (n_5613), .Y (n_872));
MX2X1 g18058(.A (n_589), .B (FP_R_23), .S0 (n_836), .Y (n_735));
NAND2X2 g17954(.A (n_611), .B (n_649), .Y (n_867));
NAND2X1 g18252(.A (n_879), .B (FP_R_20), .Y (n_732));
NAND2X2 g17933(.A (n_6096), .B (n_6097), .Y (n_865));
NAND2X2 g17919(.A (n_5627), .B (n_5628), .Y (n_853));
NAND4X1 g17906(.A (n_459), .B (n_477), .C (n_467), .D (n_260), .Y(n_828));
NAND2X2 g17909(.A (n_570), .B (n_652), .Y (n_856));
NAND2X1 g17910(.A (n_565), .B (n_659), .Y (n_868));
NAND2X2 g17915(.A (n_5677), .B (n_5678), .Y (n_849));
NAND2X2 g17922(.A (n_6043), .B (n_6044), .Y (n_793));
NAND2X2 g17929(.A (n_7585), .B (n_7586), .Y (n_785));
NAND2X2 g17930(.A (n_5658), .B (n_5659), .Y (n_877));
NAND2X2 g17935(.A (n_511), .B (n_644), .Y (n_831));
NAND2X2 g17938(.A (n_487), .B (n_657), .Y (n_797));
NAND3X1 g17943(.A (n_675), .B (n_473), .C (n_451), .Y (n_846));
NAND2X2 g17945(.A (n_532), .B (n_7511), .Y (n_858));
NAND2X2 g17949(.A (n_5690), .B (n_5691), .Y (n_902));
NAND2X2 g17952(.A (n_5966), .B (n_5967), .Y (n_888));
NAND2X2 g17953(.A (n_5662), .B (n_5663), .Y (n_786));
NAND2X1 g17956(.A (n_571), .B (n_655), .Y (n_873));
NAND2X2 g17961(.A (n_5616), .B (n_5617), .Y (n_798));
NAND2X1 g17963(.A (n_617), .B (n_612), .Y (n_779));
NAND2X1 g17959(.A (n_5707), .B (n_5708), .Y (n_861));
NAND2X2 g17958(.A (n_5647), .B (n_5648), .Y (n_792));
NAND2X1 g18119(.A (FP_R_8), .B (n_730), .Y (n_731));
NAND3X1 g18130(.A (n_658), .B (FP_R_28), .C (n_7858), .Y (n_729));
NAND2X2 g17947(.A (n_5645), .B (n_5646), .Y (n_869));
MX2X1 g18212(.A (R_100), .B (FP_R_6), .S0 (n_7858), .Y (n_728));
NAND2X1 g18215(.A (n_493), .B (n_615), .Y (n_726));
AND2X1 g18227(.A (n_755), .B (desIn[27]), .Y (n_725));
NAND2X2 g17940(.A (n_7582), .B (n_7583), .Y (n_788));
NAND2X1 g18250(.A (n_559), .B (FP_R_31), .Y (n_724));
NAND2X2 g17937(.A (n_509), .B (n_646), .Y (n_781));
NAND2X2 g17942(.A (n_5639), .B (n_5640), .Y (n_803));
NAND2X2 g17936(.A (n_5995), .B (n_5996), .Y (n_899));
NAND2X2 g17932(.A (n_7535), .B (n_7536), .Y (n_814));
MX2X1 g18205(.A (R_116), .B (FP_R_22), .S0 (n_7819), .Y (n_722));
NAND2X1 g18219(.A (n_941), .B (FP_R_2), .Y (n_721));
NAND2X1 g17925(.A (n_503), .B (n_665), .Y (n_876));
NAND2X2 g17923(.A (n_6015), .B (n_6016), .Y (n_886));
NAND2X1 g18218(.A (n_941), .B (FP_R_17), .Y (n_720));
NAND2X1 g17907(.A (n_507), .B (n_622), .Y (n_885));
NAND2X2 g17921(.A (n_7757), .B (n_7758), .Y (n_839));
INVX2 g18540(.A (n_701), .Y (n_879));
NAND2X1 g18233(.A (n_755), .B (desIn[7]), .Y (n_719));
NAND2X2 g17917(.A (n_6085), .B (n_6086), .Y (n_791));
MX2X1 g18142(.A (R_125), .B (FP_R_31), .S0 (n_7858), .Y (n_717));
MX2X1 g18201(.A (R_108), .B (FP_R_14), .S0 (n_7824), .Y (n_716));
NAND3X1 g18141(.A (n_714), .B (n_7813), .C (FP_R_24), .Y (n_715));
MX2X1 g18207(.A (n_63), .B (n_710), .S0 (n_7858), .Y (n_711));
MX2X1 g18203(.A (n_83), .B (n_689), .S0 (n_7824), .Y (n_709));
NAND2X1 g18073(.A (n_601), .B (n_835), .Y (n_707));
INVX1 g18403(.A (n_610), .Y (n_733));
NAND2X2 g17911(.A (n_533), .B (n_586), .Y (n_746));
NAND2X2 g17957(.A (n_5631), .B (n_5632), .Y (n_774));
NAND2X1 g18242(.A (n_701), .B (desIn[29]), .Y (n_702));
NAND2X2 g17960(.A (n_6019), .B (n_6020), .Y (n_778));
NAND3X1 g18121(.A (n_835), .B (R_122), .C (n_7816), .Y (n_700));
NAND2X2 g17951(.A (n_521), .B (n_438), .Y (n_770));
NAND2X2 g17950(.A (n_5651), .B (n_5652), .Y (n_742));
MX2X1 g18204(.A (n_82), .B (n_697), .S0 (n_7819), .Y (n_698));
MX2X1 g18208(.A (n_51), .B (n_695), .S0 (n_7867), .Y (n_696));
MX2X1 g18209(.A (n_6), .B (n_692), .S0 (n_7820), .Y (n_693));
OR2X1 g18220(.A (n_835), .B (n_689), .Y (n_690));
INVX2 g18238(.A (n_730), .Y (n_764));
NOR2X1 g18256(.A (n_836), .B (n_701), .Y (n_1469));
NAND2X2 g17934(.A (n_529), .B (n_592), .Y (n_768));
NAND2X1 g18217(.A (n_836), .B (FP_R_3), .Y (n_685));
MX2X1 g18214(.A (R), .B (FP_R), .S0 (n_7858), .Y (n_684));
NAND2X1 g17916(.A (n_534), .B (n_460), .Y (n_739));
NAND2X2 g17913(.A (n_524), .B (n_452), .Y (n_741));
INVX4 g18537(.A (n_559), .Y (n_755));
NAND2X2 g17908(.A (n_7779), .B (n_7780), .Y (n_767));
OR2X1 g18221(.A (n_614), .B (n_88), .Y (n_680));
NOR2X1 g18001(.A (n_339), .B (n_469), .Y (n_5967));
AOI21X1 g18179(.A0 (n_556), .A1 (kcy1[29]), .B0 (n_447), .Y (n_676));
AOI21X1 g18014(.A0 (n_411), .A1 (kcy2[8]), .B0 (n_315), .Y (n_675));
AOI22X1 g18039(.A0 (n_619), .A1 (kcy2[28]), .B0 (n_662), .B1(kcy3[28]), .Y (n_5639));
NOR2X1 g18017(.A (n_215), .B (n_434), .Y (n_6016));
AOI22X1 g18040(.A0 (n_623), .A1 (kcy2[3]), .B0 (n_664), .B1(kcy3[3]), .Y (n_5612));
AOI21X1 g18018(.A0 (n_370), .A1 (kcy2[35]), .B0 (n_219), .Y (n_5690));
AOI22X1 g18034(.A0 (n_625), .A1 (kcy2[10]), .B0 (n_636), .B1(kcy3[10]), .Y (n_5662));
AOI22X1 g18051(.A0 (n_627), .A1 (kcy2[46]), .B0 (n_664), .B1(kcy3[46]), .Y (n_666));
AOI22X1 g18025(.A0 (n_637), .A1 (kcy2[49]), .B0 (n_664), .B1(kcy3[49]), .Y (n_665));
AOI21X1 g18019(.A0 (n_662), .A1 (kcy3[39]), .B0 (n_455), .Y (n_5645));
AOI21X1 g18007(.A0 (n_408), .A1 (kcy2[15]), .B0 (n_226), .Y (n_5707));
AOI21X1 g18006(.A0 (n_375), .A1 (kcy2[18]), .B0 (n_265), .Y (n_659));
INVX1 g18397(.A (n_610), .Y (n_658));
AOI21X1 g18010(.A0 (n_654), .A1 (kcy3[33]), .B0 (n_454), .Y (n_657));
INVX4 g18298(.A (n_6957), .Y (n_884));
AOI22X1 g18047(.A0 (n_606), .A1 (kcy2[31]), .B0 (n_654), .B1(kcy3[31]), .Y (n_655));
AOI21X1 g18002(.A0 (n_392), .A1 (kcy2[34]), .B0 (n_333), .Y (n_5627));
AOI21X1 g18003(.A0 (n_422), .A1 (kcy2[16]), .B0 (n_290), .Y (n_652));
AOI21X1 g18005(.A0 (n_386), .A1 (kcy2[2]), .B0 (n_227), .Y (n_5658));
AOI21X1 g18008(.A0 (n_421), .A1 (kcy2[41]), .B0 (n_241), .Y (n_649));
AOI21X1 g18012(.A0 (n_423), .A1 (kcy2[37]), .B0 (n_276), .Y (n_7585));
AOI21X1 g18016(.A0 (n_381), .A1 (kcy2[30]), .B0 (n_245), .Y (n_646));
AOI21X1 g18021(.A0 (n_367), .A1 (kcy2[25]), .B0 (n_337), .Y (n_5677));
AOI21X1 g18022(.A0 (n_429), .A1 (kcy2[45]), .B0 (n_295), .Y (n_644));
AOI22X1 g18023(.A0 (n_632), .A1 (kcy2[17]), .B0 (n_639), .B1(kcy3[17]), .Y (n_6085));
AOI22X1 g18026(.A0 (n_630), .A1 (kcy2[0]), .B0 (n_654), .B1(kcy3[0]), .Y (n_7535));
AOI22X1 g18028(.A0 (n_634), .A1 (kcy2[55]), .B0 (n_662), .B1(kcy3[55]), .Y (n_7582));
AOI22X1 g18030(.A0 (n_621), .A1 (kcy2[23]), .B0 (n_639), .B1(kcy3[23]), .Y (n_6096));
AOI22X1 g18033(.A0 (n_637), .A1 (kcy2[22]), .B0 (n_636), .B1(kcy3[22]), .Y (n_7757));
AOI22X1 g18036(.A0 (n_634), .A1 (kcy2[51]), .B0 (n_662), .B1(kcy3[51]), .Y (n_5647));
AOI22X1 g18037(.A0 (n_632), .A1 (kcy2[43]), .B0 (n_654), .B1(kcy3[43]), .Y (n_633));
AOI22X1 g18038(.A0 (n_630), .A1 (kcy2[50]), .B0 (n_664), .B1(kcy3[50]), .Y (n_6043));
AOI22X1 g18041(.A0 (n_627), .A1 (kcy2[42]), .B0 (n_639), .B1(kcy3[42]), .Y (n_5995));
AOI22X1 g18043(.A0 (n_625), .A1 (kcy2[29]), .B0 (n_664), .B1(kcy3[29]), .Y (n_626));
AOI22X1 g18045(.A0 (n_621), .A1 (kcy2[12]), .B0 (n_636), .B1(kcy3[12]), .Y (n_622));
AOI21X1 g18176(.A0 (n_595), .A1 (kcy1[32]), .B0 (n_445), .Y (n_618));
AOI21X1 g18182(.A0 (n_483), .A1 (kcy1[24]), .B0 (n_471), .Y (n_617));
OR2X1 g18235(.A (n_46), .B (n_7858), .Y (n_615));
NAND2X1 g18240(.A (n_614), .B (n_7857), .Y (n_730));
OR2X1 g18241(.A (n_47), .B (n_7815), .Y (n_613));
AOI21X1 g18013(.A0 (n_654), .A1 (kcy3[24]), .B0 (n_464), .Y (n_612));
AOI21X1 g18186(.A0 (n_510), .A1 (kcy1[41]), .B0 (n_443), .Y (n_611));
INVX4 g18396(.A (n_610), .Y (n_714));
INVX1 g18410(.A (n_835), .Y (n_941));
INVX4 g18308(.A (n_860), .Y (n_866));
AOI22X1 g18046(.A0 (n_606), .A1 (kcy2[54]), .B0 (n_662), .B1(kcy3[54]), .Y (n_5616));
AOI22X1 g18032(.A0 (n_538), .A1 (kcy2[14]), .B0 (n_639), .B1(kcy3[14]), .Y (n_5651));
MX2X1 g18211(.A (R_106), .B (FP_R_12), .S0 (n_7858), .Y (n_602));
MX2X1 g18200(.A (R_97), .B (FP_R_3), .S0 (n_7858), .Y (n_601));
AOI22X1 g18197(.A0 (n_595), .A1 (kcy1[28]), .B0 (kcy3[28]), .B1(n_573), .Y (n_5640));
AOI21X1 g18156(.A0 (n_518), .A1 (kcy1[46]), .B0 (n_373), .Y (n_593));
AOI22X1 g18048(.A0 (n_488), .A1 (kcy2[27]), .B0 (n_662), .B1(kcy3[27]), .Y (n_592));
INVX2 g18265(.A (n_6873), .Y (n_901));
MX2X1 g18199(.A (R_117), .B (FP_R_23), .S0 (n_7821), .Y (n_589));
AOI21X1 g18173(.A0 (n_508), .A1 (kcy1[40]), .B0 (n_427), .Y (n_6015));
AOI22X1 g18169(.A0 (n_549), .A1 (kcy1[35]), .B0 (kcy3[35]), .B1(n_573), .Y (n_5691));
AOI22X1 g18027(.A0 (n_576), .A1 (kcy2[21]), .B0 (n_664), .B1(kcy3[21]), .Y (n_586));
AOI21X1 g18163(.A0 (n_528), .A1 (kcy1[20]), .B0 (n_415), .Y (n_7779));
AOI22X1 g18195(.A0 (n_485), .A1 (kcy1[42]), .B0 (kcy3[42]), .B1(n_569), .Y (n_5996));
AOI21X1 g18152(.A0 (n_7133), .A1 (kcy1[17]), .B0 (n_418), .Y(n_6086));
AOI22X1 g18162(.A0 (n_522), .A1 (kcy1[25]), .B0 (kcy3[25]), .B1(n_562), .Y (n_5678));
AOI22X1 g18153(.A0 (n_574), .A1 (kcy1[14]), .B0 (kcy3[14]), .B1(n_520), .Y (n_5652));
AOI22X1 g18031(.A0 (n_576), .A1 (kcy2[11]), .B0 (n_636), .B1(kcy3[11]), .Y (n_5631));
AOI22X1 g18166(.A0 (n_574), .A1 (kcy1[0]), .B0 (kcy3[0]), .B1(n_573), .Y (n_7536));
CLKBUFX3 g18301(.A (n_6647), .Y (n_870));
INVX4 g18266(.A (n_6873), .Y (n_815));
AOI22X1 g18172(.A0 (n_542), .A1 (kcy1[31]), .B0 (n_472), .B1(kcy3[31]), .Y (n_571));
AOI22X1 g18185(.A0 (n_500), .A1 (kcy1[16]), .B0 (kcy3[16]), .B1(n_569), .Y (n_570));
AND2X1 g18246(.A (R_118), .B (n_7857), .Y (n_568));
AOI21X1 g18191(.A0 (n_525), .A1 (kcy1[34]), .B0 (n_362), .Y (n_5628));
AOI22X1 g18183(.A0 (n_563), .A1 (kcy1[18]), .B0 (kcy3[18]), .B1(n_573), .Y (n_565));
AOI22X1 g18175(.A0 (n_563), .A1 (kcy1[9]), .B0 (kcy3[9]), .B1(n_562), .Y (n_5655));
AOI21X1 g18178(.A0 (n_7133), .A1 (kcy1[50]), .B0 (n_419), .Y(n_6044));
INVX4 g18553(.A (n_559), .Y (n_701));
AOI21X1 g18190(.A0 (n_556), .A1 (kcy1[55]), .B0 (n_372), .Y (n_7583));
NAND2X1 g18076(.A (n_346), .B (kcy2[36]), .Y (n_553));
INVX4 g18290(.A (n_552), .Y (n_790));
INVX2 g18406(.A (n_614), .Y (n_610));
AOI21X1 g18177(.A0 (n_549), .A1 (kcy1[2]), .B0 (n_404), .Y (n_5659));
INVX2 g18272(.A (n_548), .Y (n_783));
OR2X1 g18258(.A (n_26), .B (n_7869), .Y (n_544));
AOI21X1 g18188(.A0 (n_542), .A1 (kcy1[54]), .B0 (n_393), .Y (n_5617));
AOI22X1 g18024(.A0 (n_538), .A1 (kcy2[32]), .B0 (n_654), .B1(kcy3[32]), .Y (n_539));
AOI22X1 g18050(.A0 (n_536), .A1 (kcy2[53]), .B0 (n_636), .B1(kcy3[53]), .Y (n_6020));
NAND2X1 g18080(.A (n_351), .B (kcy2[47]), .Y (n_5992));
AOI22X1 g18148(.A0 (n_431), .A1 (kcy1[44]), .B0 (kcy3[44]), .B1(n_569), .Y (n_534));
AOI21X1 g18149(.A0 (n_530), .A1 (kcy1[21]), .B0 (n_430), .Y (n_533));
AOI22X1 g18150(.A0 (n_515), .A1 (kcy1[4]), .B0 (kcy3[4]), .B1(n_573), .Y (n_532));
AOI21X1 g18151(.A0 (n_530), .A1 (kcy1[11]), .B0 (n_405), .Y (n_5632));
AOI21X1 g18154(.A0 (n_528), .A1 (kcy1[27]), .B0 (n_355), .Y (n_529));
AOI21X1 g18155(.A0 (n_7133), .A1 (kcy1[43]), .B0 (n_360), .Y (n_527));
AOI22X1 g18158(.A0 (n_506), .A1 (kcy1[38]), .B0 (kcy3[38]), .B1(n_282), .Y (n_524));
AOI21X1 g18160(.A0 (n_522), .A1 (kcy1[39]), .B0 (n_359), .Y (n_5646));
AOI22X1 g18161(.A0 (n_512), .A1 (kcy1[19]), .B0 (kcy3[19]), .B1(n_520), .Y (n_521));
AOI21X1 g18164(.A0 (n_518), .A1 (kcy1[23]), .B0 (n_387), .Y (n_6097));
AOI22X1 g18165(.A0 (n_502), .A1 (kcy1[22]), .B0 (kcy3[22]), .B1(n_562), .Y (n_7758));
AOI22X1 g18168(.A0 (n_515), .A1 (kcy1[15]), .B0 (kcy3[15]), .B1(n_569), .Y (n_5708));
AOI22X1 g18170(.A0 (n_504), .A1 (kcy1[53]), .B0 (kcy3[53]), .B1(n_520), .Y (n_6019));
AOI21X1 g18171(.A0 (n_512), .A1 (kcy1[51]), .B0 (n_391), .Y (n_5648));
AOI21X1 g18174(.A0 (n_510), .A1 (kcy1[45]), .B0 (n_402), .Y (n_511));
AOI22X1 g18180(.A0 (n_508), .A1 (kcy1[30]), .B0 (n_5676), .B1(kcy3[30]), .Y (n_509));
AOI22X1 g18184(.A0 (n_506), .A1 (kcy1[12]), .B0 (kcy3[12]), .B1(n_573), .Y (n_507));
AOI21X1 g18192(.A0 (n_502), .A1 (kcy1[49]), .B0 (n_400), .Y (n_503));
AOI21X1 g18193(.A0 (n_500), .A1 (kcy1[52]), .B0 (n_388), .Y (n_5966));
AOI22X1 g18194(.A0 (n_498), .A1 (kcy1[3]), .B0 (kcy3[3]), .B1(n_356), .Y (n_5613));
NOR2X1 g18259(.A (n_358), .B (n_269), .Y (n_497));
INVX1 g18286(.A (n_852), .Y (n_855));
INVX4 g18309(.A (n_6757), .Y (n_860));
INVX4 g18313(.A (n_7348), .Y (n_881));
OR2X1 g18249(.A (n_5), .B (n_7869), .Y (n_493));
CLKBUFX1 g18408(.A (n_494), .Y (n_836));
INVX2 g18411(.A (n_494), .Y (n_835));
AOI21X1 g18196(.A0 (n_490), .A1 (kcy1[10]), .B0 (n_349), .Y (n_5663));
AOI22X1 g18042(.A0 (n_488), .A1 (kcy2[20]), .B0 (n_639), .B1(kcy3[20]), .Y (n_7780));
AOI21X1 g18167(.A0 (n_450), .A1 (kcy1[33]), .B0 (n_406), .Y (n_487));
AOI21X1 g18146(.A0 (n_483), .A1 (kcy1[37]), .B0 (n_380), .Y (n_7586));
INVX2 g18267(.A (n_6874), .Y (n_842));
INVX1 g18646(.A (n_3121), .Y (n_2813));
NAND2X1 g18251(.A (n_476), .B (kcy1[48]), .Y (n_477));
INVX2 g18274(.A (n_475), .Y (n_784));
INVX2 g18285(.A (n_449), .Y (n_852));
NAND2X1 g18429(.A (kcy3[8]), .B (n_472), .Y (n_473));
NOR2X1 g18556(.A (n_92), .B (n_446), .Y (n_471));
AOI21X1 g18078(.A0 (n_7508), .A1 (n_7505), .B0 (n_73), .Y (n_469));
INVX4 g18271(.A (n_475), .Y (n_766));
INVX2 g18289(.A (n_466), .Y (n_883));
NAND2X1 g18081(.A (n_283), .B (kcy2[48]), .Y (n_467));
INVX2 g18292(.A (n_466), .Y (n_552));
INVX2 g18275(.A (n_475), .Y (n_864));
AOI21X1 g18079(.A0 (n_463), .A1 (n_420), .B0 (n_65), .Y (n_464));
CLKBUFX1 g18415(.A (n_439), .Y (n_494));
CLKBUFX3 g18278(.A (n_475), .Y (n_871));
AOI21X1 g18011(.A0 (n_181), .A1 (kcy2[44]), .B0 (n_320), .Y (n_460));
NAND2X1 g18565(.A (kcy3[48]), .B (n_472), .Y (n_459));
INVX1 g18283(.A (n_449), .Y (n_777));
AOI21X1 g18074(.A0 (n_424), .A1 (n_416), .B0 (n_64), .Y (n_455));
AOI21X1 g18082(.A0 (n_7505), .A1 (n_463), .B0 (n_86), .Y (n_454));
AOI22X1 g18049(.A0 (n_437), .A1 (kcy2[38]), .B0 (n_199), .B1(kcy3[38]), .Y (n_452));
NAND2X1 g18254(.A (n_450), .B (kcy1[8]), .Y (n_451));
INVX2 g18273(.A (n_475), .Y (n_548));
INVX1 g18276(.A (n_475), .Y (n_448));
NOR2X1 g18418(.A (n_80), .B (n_446), .Y (n_447));
NOR2X1 g18422(.A (n_27), .B (n_446), .Y (n_445));
NOR2X1 g18561(.A (n_69), .B (n_446), .Y (n_443));
INVX1 g18677(.A (n_440), .Y (n_2811));
INVX2 g18407(.A (n_439), .Y (n_614));
INVX4 g18554(.A (n_377), .Y (n_559));
AOI22X1 g18035(.A0 (n_437), .A1 (kcy2[19]), .B0 (n_636), .B1(kcy3[19]), .Y (n_438));
AOI21X1 g18075(.A0 (n_7508), .A1 (n_7037), .B0 (n_96), .Y (n_434));
NAND2X1 g18255(.A (n_431), .B (kcy1[47]), .Y (n_432));
NOR2X1 g18423(.A (n_401), .B (n_52), .Y (n_430));
NAND2X1 g18134(.A (n_425), .B (n_278), .Y (n_429));
NOR2X1 g18428(.A (n_39), .B (n_414), .Y (n_427));
NOR2X1 g18448(.A (n_10), .B (n_221), .Y (n_426));
NAND2X1 g18128(.A (n_425), .B (n_424), .Y (n_637));
NAND2X1 g18125(.A (n_369), .B (n_424), .Y (n_423));
NAND2X1 g18118(.A (n_7040), .B (n_278), .Y (n_422));
NAND2X1 g18126(.A (n_463), .B (n_420), .Y (n_421));
NOR2X1 g18568(.A (n_35), .B (n_399), .Y (n_419));
NOR2X1 g18571(.A (n_85), .B (n_397), .Y (n_418));
NAND2X1 g18138(.A (n_424), .B (n_416), .Y (n_625));
NOR2X1 g18416(.A (n_133), .B (n_376), .Y (n_439));
NOR2X1 g18560(.A (n_61), .B (n_414), .Y (n_415));
NAND2X1 g18097(.A (n_463), .B (n_7505), .Y (n_413));
NAND2X1 g18122(.A (n_7508), .B (n_7037), .Y (n_411));
NAND2X1 g18113(.A (n_424), .B (n_416), .Y (n_606));
NAND2X1 g18108(.A (n_425), .B (n_424), .Y (n_408));
NAND2X1 g18109(.A (n_7037), .B (n_7040), .Y (n_630));
NAND2X1 g18123(.A (n_7541), .B (n_365), .Y (n_621));
NAND2X1 g18101(.A (n_424), .B (n_425), .Y (n_623));
NOR2X1 g18433(.A (n_78), .B (n_217), .Y (n_406));
NOR2X1 g18424(.A (n_48), .B (n_414), .Y (n_405));
NOR2X1 g18451(.A (n_1), .B (n_243), .Y (n_404));
CLKBUFX3 g18294(.A (n_6792), .Y (n_887));
NOR2X1 g18460(.A (n_45), .B (n_401), .Y (n_402));
NOR2X1 g18453(.A (n_97), .B (n_399), .Y (n_400));
NOR2X1 g18452(.A (n_43), .B (n_397), .Y (n_398));
NOR2X1 g18431(.A (n_77), .B (n_262), .Y (n_393));
NAND2X1 g18103(.A (n_280), .B (n_7040), .Y (n_392));
NOR2X1 g18566(.A (n_8), .B (n_401), .Y (n_391));
INVX1 g18741(.A (n_390), .Y (n_3179));
NOR2X1 g18449(.A (n_42), .B (n_401), .Y (n_388));
CLKBUFX1 g18647(.A (n_2735), .Y (n_3121));
NOR2X1 g18425(.A (n_87), .B (n_397), .Y (n_387));
NAND2X1 g18105(.A (n_7508), .B (n_7505), .Y (n_386));
NAND2X1 g18129(.A (n_463), .B (n_420), .Y (n_381));
NOR2X1 g18567(.A (n_40), .B (n_397), .Y (n_380));
NOR2X1 g18455(.A (n_12), .B (n_414), .Y (n_379));
NOR2X1 g18555(.A (n_159), .B (n_376), .Y (n_377));
INVX2 g18288(.A (n_6792), .Y (n_449));
NAND2X1 g18117(.A (n_463), .B (n_420), .Y (n_375));
NOR2X1 g18557(.A (n_95), .B (n_399), .Y (n_373));
NOR2X1 g18435(.A (n_31), .B (n_262), .Y (n_372));
NAND2X1 g18115(.A (n_424), .B (n_425), .Y (n_619));
NAND2X1 g18099(.A (n_7037), .B (n_7508), .Y (n_371));
NAND2X1 g18104(.A (n_463), .B (n_7505), .Y (n_370));
NAND2X1 g18111(.A (n_364), .B (n_369), .Y (n_632));
NAND2X1 g18131(.A (n_7037), .B (n_7040), .Y (n_367));
NAND2X1 g18135(.A (n_364), .B (n_365), .Y (n_627));
NAND2X1 g18136(.A (n_424), .B (n_416), .Y (n_634));
NOR2X1 g18430(.A (n_89), .B (n_256), .Y (n_362));
NOR2X1 g18427(.A (n_37), .B (n_399), .Y (n_360));
NOR2X1 g18436(.A (n_67), .B (n_299), .Y (n_359));
NOR2X1 g18443(.A (n_62), .B (n_232), .Y (n_358));
NAND2X1 g18447(.A (kcy3[47]), .B (n_356), .Y (n_5993));
NOR2X1 g18459(.A (n_60), .B (n_217), .Y (n_355));
INVX1 g18870(.A (n_297), .Y (n_3134));
INVX1 g18293(.A (n_6792), .Y (n_466));
NAND2X1 g18098(.A (n_365), .B (n_7541), .Y (n_351));
NOR2X1 g18446(.A (n_72), .B (n_262), .Y (n_349));
BUFX3 g18279(.A (n_6562), .Y (n_475));
NAND2X1 g18107(.A (n_364), .B (n_365), .Y (n_346));
NAND2X1 g18102(.A (n_369), .B (n_338), .Y (n_576));
NAND2X1 g18426(.A (n_341), .B (n_340), .Y (n_525));
NAND2X1 g18439(.A (n_318), .B (n_302), .Y (n_508));
NAND2X1 g18420(.A (n_324), .B (n_318), .Y (n_518));
NAND2X1 g18437(.A (n_341), .B (n_340), .Y (n_510));
NOR2X1 g18347(.A (n_332), .B (n_42), .Y (n_339));
NAND2X1 g18112(.A (n_338), .B (n_369), .Y (n_536));
NOR2X1 g18362(.A (n_332), .B (n_56), .Y (n_337));
NOR2X1 g18354(.A (n_332), .B (n_89), .Y (n_333));
NAND2X1 g18563(.A (n_318), .B (n_302), .Y (n_530));
NAND2X1 g18442(.A (n_318), .B (n_324), .Y (n_515));
NAND2X1 g18434(.A (n_303), .B (n_7127), .Y (n_506));
INVX1 g18600(.A (n_183), .Y (n_3159));
NAND2X1 g18569(.A (n_324), .B (n_318), .Y (n_476));
NAND2X1 g18356(.A (n_664), .B (kcy3[36]), .Y (n_321));
NOR2X1 g18350(.A (n_332), .B (n_53), .Y (n_320));
CLKBUFX1 g18745(.A (n_2653), .Y (n_3153));
NAND2X1 g18114(.A (n_369), .B (n_338), .Y (n_538));
NAND2X1 g18450(.A (n_318), .B (n_302), .Y (n_485));
NAND2X1 g18558(.A (n_318), .B (n_302), .Y (n_490));
NOR2X1 g18364(.A (n_332), .B (n_19), .Y (n_315));
INVX1 g18798(.A (n_7437), .Y (n_2931));
NAND2X1 g18421(.A (n_303), .B (n_7127), .Y (n_522));
NAND2X1 g18432(.A (n_318), .B (n_302), .Y (n_500));
NAND2X1 g18457(.A (n_303), .B (n_302), .Y (n_563));
NAND2X1 g18454(.A (n_341), .B (n_340), .Y (n_574));
INVX2 g18773(.A (n_356), .Y (n_446));
INVX1 g18742(.A (n_2653), .Y (n_390));
NAND2X1 g18456(.A (n_303), .B (n_302), .Y (n_549));
NAND2X1 g18441(.A (n_318), .B (n_324), .Y (n_504));
INVX1 g18768(.A (n_299), .Y (n_5676));
NAND2X1 g18444(.A (n_303), .B (n_302), .Y (n_498));
INVX1 g18872(.A (n_3106), .Y (n_297));
NAND2X1 g18440(.A (n_303), .B (n_302), .Y (n_502));
NAND2X1 g18096(.A (n_338), .B (n_365), .Y (n_488));
INVX2 g18767(.A (n_299), .Y (n_472));
NAND2X1 g18438(.A (n_341), .B (n_340), .Y (n_542));
NAND2X1 g18572(.A (n_303), .B (n_302), .Y (n_450));
NOR2X1 g18348(.A (n_332), .B (n_45), .Y (n_295));
NOR2X1 g18346(.A (n_332), .B (n_54), .Y (n_290));
NAND2X1 g18445(.A (n_7130), .B (n_174), .Y (n_431));
NAND2X1 g18559(.A (n_341), .B (n_340), .Y (n_556));
NAND2X1 g18419(.A (n_303), .B (n_302), .Y (n_595));
NAND2X1 g18458(.A (n_318), .B (n_302), .Y (n_528));
NAND2X1 g18564(.A (n_318), .B (n_324), .Y (n_483));
INVX1 g18808(.A (n_191), .Y (n_2613));
NAND2X1 g18139(.A (n_338), .B (n_365), .Y (n_283));
NAND2X1 g18570(.A (n_341), .B (n_340), .Y (n_512));
INVX2 g18766(.A (n_282), .Y (n_397));
INVX1 g18611(.A (n_281), .Y (n_2490));
INVX1 g18327(.A (n_277), .Y (n_280));
INVX1 g18653(.A (n_2735), .Y (n_329));
INVX1 g18330(.A (n_277), .Y (n_278));
NAND3X1 g18575(.A (n_7579), .B (n_7580), .C (n_34), .Y (n_376));
NOR2X1 g18363(.A (n_225), .B (n_40), .Y (n_276));
INVX2 g18666(.A (n_274), .Y (n_3044));
INVX1 g18877(.A (n_207), .Y (n_2863));
INVX4 g18320(.A (n_266), .Y (n_424));
NOR2X1 g18417(.A (n_318), .B (n_50), .Y (n_269));
INVX2 g18318(.A (n_266), .Y (n_7541));
INVX1 g18630(.A (n_136), .Y (n_2635));
NOR2X1 g18365(.A (n_248), .B (n_79), .Y (n_265));
INVX1 g18681(.A (n_1719), .Y (n_440));
INVX1 g18886(.A (n_2042), .Y (n_3194));
INVX2 g18762(.A (n_569), .Y (n_262));
INVX1 g18966(.A (n_2440), .Y (n_2281));
NAND2X1 g18366(.A (n_636), .B (kcy3[48]), .Y (n_260));
INVX2 g18776(.A (n_259), .Y (n_562));
INVX4 g18936(.A (n_6801), .Y (n_2842));
INVX1 g18901(.A (n_2067), .Y (n_2744));
INVX1 g18763(.A (n_569), .Y (n_256));
INVX2 g18317(.A (n_266), .Y (n_364));
CLKBUFX1 g18873(.A (n_2134), .Y (n_3106));
INVX1 g18656(.A (n_1750), .Y (n_2436));
NOR2X1 g18358(.A (n_248), .B (n_33), .Y (n_249));
INVX2 g18752(.A (n_223), .Y (n_414));
NOR2X1 g18355(.A (n_248), .B (n_9), .Y (n_245));
INVX1 g18755(.A (n_520), .Y (n_243));
CLKBUFX1 g18746(.A (n_2666), .Y (n_2653));
NOR2X1 g18360(.A (n_248), .B (n_69), .Y (n_241));
INVX1 g18662(.A (n_240), .Y (n_2464));
NAND4X1 g18357(.A (kcy1[36]), .B (n_105), .C (n_156), .D (n_157), .Y(n_239));
INVX1 g18867(.A (n_2134), .Y (n_234));
NAND2X1 g18345(.A (n_639), .B (kcy3[47]), .Y (n_233));
INVX1 g18770(.A (n_282), .Y (n_232));
INVX2 g18769(.A (n_282), .Y (n_299));
INVX1 g18640(.A (n_1882), .Y (n_231));
INVX1 g18663(.A (n_240), .Y (n_2412));
NAND2X1 g18120(.A (n_365), .B (n_7503), .Y (n_437));
NAND3X1 g18501(.A (n_158), .B (n_149), .C (n_132), .Y (n_296));
INVX2 g18848(.A (n_7341), .Y (n_2182));
INVX4 g18772(.A (n_259), .Y (n_573));
NOR2X1 g18349(.A (n_248), .B (n_10), .Y (n_229));
NOR2X1 g18368(.A (n_248), .B (n_1), .Y (n_227));
NOR2X1 g18351(.A (n_225), .B (n_14), .Y (n_226));
INVX2 g18751(.A (n_223), .Y (n_401));
INVX1 g18754(.A (n_520), .Y (n_221));
INVX1 g18738(.A (n_2666), .Y (n_316));
NOR2X1 g18359(.A (n_248), .B (n_11), .Y (n_219));
INVX1 g18878(.A (n_207), .Y (n_2410));
INVX2 g18757(.A (n_520), .Y (n_217));
INVX2 g18759(.A (n_569), .Y (n_399));
INVX2 g18326(.A (n_277), .Y (n_420));
INVX2 g18774(.A (n_259), .Y (n_356));
NOR2X1 g18353(.A (n_225), .B (n_39), .Y (n_215));
CLKBUFX1 g18800(.A (n_7436), .Y (n_2928));
INVX2 g18707(.A (n_7126), .Y (n_340));
INVX1 g18641(.A (n_1750), .Y (n_1882));
INVX1 g18699(.A (n_1777), .Y (n_2600));
INVX1 g18664(.A (n_1719), .Y (n_240));
INVX1 g18693(.A (n_2668), .Y (n_253));
INVX1 g18675(.A (n_1719), .Y (n_274));
INVX4 g18764(.A (n_187), .Y (n_569));
INVX1 g18833(.A (n_2122), .Y (n_3054));
INVX1 g18866(.A (n_1745), .Y (n_207));
INVX1 g18902(.A (n_2719), .Y (n_2067));
INVX1 g18887(.A (n_1745), .Y (n_2042));
INVX2 g18654(.A (n_1750), .Y (n_2735));
INVX4 g18594(.A (n_199), .Y (n_332));
INVX4 g18589(.A (n_225), .Y (n_664));
INVX1 g18782(.A (n_198), .Y (n_1760));
CLKBUFX1 g18717(.A (n_2546), .Y (n_2539));
INVX4 g18321(.A (n_7503), .Y (n_266));
INVX8 g18747(.A (n_164), .Y (n_2666));
INVX1 g18949(.A (n_2402), .Y (n_192));
INVX1 g18813(.A (n_2746), .Y (n_191));
INVX1 g18612(.A (n_2680), .Y (n_281));
INVX1 g18943(.A (n_2842), .Y (n_2036));
INVX1 g18876(.A (n_1745), .Y (n_2136));
INVX2 g18758(.A (n_187), .Y (n_520));
INVX2 g18753(.A (n_187), .Y (n_223));
INVX1 g18893(.A (n_3189), .Y (n_2488));
INVX1 g18788(.A (n_2151), .Y (n_2529));
INVX1 g18604(.A (n_183), .Y (n_2432));
CLKBUFX3 g18325(.A (n_7503), .Y (n_338));
INVX1 g18684(.A (n_1777), .Y (n_2216));
INVX4 g18960(.A (n_170), .Y (n_2440));
CLKBUFX1 g18874(.A (n_1745), .Y (n_2134));
INVX2 g18331(.A (n_7503), .Y (n_277));
INVX1 g18721(.A (n_2171), .Y (n_2907));
AOI21X1 g18095(.A0 (n_105), .A1 (n_109), .B0 (n_6132), .Y (n_181));
CLKBUFX3 g18771(.A (n_180), .Y (n_282));
INVX2 g18777(.A (n_180), .Y (n_259));
INVX1 g18695(.A (n_1777), .Y (n_2637));
INVX1 g18827(.A (n_177), .Y (n_275));
INVX1 g18787(.A (n_2151), .Y (n_2548));
INVX1 g18785(.A (n_2151), .Y (n_2913));
INVX1 g18603(.A (n_183), .Y (n_2404));
INVX1 g18705(.A (n_7126), .Y (n_174));
INVX4 g18706(.A (n_7126), .Y (n_302));
INVX1 g18730(.A (n_204), .Y (n_235));
INVX1 g18928(.A (n_200), .Y (n_172));
INVX2 g18703(.A (n_7126), .Y (n_324));
INVX1 g18636(.A (n_1750), .Y (n_2692));
INVX1 g18658(.A (n_1750), .Y (n_171));
CLKBUFX1 g18814(.A (n_2746), .Y (n_2974));
INVX1 g18913(.A (n_200), .Y (n_2695));
NAND2X1 g18748(.A (n_129), .B (n_162), .Y (n_164));
INVX1 g18786(.A (n_7436), .Y (n_2151));
INVX1 g18864(.A (n_7340), .Y (n_189));
INVX4 g18581(.A (n_7131), .Y (n_303));
INVX4 g18831(.A (n_127), .Y (n_177));
AND2X1 g18683(.A (n_162), .B (n_123), .Y (n_1719));
INVX1 g18718(.A (n_1405), .Y (n_2546));
CLKBUFX3 g18585(.A (n_155), .Y (n_639));
INVX2 g18778(.A (n_6119), .Y (n_180));
INVX4 g18597(.A (n_140), .Y (n_199));
CLKBUFX1 g18694(.A (n_6600), .Y (n_2668));
CLKBUFX3 g18765(.A (n_6119), .Y (n_187));
INVX4 g18627(.A (n_136), .Y (n_2624));
OR2X1 g18574(.A (n_106), .B (n_131), .Y (n_159));
AND2X1 g18982(.A (n_157), .B (n_156), .Y (n_158));
INVX2 g18343(.A (n_145), .Y (n_365));
INVX4 g18978(.A (n_2248), .Y (n_170));
CLKBUFX3 g18587(.A (n_155), .Y (n_662));
CLKBUFX3 g18614(.A (n_2284), .Y (n_2680));
INVX1 g18335(.A (n_7507), .Y (n_425));
INVX2 g18582(.A (n_7131), .Y (n_341));
INVX1 g18905(.A (n_2144), .Y (n_1861));
CLKBUFX1 g18615(.A (n_2284), .Y (n_3049));
INVX1 g18732(.A (n_1405), .Y (n_204));
INVX2 g18338(.A (n_135), .Y (n_463));
AND2X1 g18888(.A (n_162), .B (n_149), .Y (n_1745));
INVX1 g18336(.A (n_7507), .Y (n_416));
INVX1 g18817(.A (n_127), .Y (n_2856));
INVX1 g18700(.A (n_6600), .Y (n_1777));
INVX4 g18904(.A (n_2144), .Y (n_2719));
INVX1 g18894(.A (n_2144), .Y (n_3189));
INVX1 g18715(.A (n_1405), .Y (n_2495));
INVX4 g18815(.A (n_128), .Y (n_2746));
INVX4 g18576(.A (n_7131), .Y (n_318));
INVX1 g18784(.A (n_7436), .Y (n_198));
INVX1 g18950(.A (n_6801), .Y (n_2402));
INVX2 g18593(.A (n_140), .Y (n_636));
INVX2 g18930(.A (n_7301), .Y (n_200));
INVX1 g18710(.A (n_1405), .Y (n_139));
INVX1 g18632(.A (n_136), .Y (n_1837));
INVX1 g18723(.A (n_1405), .Y (n_2171));
INVX2 g18339(.A (n_135), .Y (n_369));
INVX1 g18907(.A (n_2144), .Y (n_2752));
INVX1 g18834(.A (n_2467), .Y (n_2122));
CLKBUFX3 g18592(.A (n_140), .Y (n_248));
INVX1 g18605(.A (n_2284), .Y (n_183));
INVX1 g18837(.A (n_127), .Y (n_2686));
NAND2X1 g18635(.A (n_132), .B (n_131), .Y (n_133));
INVX2 g18590(.A (n_155), .Y (n_225));
NAND2X2 g18660(.A (n_162), .B (n_126), .Y (n_1750));
CLKBUFX3 g18586(.A (n_155), .Y (n_654));
INVX1 g18992(.A (n_157), .Y (n_7579));
AND2X1 g18616(.A (n_129), .B (n_117), .Y (n_2284));
NAND2X1 g18816(.A (n_149), .B (n_132), .Y (n_128));
INVX2 g18840(.A (n_1880), .Y (n_127));
CLKBUFX3 g18598(.A (n_6904), .Y (n_140));
INVX2 g18591(.A (n_6904), .Y (n_155));
INVX1 g18340(.A (n_7506), .Y (n_135));
NAND2X2 g18979(.A (n_124), .B (n_123), .Y (n_2248));
NAND2X2 g18734(.A (n_123), .B (n_132), .Y (n_1405));
CLKBUFX1 g18835(.A (n_1880), .Y (n_2467));
NAND2X1 g18634(.A (n_129), .B (n_124), .Y (n_136));
NAND2X2 g18909(.A (n_126), .B (n_117), .Y (n_2144));
INVX1 g18344(.A (n_7506), .Y (n_145));
INVX1 g18993(.A (n_113), .Y (n_157));
AND2X1 g18986(.A (roundSel[2]), .B (roundSel[3]), .Y (n_162));
AND2X1 g18841(.A (n_129), .B (n_132), .Y (n_1880));
INVX1 g19050(.A (n_156), .Y (n_131));
INVX1 g18994(.A (n_6495), .Y (n_113));
NOR2X1 g18985(.A (n_104), .B (roundSel[3]), .Y (n_124));
NOR2X1 g18980(.A (roundSel[0]), .B (n_34), .Y (n_123));
INVX1 g18990(.A (n_132), .Y (n_106));
INVX1 g19025(.A (n_105), .Y (n_109));
NOR2X1 g18984(.A (roundSel[1]), .B (n_7580), .Y (n_126));
AND2X1 g18981(.A (n_104), .B (roundSel[3]), .Y (n_117));
INVX1 g19051(.A (n_103), .Y (n_156));
INVX1 g19026(.A (n_102), .Y (n_105));
NOR2X1 g18991(.A (roundSel[2]), .B (roundSel[3]), .Y (n_132));
NOR2X1 g18988(.A (roundSel[0]), .B (roundSel[1]), .Y (n_149));
INVX1 g19052(.A (n_7124), .Y (n_103));
AND2X1 g18987(.A (roundSel[0]), .B (roundSel[1]), .Y (n_129));
INVX1 g19099(.A (kcy3[49]), .Y (n_97));
INVX1 g19091(.A (kcy2[40]), .Y (n_96));
INVX1 g19092(.A (kcy3[46]), .Y (n_95));
INVX1 g19046(.A (kcy2[1]), .Y (n_93));
INVX1 g19105(.A (kcy3[24]), .Y (n_92));
INVX1 g18999(.A (desIn[26]), .Y (n_91));
INVX1 g19089(.A (desIn[12]), .Y (n_90));
INVX1 g19066(.A (kcy3[34]), .Y (n_89));
INVX1 g19044(.A (FP_R_28), .Y (n_88));
INVX1 g19030(.A (kcy3[23]), .Y (n_87));
INVX1 g19019(.A (kcy2[33]), .Y (n_86));
INVX1 g19060(.A (kcy3[17]), .Y (n_85));
INVX1 g19018(.A (R_109), .Y (n_83));
INVX1 g19041(.A (R_101), .Y (n_82));
INVX1 g19047(.A (kcy3[4]), .Y (n_81));
INVX1 g19074(.A (kcy3[29]), .Y (n_80));
INVX1 g19038(.A (kcy3[18]), .Y (n_79));
INVX1 g19003(.A (kcy3[33]), .Y (n_78));
INVX1 g19111(.A (kcy3[54]), .Y (n_77));
INVX1 g19071(.A (desIn[4]), .Y (n_76));
INVX1 g19112(.A (desIn[24]), .Y (n_74));
INVX1 g19057(.A (kcy2[52]), .Y (n_73));
INVX1 g19012(.A (FP_R_46), .Y (n_99));
INVX1 g19043(.A (roundSel[2]), .Y (n_104));
INVX1 g19029(.A (kcy3[10]), .Y (n_72));
INVX1 g19095(.A (desIn[58]), .Y (n_70));
INVX1 g19013(.A (kcy3[41]), .Y (n_69));
INVX1 g19086(.A (kcy3[39]), .Y (n_67));
INVX1 g19100(.A (R_110), .Y (n_66));
INVX1 g19010(.A (FP_R_19), .Y (n_695));
INVX2 g19027(.A (decrypt), .Y (n_102));
INVX1 g19045(.A (kcy2[24]), .Y (n_65));
INVX1 g19031(.A (kcy2[39]), .Y (n_64));
INVX1 g19078(.A (R_121), .Y (n_63));
INVX1 g19056(.A (kcy3[36]), .Y (n_62));
INVX1 g19104(.A (kcy3[20]), .Y (n_61));
INVX1 g19000(.A (kcy3[27]), .Y (n_60));
INVX1 g19098(.A (kcy3[25]), .Y (n_56));
INVX1 g19039(.A (roundSel[0]), .Y (n_7580));
INVX1 g19007(.A (kcy3[16]), .Y (n_54));
INVX1 g19017(.A (kcy3[44]), .Y (n_53));
INVX1 g19032(.A (kcy3[21]), .Y (n_52));
INVX1 g19110(.A (R_113), .Y (n_51));
INVX1 g19090(.A (kcy1[36]), .Y (n_50));
INVX1 g19106(.A (desIn[40]), .Y (n_49));
INVX1 g19077(.A (FP_R_11), .Y (n_692));
INVX1 g19076(.A (kcy3[11]), .Y (n_48));
INVX1 g19065(.A (R_112), .Y (n_47));
INVX1 g19109(.A (R_98), .Y (n_46));
INVX1 g19093(.A (kcy3[45]), .Y (n_45));
INVX1 g19085(.A (kcy3[1]), .Y (n_43));
INVX1 g19082(.A (kcy3[52]), .Y (n_42));
INVX1 g19103(.A (FP_R_16), .Y (n_41));
INVX1 g19101(.A (kcy3[37]), .Y (n_40));
INVX1 g19062(.A (kcy3[40]), .Y (n_39));
INVX1 g19035(.A (FP_R_47), .Y (n_38));
INVX1 g19034(.A (kcy3[43]), .Y (n_37));
INVX1 g19004(.A (kcy3[50]), .Y (n_35));
INVX1 g19108(.A (roundSel[1]), .Y (n_34));
INVX1 g19087(.A (kcy3[5]), .Y (n_33));
INVX1 g19009(.A (kcy3[9]), .Y (n_32));
INVX1 g19058(.A (kcy3[55]), .Y (n_31));
INVX1 g19006(.A (desIn[38]), .Y (n_30));
INVX1 g19064(.A (kcy3[32]), .Y (n_27));
INVX1 g19037(.A (FP_R_27), .Y (n_710));
INVX1 g19049(.A (FP_R_18), .Y (n_26));
INVX1 g19113(.A (desIn[60]), .Y (n_25));
INVX1 g19088(.A (desIn[36]), .Y (n_24));
INVX1 g19073(.A (desIn[2]), .Y (n_23));
INVX1 g19063(.A (kcy3[8]), .Y (n_19));
INVX1 g19083(.A (desIn[52]), .Y (n_18));
INVX1 g19002(.A (desIn[50]), .Y (n_17));
INVX1 g19072(.A (desIn[42]), .Y (n_15));
INVX1 g19079(.A (kcy3[15]), .Y (n_14));
INVX1 g19070(.A (kcy3[7]), .Y (n_12));
INVX1 g19008(.A (kcy3[35]), .Y (n_11));
INVX1 g19068(.A (kcy3[6]), .Y (n_10));
INVX1 g19059(.A (kcy3[30]), .Y (n_9));
INVX1 g19080(.A (kcy3[51]), .Y (n_8));
INVX1 g19015(.A (FP_R_34), .Y (n_7));
INVX1 g19001(.A (R_105), .Y (n_6));
INVX1 g19005(.A (FP_R_4), .Y (n_5));
INVX1 g19048(.A (FP_R_15), .Y (n_689));
INVX1 g19096(.A (kcy3[2]), .Y (n_1));
INVX1 g19075(.A (desIn[14]), .Y (n_0));
INVX1 g19033(.A (FP_R_7), .Y (n_697));
INVX1 g19243(.A (n_5713), .Y (n_5711));
INVX1 g19245(.A (n_6583), .Y (n_5713));
INVX1 g19252(.A (n_5726), .Y (n_5722));
INVX4 g19260(.A (n_5726), .Y (n_5732));
INVX2 g19261(.A (n_1349), .Y (n_5726));
CLKBUFX3 g19340(.A (n_5836), .Y (n_5835));
CLKBUFX1 g19342(.A (n_5836), .Y (n_5838));
CLKBUFX3 g19384(.A (n_5912), .Y (n_5908));
CLKBUFX3 g19389(.A (n_6567), .Y (n_5921));
CLKBUFX3 g19391(.A (n_5927), .Y (n_5924));
CLKBUFX1 g19394(.A (n_5927), .Y (n_5929));
INVX4 g19395(.A (n_5935), .Y (n_5931));
CLKBUFX3 g19398(.A (n_7416), .Y (n_5935));
INVX2 g19401(.A (n_7426), .Y (n_5938));
INVX2 g19408(.A (n_7417), .Y (n_5948));
CLKBUFX1 g19424(.A (n_6673), .Y (n_5977));
CLKBUFX2 g19437(.A (n_6023), .Y (n_6022));
CLKBUFX2 g19438(.A (n_6759), .Y (n_6023));
CLKBUFX3 g19439(.A (n_6759), .Y (n_6025));
CLKBUFX1 g19440(.A (n_6759), .Y (n_6027));
INVX1 g19452(.A (n_6048), .Y (n_6047));
INVX1 g19453(.A (n_6049), .Y (n_6048));
INVX2 g19454(.A (n_3786), .Y (n_6049));
CLKBUFX3 g19455(.A (n_3786), .Y (n_6050));
CLKBUFX1 g19456(.A (n_6053), .Y (n_6052));
CLKBUFX3 g19460(.A (n_6060), .Y (n_6058));
INVX4 g19462(.A (n_6056), .Y (n_6060));
INVX2 g19463(.A (n_6053), .Y (n_6056));
CLKBUFX2 g19466(.A (n_6070), .Y (n_6065));
NAND2X2 g14(.A (n_6117), .B (n_6118), .Y (n_6119));
INVX2 g17(.A (n_7128), .Y (n_6117));
NOR2X1 g15(.A (decrypt), .B (roundSel[4]), .Y (n_6118));
MX2X1 g28(.A (n_6121), .B (n_6120), .S0 (n_7178), .Y (desOut[30]));
INVX1 g29(.A (n_6120), .Y (n_6121));
AOI22X1 g30(.A0 (desIn[30]), .A1 (n_3668), .B0 (n_2787), .B1(n_3625), .Y (n_6120));
NAND2X1 g12_dup(.A (n_6129), .B (roundSel[4]), .Y (n_6130));
INVX2 g19487(.A (roundSel[5]), .Y (n_6129));
NAND2X1 g12(.A (n_6129), .B (roundSel[4]), .Y (n_6132));
NAND2X1 g58(.A (n_5597), .B (n_5598), .Y (n_6136));
NAND2X1 g59(.A (n_4807), .B (n_4689), .Y (n_6137));
INVX1 g76(.A (n_6209), .Y (n_6151));
NAND3X1 g72(.A (n_4775), .B (n_5042), .C (n_5092), .Y (n_6153));
AND2X1 g69(.A (n_5203), .B (n_6209), .Y (n_6154));
NAND3X1 g71(.A (n_5045), .B (n_4503), .C (n_5140), .Y (n_6156));
MX2X1 g19488(.A (n_6159), .B (n_6160), .S0 (n_6165), .Y (desOut[0]));
AOI22X1 g32(.A0 (desIn[0]), .A1 (n_3631), .B0 (n_3532), .B1 (n_3625),.Y (n_6159));
INVX1 g19489(.A (n_6159), .Y (n_6160));
NOR2X1 g19490(.A (n_6164), .B (n_5447), .Y (n_6165));
NAND3X1 g19491(.A (n_6161), .B (n_6162), .C (n_6163), .Y (n_6164));
INVX1 g34(.A (n_5349), .Y (n_6161));
INVX1 g33(.A (n_5026), .Y (n_6162));
INVX1 g35(.A (n_4691), .Y (n_6163));
MX2X1 g21(.A (n_6168), .B (n_6167), .S0 (n_6169), .Y (desOut[8]));
INVX1 g22(.A (n_6167), .Y (n_6168));
AOI22X1 g23(.A0 (desIn[8]), .A1 (n_3668), .B0 (n_3534), .B1 (n_3628),.Y (n_6167));
NAND2X1 g19492(.A (n_5443), .B (n_5019), .Y (n_6169));
MX2X1 g19493(.A (n_6172), .B (n_6171), .S0 (n_6176), .Y (desOut[48]));
INVX1 g19494(.A (n_6171), .Y (n_6172));
AOI22X1 g19495(.A0 (desIn[48]), .A1 (n_3668), .B0 (n_3553), .B1(n_3625), .Y (n_6171));
OR2X1 g19496(.A (n_5400), .B (n_6175), .Y (n_6176));
NAND2X1 g19497(.A (n_5364), .B (n_6174), .Y (n_6175));
NOR2X1 g19499(.A (n_6267), .B (n_4778), .Y (n_6174));
AND2X1 g48(.A (n_6179), .B (n_2415), .Y (n_6180));
NOR2X1 g19500(.A (n_2120), .B (n_6178), .Y (n_6179));
INVX1 g54(.A (n_1806), .Y (n_6178));
AOI21X1 g19501(.A0 (n_1632), .A1 (n_2680), .B0 (n_2785), .Y (n_6181));
AOI21X1 g19502(.A0 (n_1814), .A1 (n_2412), .B0 (n_6182), .Y (n_6183));
NAND2X1 g19503(.A (n_2562), .B (n_2516), .Y (n_6182));
NOR2X1 g19504(.A (n_2121), .B (n_2786), .Y (n_6184));
MX2X1 g19505(.A (n_6187), .B (n_6186), .S0 (n_6188), .Y (desOut[6]));
INVX1 g19506(.A (n_6186), .Y (n_6187));
AOI22X1 g19507(.A0 (desIn[6]), .A1 (n_3677), .B0 (n_3548), .B1(n_3625), .Y (n_6186));
NAND3X1 g19508(.A (n_5391), .B (n_5402), .C (n_5370), .Y (n_6188));
NAND2X1 g19511(.A (n_6190), .B (n_6191), .Y (n_6192));
NAND2X1 g63(.A (n_4859), .B (n_4578), .Y (n_6190));
INVX1 g19512(.A (n_6676), .Y (n_6191));
INVX1 g19514(.A (n_7121), .Y (n_6195));
NAND2X1 g61(.A (n_6197), .B (n_6198), .Y (n_6199));
NAND2X1 g64(.A (n_4687), .B (n_7714), .Y (n_6197));
NAND2X1 g62(.A (n_5977), .B (n_4237), .Y (n_6198));
OAI21X1 g45(.A0 (n_5288), .A1 (n_5161), .B0 (n_5404), .Y (n_7906));
OAI21X1 g44(.A0 (n_6206), .A1 (n_6208), .B0 (n_6151), .Y (n_7905));
NAND2X1 g52(.A (n_5242), .B (n_5017), .Y (n_6206));
NAND2X1 g46(.A (n_5162), .B (n_6207), .Y (n_6208));
NAND2X1 g51(.A (n_7738), .B (n_7490), .Y (n_6207));
MX2X1 g50(.A (desOut[31]), .B (n_3585), .S0 (n_3752), .Y (n_6209));
NAND2X1 g19520(.A (n_5203), .B (n_5151), .Y (n_6212));
INVX1 g60(.A (desOut[25]), .Y (n_6215));
MX2X1 g19521(.A (n_929), .B (desIn[25]), .S0 (n_701), .Y(desOut[25]));
NAND4X1 g19522(.A (n_7786), .B (n_7787), .C (n_6220), .D (n_6221), .Y(n_6222));
AND2X1 g19523(.A (n_6216), .B (n_6217), .Y (n_7787));
NAND2X1 g19524(.A (n_1971), .B (n_3054), .Y (n_6216));
NAND2X1 g19525(.A (n_1556), .B (n_7301), .Y (n_6217));
NOR2X1 g19526(.A (n_3010), .B (n_3320), .Y (n_7786));
NOR2X1 g19527(.A (n_3276), .B (n_3275), .Y (n_6220));
NOR2X1 g19528(.A (n_2102), .B (n_2191), .Y (n_6221));
NAND3X1 g19529(.A (n_6226), .B (n_6227), .C (n_6228), .Y (n_6229));
NOR2X1 g19530(.A (n_6224), .B (n_6225), .Y (n_6226));
NAND3X1 g19531(.A (n_2640), .B (n_1841), .C (n_1826), .Y (n_6224));
NAND3X1 g49(.A (n_2487), .B (n_2556), .C (n_2486), .Y (n_6225));
AOI21X1 g19532(.A0 (n_1540), .A1 (n_1882), .B0 (n_3068), .Y (n_6227));
NOR2X1 g19533(.A (n_3053), .B (n_2133), .Y (n_6228));
MX2X1 g19543(.A (n_6243), .B (n_6242), .S0 (n_6244), .Y (desOut[38]));
INVX1 g19544(.A (n_6242), .Y (n_6243));
OAI21X1 g19545(.A0 (n_3530), .A1 (n_3677), .B0 (n_6241), .Y (n_6242));
OR2X1 g19546(.A (n_30), .B (n_1776), .Y (n_6241));
NAND3X1 g19547(.A (n_5425), .B (n_5417), .C (n_5158), .Y (n_6244));
AOI21X1 g19560(.A0 (n_6156), .A1 (n_6209), .B0 (n_6262), .Y (n_6263));
AND2X1 g19561(.A (n_5134), .B (n_7490), .Y (n_6262));
OAI21X1 g19562(.A0 (n_5187), .A1 (n_5067), .B0 (n_6151), .Y (n_6264));
AOI21X1 g19563(.A0 (n_6154), .A1 (n_6153), .B0 (n_6265), .Y (n_6266));
NOR3X1 g19564(.A (n_4823), .B (n_4727), .C (n_7735), .Y (n_6265));
NOR2X1 g19565(.A (n_6267), .B (n_5185), .Y (n_6268));
NOR3X1 g19566(.A (n_4134), .B (n_4055), .C (n_4384), .Y (n_6267));
NAND4X1 g19567(.A (n_6271), .B (n_6273), .C (n_6274), .D (n_6275), .Y(n_6276));
INVX1 g19568(.A (n_6270), .Y (n_6271));
AOI21X1 g19569(.A0 (n_6040), .A1 (n_5062), .B0 (n_4814), .Y (n_6270));
AOI21X1 g19570(.A0 (n_7322), .A1 (n_4866), .B0 (n_6272), .Y (n_6273));
NOR3X1 g19571(.A (n_4289), .B (n_7321), .C (n_6441), .Y (n_6272));
NAND2X1 g19572(.A (n_4635), .B (n_4634), .Y (n_6274));
NAND3X1 g19573(.A (n_4577), .B (n_6534), .C (n_4781), .Y (n_6275));
INVX1 g19575(.A (n_6277), .Y (n_6278));
OAI21X1 g19576(.A0 (n_3565), .A1 (n_3677), .B0 (n_2712), .Y (n_6277));
NAND4X1 g19577(.A (n_5698), .B (n_5440), .C (n_5699), .D (n_5293), .Y(n_6279));
NAND4X1 g19578(.A (n_6285), .B (n_6287), .C (n_6289), .D (n_6290), .Y(n_6291));
INVX1 g19579(.A (n_6284), .Y (n_6285));
NAND2X1 g19580(.A (n_6281), .B (n_6283), .Y (n_6284));
NAND2X1 g19581(.A (n_1671), .B (n_177), .Y (n_6281));
NOR2X1 g19582(.A (n_6282), .B (n_2509), .Y (n_6283));
NAND2X1 g19583(.A (n_2585), .B (n_2587), .Y (n_6282));
NOR2X1 g55(.A (n_6286), .B (n_3207), .Y (n_6287));
NAND2X1 g19584(.A (n_2700), .B (n_2658), .Y (n_6286));
NOR2X1 g19585(.A (n_2916), .B (n_6288), .Y (n_6289));
INVX1 g19586(.A (n_2699), .Y (n_6288));
AOI21X1 g56(.A0 (n_1920), .A1 (n_2811), .B0 (n_3168), .Y (n_6290));
MX2X1 g19591(.A (n_6297), .B (n_6296), .S0 (n_6299), .Y (desOut[32]));
INVX1 g19592(.A (n_6296), .Y (n_6297));
OAI21X1 g19593(.A0 (n_3485), .A1 (n_3677), .B0 (n_2715), .Y (n_6296));
NAND3X1 g19594(.A (n_6090), .B (n_6089), .C (n_6298), .Y (n_6299));
AND2X1 g19595(.A (n_5055), .B (n_5365), .Y (n_6298));
INVX1 g74(.A (n_6301), .Y (n_6302));
AOI21X1 g75(.A0 (n_1654), .A1 (n_1670), .B0 (n_7437), .Y (n_6301));
INVX1 g78(.A (n_2427), .Y (n_7594));
NAND2X1 g70(.A (n_3123), .B (n_6306), .Y (n_6307));
AOI21X1 g73(.A0 (n_1950), .A1 (n_3179), .B0 (n_2425), .Y (n_6306));
NAND2X1 g19600(.A (n_2789), .B (n_2735), .Y (n_6311));
INVX1 g77(.A (n_2909), .Y (n_7598));
NAND3X1 g19601(.A (n_6321), .B (n_6322), .C (n_6323), .Y (n_6324));
OAI21X1 g19602(.A0 (n_6316), .A1 (n_6317), .B0 (n_6320), .Y (n_6321));
NAND4X1 g19603(.A (n_7522), .B (n_5975), .C (n_6451), .D (n_5188), .Y(n_6316));
NAND2X1 g19604(.A (n_6062), .B (n_5974), .Y (n_6317));
INVX2 g19605(.A (n_7375), .Y (n_6320));
NAND2X1 g19608(.A (n_6276), .B (n_7375), .Y (n_6322));
AOI21X1 g19609(.A0 (n_5037), .A1 (n_7323), .B0 (n_5218), .Y (n_6323));
NAND4X1 g19610(.A (n_6325), .B (n_6328), .C (n_6331), .D (n_6332), .Y(n_6333));
NAND2X1 g19611(.A (n_5340), .B (n_4172), .Y (n_6325));
NAND2X1 g19612(.A (n_6326), .B (n_6327), .Y (n_6328));
NAND4X1 g19613(.A (n_4959), .B (n_5891), .C (n_5892), .D (n_4450), .Y(n_6326));
NAND2X2 g19614(.A (n_3864), .B (n_3865), .Y (n_6327));
NAND2X1 g19615(.A (n_6329), .B (n_4449), .Y (n_6331));
INVX1 g19616(.A (n_4452), .Y (n_6329));
AOI21X1 g19618(.A0 (n_4387), .A1 (n_4393), .B0 (n_5307), .Y (n_6332));
INVX1 g19620(.A (n_6334), .Y (n_6335));
AOI22X1 g19621(.A0 (desIn[16]), .A1 (n_3631), .B0 (n_3563), .B1(n_3625), .Y (n_6334));
NOR2X1 g19624(.A (n_6338), .B (n_2441), .Y (n_6339));
NAND2X1 g19625(.A (n_2444), .B (n_2226), .Y (n_6338));
NOR2X1 g19626(.A (n_6340), .B (n_3271), .Y (n_6341));
NAND2X1 g19627(.A (n_2532), .B (n_1819), .Y (n_6340));
NOR2X1 g19628(.A (n_6342), .B (n_3270), .Y (n_6343));
NAND2X1 g19629(.A (n_2443), .B (n_1818), .Y (n_6342));
NAND2X1 g19630(.A (n_2343), .B (n_3189), .Y (n_6344));
INVX1 g19635(.A (n_6802), .Y (n_6347));
NAND2X1 g19637(.A (n_6350), .B (n_6351), .Y (n_6352));
INVX1 g19638(.A (n_2070), .Y (n_6350));
NAND2X1 g19639(.A (n_1951), .B (n_2624), .Y (n_6351));
NAND2X1 g19641(.A (n_2912), .B (n_6354), .Y (n_6355));
NAND2X1 g19642(.A (n_1953), .B (n_1882), .Y (n_6354));
AOI21X1 g19644(.A0 (n_1739), .A1 (n_2856), .B0 (n_2926), .Y (n_6358));
AOI21X1 g19645(.A0 (n_1764), .A1 (n_2913), .B0 (n_6359), .Y (n_6360));
NAND2X1 g19646(.A (n_2748), .B (n_2471), .Y (n_6359));
NOR2X1 g19647(.A (n_6361), .B (n_2749), .Y (n_6362));
NAND2X1 g19648(.A (n_1884), .B (n_1740), .Y (n_6361));
NOR2X1 g19649(.A (n_2986), .B (n_2058), .Y (n_6363));
NAND3X1 g19650(.A (n_6372), .B (n_6376), .C (n_6377), .Y (n_6378));
AOI21X1 g19651(.A0 (n_5170), .A1 (n_4574), .B0 (n_6371), .Y (n_6372));
AOI21X1 g19652(.A0 (n_4867), .A1 (n_6451), .B0 (n_6320), .Y (n_6371));
AOI21X1 g19659(.A0 (n_4844), .A1 (n_7323), .B0 (n_6375), .Y (n_6376));
NOR2X1 g19660(.A (n_6373), .B (n_6374), .Y (n_6375));
NOR2X1 g19661(.A (n_4634), .B (n_4270), .Y (n_6373));
NAND2X1 g19662(.A (n_5059), .B (n_7375), .Y (n_6374));
NAND2X1 g19663(.A (n_5356), .B (n_6320), .Y (n_6377));
NAND2X1 g19664(.A (n_6382), .B (n_6384), .Y (n_6385));
MX2X1 g19665(.A (n_6379), .B (desOut[3]), .S0 (n_6381), .Y (n_6382));
AND2X1 g41(.A (n_1003), .B (n_748), .Y (n_6379));
NAND4X1 g19666(.A (n_6180), .B (n_6181), .C (n_6183), .D (n_6184), .Y(n_6381));
INVX2 g42(.A (n_6383), .Y (n_6384));
NAND2X2 g38(.A (n_3692), .B (n_3651), .Y (n_6383));
MX2X1 g19667(.A (desOut[3]), .B (n_6379), .S0 (n_6381), .Y (n_6386));
NAND2X1 g19668(.A (n_6389), .B (n_6393), .Y (n_6394));
AND2X1 g19669(.A (n_6387), .B (n_6388), .Y (n_6389));
NAND2X2 g19670(.A (n_5325), .B (n_6965), .Y (n_6387));
NAND2X1 g19671(.A (n_5267), .B (n_6966), .Y (n_6388));
NOR2X1 g19672(.A (n_6390), .B (n_5304), .Y (n_6393));
NAND2X1 g19673(.A (n_6872), .B (n_7250), .Y (n_6390));
NAND2X1 g19675(.A (n_5132), .B (n_7465), .Y (n_6391));
NAND2X1 g19676(.A (n_6387), .B (n_6388), .Y (n_6395));
NAND2X1 g19677(.A (n_6707), .B (n_6402), .Y (n_6403));
INVX2 g19679(.A (n_4539), .Y (n_6402));
CLKBUFX3 g19681(.A (n_7357), .Y (n_6400));
MX2X1 g19685(.A (n_6405), .B (n_6404), .S0 (n_6412), .Y (desOut[14]));
INVX1 g19686(.A (n_6404), .Y (n_6405));
OAI22X1 g19687(.A0 (n_1776), .A1 (n_0), .B0 (n_3522), .B1 (n_3677),.Y (n_6404));
NOR2X1 g19688(.A (n_6406), .B (n_7374), .Y (n_6412));
AOI21X1 g19689(.A0 (n_5375), .A1 (n_6062), .B0 (n_6320), .Y (n_6406));
NAND3X1 g19695(.A (n_6416), .B (n_6418), .C (n_6420), .Y (n_6421));
NOR2X1 g19696(.A (n_6415), .B (n_3181), .Y (n_6416));
NAND4X1 g19697(.A (n_2964), .B (n_2762), .C (n_2661), .D (n_6414), .Y(n_6415));
NAND2X1 g19698(.A (n_1998), .B (n_177), .Y (n_6414));
NOR2X1 g19699(.A (n_3243), .B (n_6417), .Y (n_6418));
OR2X1 g19700(.A (n_3119), .B (n_2566), .Y (n_6417));
AOI21X1 g19701(.A0 (n_2346), .A1 (n_7301), .B0 (n_6419), .Y (n_6420));
NAND2X1 g19702(.A (n_3071), .B (n_2643), .Y (n_6419));
NOR2X1 g36(.A (n_6432), .B (n_6541), .Y (n_6435));
NAND3X1 g37(.A (n_5620), .B (n_6430), .C (n_6431), .Y (n_6432));
AOI21X1 g19709(.A0 (n_1415), .A1 (n_2600), .B0 (n_2043), .Y (n_6430));
INVX1 g19710(.A (n_2152), .Y (n_6431));
NAND4X1 g19713(.A (n_6534), .B (n_6441), .C (n_6529), .D (n_6450), .Y(n_6451));
INVX4 g19714(.A (n_6989), .Y (n_6441));
NAND2X1 g19718(.A (n_3635), .B (desOut[47]), .Y (n_6436));
NAND2X1 g19719(.A (n_2293), .B (n_3634), .Y (n_6437));
INVX1 g19725(.A (n_6992), .Y (n_6450));
INVX2 g19731(.A (n_6529), .Y (n_6454));
NAND2X1 g19736(.A (n_3602), .B (desOut[39]), .Y (n_6457));
NAND2X1 g19737(.A (n_1980), .B (n_3601), .Y (n_6458));
INVX1 g19738(.A (n_6614), .Y (n_6461));
NAND3X1 g19739(.A (n_6472), .B (n_6464), .C (n_6477), .Y (n_6478));
CLKBUFX1 g19740(.A (n_6463), .Y (n_6464));
INVX1 g19741(.A (n_6583), .Y (n_6463));
INVX2 g19743(.A (n_6471), .Y (n_6472));
INVX2 g19744(.A (n_6470), .Y (n_6471));
INVX2 g19745(.A (n_6469), .Y (n_6470));
INVX2 g19746(.A (n_6468), .Y (n_6469));
MX2X1 g19747(.A (n_6466), .B (desOut[5]), .S0 (n_6467), .Y (n_6468));
INVX1 g19748(.A (desOut[5]), .Y (n_6466));
MX2X1 g19749(.A (n_735), .B (desIn[5]), .S0 (n_755), .Y (desOut[5]));
NAND4X1 g19750(.A (n_3405), .B (n_3321), .C (n_3446), .D (n_3193), .Y(n_6467));
INVX1 g19751(.A (n_6476), .Y (n_6477));
INVX2 g19752(.A (n_6475), .Y (n_6476));
INVX1 g19753(.A (n_6474), .Y (n_6475));
INVX2 g19754(.A (n_6473), .Y (n_6474));
MX2X1 g19755(.A (n_2544), .B (desOut[37]), .S0 (n_3578), .Y (n_6473));
CLKBUFX1 g1(.A (n_6469), .Y (n_6479));
INVX1 g19757(.A (n_6480), .Y (n_6481));
AOI22X1 g19758(.A0 (desIn[62]), .A1 (n_3631), .B0 (n_3529), .B1(n_3625), .Y (n_6480));
NAND2X1 g19762(.A (n_2824), .B (n_6485), .Y (n_6486));
AOI22X1 g19763(.A0 (n_3044), .A1 (n_1542), .B0 (n_2747), .B1(n_2668), .Y (n_6485));
INVX1 g19767(.A (n_2825), .Y (n_6488));
INVX1 g19768(.A (n_2398), .Y (n_6491));
INVX2 g19770(.A (n_7128), .Y (n_6495));
NAND3X1 g19777(.A (n_6500), .B (n_2911), .C (n_6501), .Y (n_6502));
NOR2X1 g19778(.A (n_2423), .B (n_2852), .Y (n_6500));
NAND2X1 g19779(.A (n_2334), .B (n_2402), .Y (n_6501));
NAND2X1 g19782(.A (n_2332), .B (n_2613), .Y (n_6504));
MX2X1 g19784(.A (desOut[33]), .B (n_7021), .S0 (n_6511), .Y (n_7615));
NOR2X1 g19788(.A (n_3379), .B (n_3501), .Y (n_6511));
NAND4X1 g19789(.A (n_7321), .B (n_6441), .C (n_6534), .D (n_6531), .Y(n_6532));
CLKBUFX1 g19801(.A (n_6985), .Y (n_6526));
INVX2 g19804(.A (n_6530), .Y (n_6531));
CLKBUFX1 g68(.A (n_6529), .Y (n_6530));
INVX2 g19805(.A (n_6528), .Y (n_6529));
NAND2X1 g70_dup(.A (n_6881), .B (n_3586), .Y (n_6528));
NAND2X1 g19806(.A (n_6882), .B (n_3586), .Y (n_6533));
INVX2 g19807(.A (n_6526), .Y (n_6534));
NAND4X1 g19808(.A (n_6536), .B (n_6537), .C (n_6538), .D (n_6540), .Y(n_6541));
NOR2X1 g19809(.A (n_6535), .B (n_2276), .Y (n_6536));
NAND2X1 g19810(.A (n_1702), .B (n_1369), .Y (n_6535));
NAND2X1 g19811(.A (n_1493), .B (n_204), .Y (n_6537));
NOR2X1 g19812(.A (n_2267), .B (n_2019), .Y (n_6538));
NOR2X1 g19813(.A (n_6539), .B (n_2030), .Y (n_6540));
NAND2X1 g19814(.A (n_1810), .B (n_1723), .Y (n_6539));
NAND2X2 g19831(.A (n_7805), .B (n_6560), .Y (n_6567));
NAND2X2 g19832(.A (n_6558), .B (n_6559), .Y (n_6560));
AOI21X1 g19833(.A0 (n_413), .A1 (kcy2[6]), .B0 (n_426), .Y (n_6558));
AOI21X1 g19834(.A0 (n_525), .A1 (kcy1[6]), .B0 (n_229), .Y (n_6559));
INVX2 g19836(.A (n_6563), .Y (n_6564));
INVX2 g19837(.A (n_6562), .Y (n_6563));
INVX2 g19838(.A (n_7345), .Y (n_6562));
NAND4X1 g19841(.A (n_6865), .B (n_6866), .C (n_6574), .D (n_6575), .Y(n_6576));
NOR2X1 g19842(.A (n_1738), .B (n_2125), .Y (n_6866));
INVX1 g19843(.A (n_6570), .Y (n_6865));
NAND3X1 g19844(.A (n_1836), .B (n_1839), .C (n_1840), .Y (n_6570));
NOR2X1 g19845(.A (n_6572), .B (n_6573), .Y (n_6574));
NAND2X1 g19846(.A (n_2126), .B (n_1747), .Y (n_6572));
INVX1 g19847(.A (n_1746), .Y (n_6573));
NOR2X1 g19848(.A (n_2280), .B (n_2757), .Y (n_6575));
INVX2 g19849(.A (n_6582), .Y (n_6583));
MX2X1 g19850(.A (n_6579), .B (n_6580), .S0 (n_6581), .Y (n_6582));
AND2X1 g19851(.A (n_6577), .B (n_6578), .Y (n_6579));
NAND2X1 g19852(.A (n_935), .B (n_559), .Y (n_6577));
NAND2X1 g19853(.A (n_701), .B (desIn[63]), .Y (n_6578));
INVX1 g19854(.A (n_6579), .Y (n_6580));
NAND4X1 g19855(.A (n_3422), .B (n_3445), .C (n_3245), .D (n_2743), .Y(n_6581));
MX2X1 g19856(.A (n_6584), .B (n_6585), .S0 (n_6594), .Y (desOut[26]));
OAI22X1 g19857(.A0 (n_1776), .A1 (n_91), .B0 (n_3515), .B1 (n_3677),.Y (n_6584));
INVX1 g19858(.A (n_6584), .Y (n_6585));
NAND2X1 g19859(.A (n_6588), .B (n_6593), .Y (n_6594));
NOR2X1 g19860(.A (n_6586), .B (n_6587), .Y (n_6588));
AOI21X1 g19861(.A0 (n_6011), .A1 (n_6012), .B0 (n_6786), .Y (n_6586));
NOR2X1 g19862(.A (n_6999), .B (n_5345), .Y (n_6587));
NOR2X1 g19863(.A (n_6589), .B (n_6592), .Y (n_6593));
NOR2X1 g19864(.A (n_4784), .B (n_4478), .Y (n_6589));
NAND2X1 g19865(.A (n_5239), .B (n_6591), .Y (n_6592));
INVX1 g19866(.A (n_6590), .Y (n_6591));
NOR2X1 g19867(.A (n_4739), .B (n_4813), .Y (n_6590));
NAND4X1 g19868(.A (n_6596), .B (n_6598), .C (n_6599), .D (n_6603), .Y(n_6604));
NOR2X1 g19869(.A (n_3255), .B (n_3383), .Y (n_6596));
NOR2X1 g19870(.A (n_6597), .B (n_2195), .Y (n_6598));
AOI21X1 g19871(.A0 (n_2542), .A1 (n_2250), .B0 (n_281), .Y (n_6597));
NOR2X1 g19872(.A (n_3013), .B (n_3014), .Y (n_6599));
AOI21X1 g19873(.A0 (n_1650), .A1 (n_2686), .B0 (n_6602), .Y (n_6603));
AOI21X1 g19874(.A0 (n_2060), .A1 (n_1616), .B0 (n_1777), .Y (n_6602));
AND2X1 g19876(.A (n_117), .B (n_149), .Y (n_6600));
NAND2X1 g19877(.A (n_6613), .B (n_6614), .Y (n_6615));
NAND2X2 g19878(.A (n_6610), .B (n_6612), .Y (n_6613));
NAND2X2 g19879(.A (n_6607), .B (n_6609), .Y (n_6610));
NAND3X1 g19880(.A (n_6611), .B (n_3414), .C (n_3487), .Y (n_6607));
NAND2X1 g19882(.A (n_3042), .B (n_2726), .Y (n_6605));
INVX1 g19883(.A (desOut[57]), .Y (n_6609));
MX2X1 g19884(.A (n_848), .B (desIn[57]), .S0 (n_701), .Y(desOut[57]));
NAND4X1 g19885(.A (n_6611), .B (n_3414), .C (n_3487), .D(desOut[57]), .Y (n_6612));
INVX1 g19886(.A (n_6605), .Y (n_6611));
NAND2X2 g19887(.A (n_6458), .B (n_6457), .Y (n_6614));
AND2X1 g19896(.A (n_639), .B (kcy3[7]), .Y (n_6621));
INVX2 g19907(.A (n_6639), .Y (n_6640));
MX2X1 g19908(.A (n_6636), .B (n_6635), .S0 (n_6638), .Y (n_6639));
INVX1 g19909(.A (n_6635), .Y (n_6636));
OAI21X1 g19910(.A0 (n_1027), .A1 (n_755), .B0 (n_924), .Y (n_6635));
NAND4X1 g19912(.A (n_3349), .B (n_3432), .C (n_3200), .D (n_3015), .Y(n_6638));
NAND2X2 g19915(.A (n_7893), .B (n_7894), .Y (n_6643));
AOI21X1 g19916(.A0 (n_490), .A1 (kcy1[7]), .B0 (n_6621), .Y (n_7894));
AOI21X1 g19917(.A0 (n_536), .A1 (kcy2[7]), .B0 (n_379), .Y (n_7893));
INVX1 g19918(.A (n_6647), .Y (n_6648));
INVX2 g19932(.A (n_6660), .Y (n_6661));
NAND2X1 g40_dup(.A (n_3748), .B (n_7022), .Y (n_6660));
NOR2X1 g20(.A (n_7227), .B (n_6675), .Y (n_6676));
NAND2X1 g21_dup(.A (n_6673), .B (n_6674), .Y (n_6675));
AND2X1 g19943(.A (n_6463), .B (n_6474), .Y (n_6673));
AND2X1 g19944(.A (n_3798), .B (n_6469), .Y (n_6674));
NAND2X1 g19945(.A (n_6673), .B (n_6674), .Y (n_6677));
NAND2X1 g19949(.A (n_3521), .B (n_1776), .Y (n_6679));
NAND2X1 g19950(.A (n_3677), .B (desIn[28]), .Y (n_6680));
NAND4X1 g19952(.A (n_7782), .B (n_7596), .C (n_7783), .D (n_6689), .Y(n_6690));
AOI21X1 g19953(.A0 (n_2350), .A1 (n_3194), .B0 (n_6684), .Y (n_7596));
NAND2X1 g53(.A (n_2638), .B (n_2479), .Y (n_6684));
AOI21X1 g19954(.A0 (n_1628), .A1 (n_2680), .B0 (n_6686), .Y (n_7783));
NAND2X1 g19955(.A (n_2929), .B (n_2477), .Y (n_6686));
NOR2X1 g19956(.A (n_3281), .B (n_3280), .Y (n_7782));
NOR2X1 g19957(.A (n_2561), .B (n_2384), .Y (n_6689));
NAND3X1 g19958(.A (n_6694), .B (n_6697), .C (n_6699), .Y (n_6700));
NOR2X1 g19959(.A (n_6693), .B (n_6307), .Y (n_6694));
NAND2X1 g19960(.A (n_6692), .B (n_6302), .Y (n_6693));
AOI21X1 g19961(.A0 (n_2373), .A1 (n_2490), .B0 (n_2420), .Y (n_6692));
INVX1 g19963(.A (n_6696), .Y (n_6697));
NAND4X1 g19964(.A (n_7597), .B (n_7598), .C (n_6311), .D (n_7594), .Y(n_6696));
INVX1 g19965(.A (n_2855), .Y (n_7597));
NOR2X1 g19966(.A (n_6698), .B (n_6502), .Y (n_6699));
NAND2X1 g57(.A (n_3138), .B (n_6504), .Y (n_6698));
NOR2X1 g19967(.A (n_7382), .B (n_6706), .Y (n_6707));
NAND2X2 g19969(.A (n_6703), .B (n_6705), .Y (n_6706));
INVX1 g19970(.A (n_7804), .Y (n_6703));
CLKBUFX3 g19972(.A (n_7376), .Y (n_6705));
MX2X1 g19991(.A (n_6727), .B (n_6726), .S0 (n_6728), .Y (desOut[40]));
INVX1 g19992(.A (n_6726), .Y (n_6727));
OAI21X1 g19993(.A0 (n_3557), .A1 (n_3677), .B0 (n_6725), .Y (n_6726));
OR2X1 g19994(.A (n_49), .B (n_1776), .Y (n_6725));
NAND3X1 g19995(.A (n_5389), .B (n_5354), .C (n_4994), .Y (n_6728));
NAND2X1 g20004(.A (n_6741), .B (n_6744), .Y (n_7600));
NAND3X1 g20005(.A (n_4668), .B (n_4479), .C (n_6740), .Y (n_6741));
NAND3X1 g20006(.A (n_4126), .B (n_6738), .C (n_7603), .Y (n_6740));
CLKBUFX1 g20007(.A (n_6940), .Y (n_6738));
CLKBUFX1 g20009(.A (n_6743), .Y (n_6744));
INVX4 g20010(.A (n_6742), .Y (n_6743));
NAND2X2 g20011(.A (n_3815), .B (n_3776), .Y (n_6742));
INVX1 g20012(.A (n_6740), .Y (n_6746));
NAND2X1 g20014(.A (n_4126), .B (n_6738), .Y (n_6748));
NAND2X2 g20015(.A (n_6753), .B (n_6758), .Y (n_6759));
NAND2X2 g20016(.A (n_6749), .B (n_6752), .Y (n_6753));
AOI21X1 g20017(.A0 (n_371), .A1 (kcy2[5]), .B0 (n_249), .Y (n_6749));
AND2X1 g20018(.A (n_6750), .B (n_6751), .Y (n_6752));
NAND2X1 g20019(.A (n_476), .B (kcy1[5]), .Y (n_6750));
NAND2X1 g20020(.A (n_562), .B (kcy3[5]), .Y (n_6751));
INVX2 g20021(.A (n_6757), .Y (n_6758));
INVX2 g20022(.A (n_7347), .Y (n_6757));
MX2X1 g20039(.A (n_6776), .B (n_6775), .S0 (n_6777), .Y (desOut[44]));
INVX1 g20040(.A (n_6775), .Y (n_6776));
AOI22X1 g20041(.A0 (desIn[44]), .A1 (n_3668), .B0 (n_3513), .B1(n_3628), .Y (n_6775));
NAND2X1 g20042(.A (n_5444), .B (n_5433), .Y (n_6777));
NAND3X1 g20043(.A (n_6779), .B (n_6782), .C (n_6788), .Y (n_6789));
NAND2X1 g20044(.A (n_5320), .B (n_5361), .Y (n_6779));
AND2X1 g20045(.A (n_6780), .B (n_6781), .Y (n_6782));
OAI21X1 g20046(.A0 (n_4819), .A1 (n_5194), .B0 (n_4955), .Y (n_6780));
NOR2X1 g20047(.A (n_4522), .B (n_6590), .Y (n_6781));
NAND2X1 g20048(.A (n_4356), .B (n_7653), .Y (n_6788));
NAND4X1 g20049(.A (n_5172), .B (n_5014), .C (n_4983), .D (n_6783), .Y(n_7653));
AND2X1 g20050(.A (n_4235), .B (n_4524), .Y (n_6783));
INVX1 g20052(.A (n_6999), .Y (n_6786));
AOI21X1 g20054(.A0 (n_6797), .A1 (n_6800), .B0 (n_6801), .Y (n_6802));
CLKBUFX1 g20055(.A (n_6796), .Y (n_6797));
NAND2X2 g20056(.A (n_6790), .B (n_6795), .Y (n_6796));
NAND2X2 g20057(.A (n_618), .B (n_539), .Y (n_6790));
INVX1 g20058(.A (n_6794), .Y (n_6795));
INVX1 g20059(.A (n_449), .Y (n_6794));
INVX2 g20061(.A (n_7345), .Y (n_6792));
INVX2 g20063(.A (n_6799), .Y (n_6800));
INVX1 g20064(.A (n_6963), .Y (n_6799));
NAND2X2 g20066(.A (n_117), .B (n_123), .Y (n_6801));
INVX1 g20069(.A (n_6801), .Y (n_6805));
CLKBUFX3 g20080(.A (n_7804), .Y (n_6816));
INVX2 g20081(.A (n_7382), .Y (n_6817));
INVX1 g20082(.A (n_7377), .Y (n_6818));
NAND3X1 g20083(.A (n_6819), .B (n_6820), .C (n_6827), .Y (n_6828));
OAI21X1 g20084(.A0 (n_4481), .A1 (n_4932), .B0 (n_4908), .Y (n_6819));
NAND2X1 g20085(.A (n_4766), .B (n_4554), .Y (n_6820));
NOR2X1 g20086(.A (n_6824), .B (n_6826), .Y (n_6827));
AND2X1 g20087(.A (n_6746), .B (n_6823), .Y (n_6824));
INVX2 g20088(.A (n_6822), .Y (n_6823));
INVX1 g20089(.A (n_6821), .Y (n_6822));
NAND2X2 g20090(.A (n_3691), .B (n_3650), .Y (n_6821));
AOI21X1 g20091(.A0 (n_4330), .A1 (n_4737), .B0 (n_6823), .Y (n_6826));
INVX1 g20093(.A (n_6824), .Y (n_6829));
INVX1 g20094(.A (n_6823), .Y (n_6830));
NAND2X1 g20095(.A (n_6831), .B (n_6837), .Y (n_6838));
NAND2X1 g20096(.A (n_593), .B (n_666), .Y (n_6831));
CLKBUFX3 g20097(.A (n_6956), .Y (n_6837));
NAND2X1 g20101(.A (n_6132), .B (n_105), .Y (n_6832));
NAND3X1 g20102(.A (n_113), .B (n_103), .C (n_102), .Y (n_6833));
INVX1 g20103(.A (n_7346), .Y (n_6647));
NAND4X1 g20104(.A (n_6842), .B (n_6843), .C (n_6845), .D (n_6847), .Y(n_6848));
AOI21X1 g20105(.A0 (n_1523), .A1 (n_3049), .B0 (n_6841), .Y (n_6842));
NAND2X1 g20106(.A (n_2678), .B (n_6840), .Y (n_6841));
INVX1 g20107(.A (n_1704), .Y (n_6840));
NOR2X1 g20108(.A (n_2652), .B (n_3009), .Y (n_6843));
AOI21X1 g20109(.A0 (n_1496), .A1 (n_2695), .B0 (n_6844), .Y (n_6845));
NAND2X1 g20110(.A (n_1852), .B (n_1863), .Y (n_6844));
NOR2X1 g20111(.A (n_6846), .B (n_2129), .Y (n_6847));
NAND2X1 g20112(.A (n_1787), .B (n_1789), .Y (n_6846));
NOR2X1 g20113(.A (n_6853), .B (n_7343), .Y (n_6857));
NAND3X1 g20114(.A (n_7589), .B (n_7590), .C (n_6852), .Y (n_6853));
INVX1 g20115(.A (n_2983), .Y (n_7590));
AOI21X1 g20116(.A0 (n_2233), .A1 (n_2974), .B0 (n_3059), .Y (n_7589));
NOR2X1 g20117(.A (n_6851), .B (n_3000), .Y (n_6852));
INVX1 g20118(.A (n_1827), .Y (n_6851));
CLKBUFX3 g20129(.A (n_6563), .Y (n_6873));
CLKBUFX1 g18269_dup(.A (n_6563), .Y (n_6874));
NAND2X1 g20130(.A (n_3758), .B (n_3736), .Y (n_6875));
NAND2X1 g15155_dup(.A (n_3758), .B (n_3736), .Y (n_6876));
MX2X1 g19931_dup(.A (n_6215), .B (desOut[25]), .S0 (n_6222), .Y(n_6878));
MX2X1 g20132(.A (n_6335), .B (n_6334), .S0 (n_7148), .Y (desOut[16]));
MX2X1 g19619_dup(.A (n_6335), .B (n_6334), .S0 (n_7148), .Y (n_6880));
NAND2X1 g20133(.A (n_7081), .B (n_3585), .Y (n_6881));
NAND2X1 g15322_dup(.A (n_7081), .B (n_3585), .Y (n_6882));
NAND2X1 g14992_dup(.A (n_7309), .B (n_7307), .Y (n_4097));
NOR2X1 g15335_dup(.A (n_7023), .B (n_7024), .Y (n_6886));
INVX1 g20137(.A (n_6890), .Y (n_6888));
INVX2 g20139(.A (n_6891), .Y (n_6890));
INVX2 g20140(.A (n_3879), .Y (n_6891));
NAND3X1 g20150(.A (n_7128), .B (n_6903), .C (decrypt), .Y (n_6904));
INVX1 g20152(.A (roundSel[4]), .Y (n_6903));
NAND3X1 g20153(.A (n_7781), .B (n_6905), .C (n_6911), .Y (n_6912));
AOI21X1 g20154(.A0 (n_4585), .A1 (n_4133), .B0 (n_5082), .Y (n_6905));
NAND2X1 g32_dup(.A (n_6906), .B (n_6909), .Y (n_7781));
NAND2X1 g20155(.A (n_5070), .B (n_5202), .Y (n_6906));
INVX1 g20156(.A (n_7122), .Y (n_6909));
NAND2X1 g34_dup(.A (n_7122), .B (n_5308), .Y (n_6911));
NAND2X1 g20159(.A (n_6909), .B (n_6906), .Y (n_6913));
NAND2X1 g20160(.A (n_7122), .B (n_5308), .Y (n_6914));
OR2X1 g20169(.A (n_6923), .B (n_7450), .Y (n_6928));
NAND4X1 g20170(.A (n_2848), .B (n_2847), .C (n_2850), .D (n_2599), .Y(n_6923));
NAND2X1 g20178(.A (n_3139), .B (n_6347), .Y (n_6930));
NAND2X1 g20179(.A (n_3125), .B (n_3126), .Y (n_6931));
NOR2X1 g20181(.A (n_7603), .B (n_7707), .Y (n_6942));
NAND2X1 g20182(.A (n_3748), .B (n_7022), .Y (n_6935));
MX2X1 g20185(.A (desOut[7]), .B (n_7305), .S0 (n_6857), .Y (n_6936));
MX2X1 g20186(.A (desOut[25]), .B (n_6215), .S0 (n_6222), .Y (n_6940));
INVX1 g20189(.A (n_6940), .Y (n_6943));
INVX2 g20190(.A (n_6936), .Y (n_6944));
NAND2X2 g20200(.A (n_884), .B (n_6962), .Y (n_6963));
INVX2 g20202(.A (n_6956), .Y (n_6957));
CLKBUFX2 g20203(.A (n_7346), .Y (n_6956));
NAND3X1 g20206(.A (n_6959), .B (n_6960), .C (n_6961), .Y (n_6962));
AOI22X1 g20207(.A0 (kcy3[13]), .A1 (n_573), .B0 (n_662), .B1(kcy3[13]), .Y (n_6959));
NAND2X1 g20208(.A (n_623), .B (kcy2[13]), .Y (n_6960));
NAND2X1 g20209(.A (n_498), .B (kcy1[13]), .Y (n_6961));
NAND4X1 g20210(.A (n_6968), .B (n_6969), .C (n_7470), .D (n_7250), .Y(n_6972));
NAND2X1 g20211(.A (n_6964), .B (n_6966), .Y (n_6968));
NAND2X1 g20212(.A (n_5280), .B (n_4796), .Y (n_6964));
INVX2 g20214(.A (n_6965), .Y (n_6966));
NAND2X2 g20215(.A (n_3814), .B (n_3775), .Y (n_6965));
NAND2X1 g20216(.A (n_6965), .B (n_7556), .Y (n_6969));
MX2X1 g20220(.A (n_6974), .B (n_6975), .S0 (n_6976), .Y (desOut[28]));
NAND2X1 g18(.A (n_6679), .B (n_6680), .Y (n_6974));
INVX1 g20221(.A (n_6974), .Y (n_6975));
NAND2X1 g16(.A (n_5430), .B (n_5407), .Y (n_6976));
NAND4X1 g20222(.A (n_6983), .B (n_6986), .C (n_6989), .D (n_6992), .Y(n_6993));
INVX1 g20223(.A (n_7320), .Y (n_6983));
AOI21X1 g67(.A0 (n_820), .A1 (n_1469), .B0 (n_1345), .Y (n_6978));
NOR2X1 g20225(.A (n_3404), .B (n_3592), .Y (n_6980));
CLKBUFX3 g20226(.A (n_6985), .Y (n_6986));
INVX4 g20227(.A (n_6984), .Y (n_6985));
MX2X1 g20228(.A (n_1980), .B (desOut[39]), .S0 (n_6291), .Y (n_6984));
INVX2 g20229(.A (n_6988), .Y (n_6989));
INVX4 g20230(.A (n_6987), .Y (n_6988));
NAND2X2 g20231(.A (n_6436), .B (n_6437), .Y (n_6987));
INVX2 g20232(.A (n_6991), .Y (n_6992));
INVX1 g20233(.A (n_6990), .Y (n_6991));
MX2X1 g20234(.A (n_6466), .B (desOut[5]), .S0 (n_7192), .Y (n_6990));
INVX1 g20235(.A (n_6992), .Y (n_6994));
XOR2X1 g20236(.A (desOut[61]), .B (n_6998), .Y (n_6999));
NAND3X1 g20239(.A (n_3568), .B (n_6997), .C (n_3423), .Y (n_6998));
AND2X1 g20240(.A (n_3341), .B (n_3342), .Y (n_6997));
NAND3X1 g20245(.A (n_7006), .B (n_6081), .C (n_3244), .Y (n_7004));
NAND2X1 g20247(.A (n_6082), .B (n_2701), .Y (n_7002));
INVX2 g20249(.A (n_7002), .Y (n_7006));
NAND2X2 g20250(.A (n_1208), .B (n_817), .Y (desOut[61]));
OAI21X1 g20259(.A0 (n_7018), .A1 (n_7020), .B0 (n_7021), .Y (n_7022));
NAND4X1 g20260(.A (n_6360), .B (n_2751), .C (n_6362), .D (n_6363), .Y(n_7018));
NAND2X1 g20261(.A (n_7019), .B (n_6358), .Y (n_7020));
AND2X1 g20262(.A (n_2628), .B (n_2473), .Y (n_7019));
AOI22X1 g20263(.A0 (n_879), .A1 (n_763), .B0 (n_755), .B1(desIn[33]), .Y (n_7021));
NAND3X1 g20264(.A (n_2751), .B (n_2628), .C (n_2473), .Y (n_7023));
NAND4X1 g20265(.A (n_6360), .B (n_6358), .C (n_6362), .D (n_6363), .Y(n_7024));
INVX1 g20269(.A (n_2474), .Y (n_7026));
NAND2X1 g20271(.A (n_2492), .B (n_2620), .Y (n_7028));
AOI21X1 g20275(.A0 (n_7041), .A1 (kcy2[9]), .B0 (n_7042), .Y(n_7043));
NAND2X1 g20276(.A (n_7037), .B (n_7040), .Y (n_7041));
INVX2 g20277(.A (n_7504), .Y (n_7037));
INVX1 g20281(.A (n_7507), .Y (n_7040));
NOR2X1 g20284(.A (n_32), .B (n_332), .Y (n_7042));
MX2X1 g20285(.A (n_7045), .B (n_7044), .S0 (n_7050), .Y (desOut[34]));
INVX1 g20286(.A (n_7044), .Y (n_7045));
AOI22X1 g20287(.A0 (n_3625), .A1 (n_3527), .B0 (n_3631), .B1(desIn[34]), .Y (n_7044));
NAND3X1 g20288(.A (n_7888), .B (n_7889), .C (n_7049), .Y (n_7050));
NAND2X1 g20289(.A (n_6828), .B (n_3899), .Y (n_7889));
NAND2X1 g20290(.A (n_5351), .B (n_5419), .Y (n_7888));
AOI21X1 g20291(.A0 (n_5129), .A1 (n_5121), .B0 (n_7048), .Y (n_7049));
AND2X1 g20292(.A (n_4909), .B (n_4561), .Y (n_7048));
MX2X1 g20302(.A (n_7062), .B (n_7061), .S0 (n_7069), .Y (desOut[46]));
INVX1 g20303(.A (n_7061), .Y (n_7062));
AOI22X1 g20304(.A0 (n_3628), .A1 (n_3531), .B0 (n_3668), .B1(desIn[46]), .Y (n_7061));
NAND3X1 g20305(.A (n_7527), .B (n_7528), .C (n_7068), .Y (n_7069));
INVX1 g20311(.A (n_5269), .Y (n_7068));
NAND2X1 g20312(.A (n_7077), .B (n_7080), .Y (n_7081));
INVX1 g20313(.A (n_7076), .Y (n_7077));
NAND4X1 g20314(.A (n_7071), .B (n_7072), .C (n_7074), .D (n_7075), .Y(n_7076));
NOR2X1 g20315(.A (n_2275), .B (n_2273), .Y (n_7071));
AND2X1 g20316(.A (n_1420), .B (n_1800), .Y (n_7072));
AOI21X1 g20317(.A0 (n_1714), .A1 (n_139), .B0 (n_7073), .Y (n_7074));
AND2X1 g20318(.A (n_6600), .B (n_1817), .Y (n_7073));
NOR2X1 g20319(.A (n_1712), .B (n_2162), .Y (n_7075));
NOR2X1 g20320(.A (n_7078), .B (n_7079), .Y (n_7080));
NAND2X1 g70_dup20321(.A (n_2845), .B (n_2394), .Y (n_7078));
NAND3X1 g20322(.A (n_7886), .B (n_7887), .C (n_2163), .Y (n_7079));
NAND2X1 g20323(.A (n_2394), .B (n_2845), .Y (n_7082));
OR2X1 g20324(.A (n_2294), .B (n_7092), .Y (n_7093));
NAND2X2 g20326(.A (n_1018), .B (n_756), .Y (desOut[35]));
NAND4X1 g20327(.A (n_7678), .B (n_7679), .C (n_7090), .D (n_7091), .Y(n_7092));
NOR2X1 g20328(.A (n_2777), .B (n_3043), .Y (n_7679));
NOR2X1 g20329(.A (n_2995), .B (n_7088), .Y (n_7678));
NAND2X1 g20330(.A (n_7086), .B (n_7087), .Y (n_7088));
INVX1 g20331(.A (n_1771), .Y (n_7086));
NAND2X1 g20332(.A (n_2763), .B (n_2624), .Y (n_7087));
NAND2X1 g20333(.A (n_1946), .B (n_2436), .Y (n_7090));
NOR2X1 g20334(.A (n_2597), .B (n_3093), .Y (n_7091));
OR2X1 g20339(.A (n_76), .B (n_3673), .Y (n_7095));
NAND2X1 g20351(.A (n_7120), .B (n_7122), .Y (n_7527));
NAND3X1 g20352(.A (n_7114), .B (n_7118), .C (n_7119), .Y (n_7120));
NOR2X1 g20353(.A (n_7112), .B (n_7113), .Y (n_7114));
NAND2X1 g20354(.A (n_7110), .B (n_7111), .Y (n_7112));
NAND4X1 g20355(.A (n_4504), .B (n_4849), .C (n_7712), .D (n_4092), .Y(n_7110));
NAND3X1 g20356(.A (n_4241), .B (n_7227), .C (n_4558), .Y (n_7111));
NAND3X1 g20357(.A (n_4952), .B (n_6677), .C (n_4678), .Y (n_7113));
NAND3X1 g20358(.A (n_4570), .B (n_4504), .C (n_7117), .Y (n_7118));
INVX1 g20361(.A (n_6464), .Y (n_7117));
OR2X1 g20362(.A (n_4677), .B (n_4454), .Y (n_7119));
CLKBUFX3 g20363(.A (n_7121), .Y (n_7122));
NAND2X1 g20364(.A (n_3893), .B (n_3894), .Y (n_7121));
NAND2X1 g20365(.A (n_7127), .B (n_303), .Y (n_7133));
INVX2 g20366(.A (n_7126), .Y (n_7127));
INVX4 g20367(.A (n_7125), .Y (n_7126));
NAND3X1 g20368(.A (n_6495), .B (n_7124), .C (decrypt), .Y (n_7125));
INVX2 g20369(.A (roundSel[4]), .Y (n_7124));
INVX4 g20371(.A (n_7130), .Y (n_7131));
NAND3X1 g20372(.A (n_7128), .B (n_7124), .C (n_7129), .Y (n_7130));
INVX2 g20373(.A (roundSel[5]), .Y (n_7128));
INVX2 g20374(.A (decrypt), .Y (n_7129));
NAND4X1 g20382(.A (n_7144), .B (n_7146), .C (n_7147), .D (n_5686), .Y(n_7148));
NAND2X1 g20383(.A (n_7141), .B (n_3899), .Y (n_7144));
NAND4X1 g20384(.A (n_5696), .B (n_5124), .C (n_5697), .D (n_4931), .Y(n_7141));
NAND2X2 g20386(.A (n_3755), .B (n_3759), .Y (n_7142));
NOR2X1 g20387(.A (n_7145), .B (n_5157), .Y (n_7146));
NAND2X1 g20388(.A (n_5687), .B (n_5212), .Y (n_7145));
NAND2X1 g20389(.A (n_5101), .B (n_4554), .Y (n_7147));
MX2X1 g20390(.A (n_7149), .B (n_7150), .S0 (n_7154), .Y (desOut[2]));
OAI22X1 g20391(.A0 (n_3561), .A1 (n_3677), .B0 (n_1776), .B1 (n_23),.Y (n_7149));
INVX1 g20392(.A (n_7149), .Y (n_7150));
NAND3X1 g20393(.A (n_7151), .B (n_7152), .C (n_7153), .Y (n_7154));
NAND2X1 g20394(.A (n_5404), .B (n_5355), .Y (n_7151));
AOI21X1 g20395(.A0 (n_5223), .A1 (n_3994), .B0 (n_5306), .Y (n_7152));
NAND2X1 g20396(.A (n_5245), .B (n_6151), .Y (n_7153));
NAND2X1 g26(.A (n_7156), .B (n_7157), .Y (n_7158));
AOI22X1 g20397(.A0 (desIn[10]), .A1 (n_3668), .B0 (n_3535), .B1(n_3628), .Y (n_7156));
NAND4X1 g20398(.A (n_5372), .B (n_5241), .C (n_5369), .D (n_4656), .Y(n_7157));
INVX1 g27(.A (n_7157), .Y (n_7159));
INVX1 g20401(.A (desOut[11]), .Y (n_7161));
OAI21X1 g20402(.A0 (n_977), .A1 (n_755), .B0 (n_808), .Y(desOut[11]));
NOR2X1 g20404(.A (n_3419), .B (n_3593), .Y (n_7163));
NAND3X1 g20405(.A (n_7166), .B (n_7176), .C (n_7177), .Y (n_7178));
NAND2X1 g20406(.A (n_5366), .B (n_5428), .Y (n_7166));
INVX1 g20407(.A (n_7175), .Y (n_7176));
NAND2X1 g20408(.A (n_7172), .B (n_7174), .Y (n_7175));
NAND2X1 g20409(.A (n_7167), .B (n_7171), .Y (n_7172));
NAND2X1 g20410(.A (n_4964), .B (n_4466), .Y (n_7167));
INVX4 g20411(.A (n_7170), .Y (n_7171));
CLKBUFX3 g20412(.A (n_7169), .Y (n_7170));
INVX2 g20413(.A (n_7168), .Y (n_7169));
MX2X1 g20414(.A (desOut[51]), .B (n_2783), .S0 (n_3683), .Y (n_7168));
NAND3X1 g20415(.A (n_5081), .B (n_4551), .C (n_7173), .Y (n_7174));
INVX1 g20416(.A (n_7171), .Y (n_7173));
OAI21X1 g20417(.A0 (n_5181), .A1 (n_5193), .B0 (n_4142), .Y (n_7177));
MX2X1 g20418(.A (n_7181), .B (n_7180), .S0 (n_7182), .Y (desOut[50]));
INVX1 g20419(.A (n_7180), .Y (n_7181));
OAI21X1 g20420(.A0 (n_3558), .A1 (n_3631), .B0 (n_7179), .Y (n_7180));
OR2X1 g20421(.A (n_17), .B (n_1776), .Y (n_7179));
NAND4X1 g20422(.A (n_6263), .B (n_6264), .C (n_6266), .D (n_6268), .Y(n_7182));
NAND4X1 g20423(.A (n_7186), .B (n_7187), .C (n_7189), .D (n_7191), .Y(n_7192));
NOR2X1 g20424(.A (n_2392), .B (n_7185), .Y (n_7186));
NAND2X1 g20425(.A (n_7184), .B (n_2694), .Y (n_7185));
INVX1 g20426(.A (n_2044), .Y (n_7184));
NOR2X1 g20427(.A (n_2656), .B (n_3019), .Y (n_7187));
AOI21X1 g20428(.A0 (n_1513), .A1 (n_2695), .B0 (n_7188), .Y (n_7189));
NAND2X1 g20429(.A (n_2258), .B (n_1865), .Y (n_7188));
AOI21X1 g20430(.A0 (n_2009), .A1 (n_204), .B0 (n_7190), .Y (n_7191));
NAND2X1 g20431(.A (n_1796), .B (n_2232), .Y (n_7190));
NAND4X1 g20432(.A (n_7194), .B (n_7195), .C (n_7197), .D (n_7198), .Y(n_7199));
INVX1 g20433(.A (n_7193), .Y (n_7194));
OAI21X1 g20434(.A0 (n_4939), .A1 (n_5948), .B0 (n_4869), .Y (n_7193));
OAI21X1 g43(.A0 (n_5300), .A1 (n_4938), .B0 (n_4172), .Y (n_7195));
INVX1 g20435(.A (n_7196), .Y (n_7197));
AOI21X1 g45_dup(.A0 (n_5111), .A1 (n_4714), .B0 (n_5426), .Y(n_7196));
NAND2X1 g20436(.A (n_5296), .B (n_6327), .Y (n_7198));
NAND2X1 g20437(.A (n_7195), .B (n_7198), .Y (n_7200));
AOI21X1 g20438(.A0 (n_4714), .A1 (n_5111), .B0 (n_5426), .Y (n_7201));
MX2X1 g20451(.A (n_7217), .B (n_7216), .S0 (n_7222), .Y (desOut[56]));
INVX1 g20452(.A (n_7216), .Y (n_7217));
AOI22X1 g20453(.A0 (n_3628), .A1 (n_3536), .B0 (n_3668), .B1(desIn[56]), .Y (n_7216));
NAND3X1 g20454(.A (n_7218), .B (n_7219), .C (n_7221), .Y (n_7222));
NAND2X1 g20455(.A (n_5426), .B (n_5333), .Y (n_7218));
NAND2X1 g20456(.A (n_6327), .B (n_5324), .Y (n_7219));
AOI21X1 g20457(.A0 (n_7426), .A1 (n_4462), .B0 (n_7220), .Y (n_7221));
AND2X1 g20458(.A (n_5938), .B (n_4872), .Y (n_7220));
AOI21X1 g31(.A0 (n_7224), .A1 (n_7225), .B0 (n_7231), .Y (n_7528));
OR2X1 g20459(.A (n_4199), .B (n_5089), .Y (n_7224));
NOR2X1 g20460(.A (n_7714), .B (n_7121), .Y (n_7225));
AOI21X1 g20461(.A0 (n_4649), .A1 (n_3960), .B0 (n_7227), .Y (n_7231));
INVX4 g20464(.A (n_7227), .Y (n_7228));
CLKBUFX3 g20465(.A (n_7226), .Y (n_7227));
NAND2X1 g37_dup(.A (n_3780), .B (n_3756), .Y (n_7226));
NAND2X1 g20466(.A (n_3780), .B (n_3756), .Y (n_7233));
NAND4X1 g20467(.A (n_7237), .B (n_7239), .C (n_7362), .D (n_7249), .Y(n_7250));
INVX4 g20468(.A (n_4443), .Y (n_7237));
INVX2 g20472(.A (n_7381), .Y (n_7239));
INVX1 g20478(.A (n_7248), .Y (n_7249));
CLKBUFX3 g20479(.A (n_7247), .Y (n_7248));
INVX2 g20480(.A (n_7803), .Y (n_7247));
NAND2X1 g20482(.A (n_3604), .B (desOut[3]), .Y (n_7244));
NAND2X1 g20483(.A (n_6379), .B (n_3603), .Y (n_7245));
INVX1 g20484(.A (n_7249), .Y (n_7251));
INVX1 g20485(.A (n_7247), .Y (n_7252));
INVX1 g20486(.A (n_7239), .Y (n_7253));
NAND2X1 g20520(.A (n_818), .B (n_1469), .Y (n_7284));
INVX1 g20521(.A (n_1025), .Y (n_7285));
NOR2X1 g20524(.A (n_3357), .B (n_6931), .Y (n_7289));
NOR2X1 g20525(.A (n_6355), .B (n_3358), .Y (n_7290));
NAND4X1 g20526(.A (n_7901), .B (n_7902), .C (n_7897), .D (n_7299), .Y(n_7300));
AOI21X1 g20527(.A0 (n_1661), .A1 (n_3049), .B0 (n_7294), .Y (n_7897));
AOI21X1 g20528(.A0 (n_1163), .A1 (n_2794), .B0 (n_2050), .Y (n_7294));
NAND2X2 g20529(.A (n_124), .B (n_126), .Y (n_2050));
NOR2X1 g20530(.A (n_3285), .B (n_3372), .Y (n_7901));
NOR2X1 g20531(.A (n_2999), .B (n_3067), .Y (n_7902));
NOR2X1 g20532(.A (n_7298), .B (n_2480), .Y (n_7299));
AOI21X1 g20533(.A0 (n_1724), .A1 (n_5835), .B0 (n_2907), .Y (n_7298));
INVX4 g20534(.A (n_2050), .Y (n_7301));
NAND2X2 g20535(.A (n_7303), .B (n_7307), .Y (n_7308));
NAND2X1 g20536(.A (n_2286), .B (n_7302), .Y (n_7303));
NAND4X1 g20537(.A (n_6339), .B (n_6343), .C (n_6341), .D (n_6344), .Y(n_7302));
NAND4X1 g20538(.A (n_7304), .B (n_6339), .C (n_6341), .D (desOut[7]),.Y (n_7307));
AND2X1 g20539(.A (n_6344), .B (n_6343), .Y (n_7304));
INVX1 g20540(.A (n_7305), .Y (desOut[7]));
AOI21X1 g20541(.A0 (n_717), .A1 (n_1469), .B0 (n_928), .Y (n_7305));
NAND2X1 g20542(.A (n_2286), .B (n_7302), .Y (n_7309));
INVX1 g25(.A (n_7382), .Y (n_7311));
AND2X1 g20545(.A (n_7803), .B (n_7376), .Y (n_7314));
NAND4X1 g20551(.A (n_6526), .B (n_4594), .C (n_4660), .D (n_6450), .Y(n_7317));
NAND2X1 g20552(.A (n_4635), .B (n_4049), .Y (n_7318));
INVX1 g20553(.A (n_7322), .Y (n_7323));
INVX4 g20554(.A (n_7321), .Y (n_7322));
INVX4 g20555(.A (n_7320), .Y (n_7321));
INVX2 g20556(.A (n_7319), .Y (n_7320));
MX2X1 g20557(.A (n_6978), .B (desOut[55]), .S0 (n_6980), .Y (n_7319));
NAND2X2 g20562(.A (n_7332), .B (n_7334), .Y (n_7335));
AOI21X1 g20563(.A0 (n_504), .A1 (kcy1[1]), .B0 (n_7331), .Y (n_7332));
AOI21X1 g20564(.A0 (n_280), .A1 (n_463), .B0 (n_93), .Y (n_7331));
NOR2X1 g20565(.A (n_7333), .B (n_398), .Y (n_7334));
NOR2X1 g20566(.A (n_225), .B (n_43), .Y (n_7333));
NAND4X1 g20567(.A (n_7336), .B (n_7337), .C (n_7338), .D (n_7342), .Y(n_7343));
NOR2X1 g20568(.A (n_2108), .B (n_3058), .Y (n_7336));
AOI21X1 g20569(.A0 (n_1610), .A1 (n_2744), .B0 (n_2112), .Y (n_7337));
NOR2X1 g20570(.A (n_2617), .B (n_3090), .Y (n_7338));
NAND2X1 g20571(.A (n_7339), .B (n_7341), .Y (n_7342));
NAND2X1 g20572(.A (n_1607), .B (n_2024), .Y (n_7339));
INVX4 g20573(.A (n_7340), .Y (n_7341));
NAND2X2 g20574(.A (n_124), .B (n_149), .Y (n_7340));
INVX1 g20575(.A (n_7340), .Y (n_7344));
NAND2X2 g20576(.A (n_7349), .B (n_7353), .Y (n_7354));
INVX2 g20577(.A (n_7348), .Y (n_7349));
INVX2 g20578(.A (n_7347), .Y (n_7348));
INVX2 g20579(.A (n_7346), .Y (n_7347));
INVX2 g20580(.A (n_7345), .Y (n_7346));
NAND2X2 g20581(.A (n_6832), .B (n_6833), .Y (n_7345));
NAND3X1 g20582(.A (n_7350), .B (n_7351), .C (n_7352), .Y (n_7353));
AOI22X1 g20583(.A0 (kcy3[26]), .A1 (n_573), .B0 (n_654), .B1(kcy3[26]), .Y (n_7350));
NAND2X1 g20584(.A (n_619), .B (kcy2[26]), .Y (n_7351));
NAND2X1 g20585(.A (n_485), .B (kcy1[26]), .Y (n_7352));
INVX4 g20587(.A (n_7358), .Y (n_7359));
INVX2 g20588(.A (n_7357), .Y (n_7358));
NAND2X2 g20589(.A (n_7652), .B (n_7651), .Y (n_7357));
NAND2X1 g20590(.A (n_7163), .B (desOut[11]), .Y (n_7651));
OAI21X1 g20591(.A0 (n_3593), .A1 (n_3419), .B0 (n_7161), .Y (n_7652));
NAND2X2 g20592(.A (n_7314), .B (n_7311), .Y (n_7360));
INVX4 g20593(.A (n_7359), .Y (n_7362));
NAND4X1 g20594(.A (n_7368), .B (n_7371), .C (n_7372), .D (n_7373), .Y(n_7374));
NAND3X1 g20595(.A (n_7364), .B (n_7321), .C (n_7367), .Y (n_7368));
INVX1 g20596(.A (n_7363), .Y (n_7364));
AOI21X1 g20597(.A0 (n_4245), .A1 (n_4515), .B0 (n_4228), .Y (n_7363));
MX2X1 g20598(.A (n_6579), .B (n_6580), .S0 (n_3751), .Y (n_7367));
NAND2X1 g20601(.A (n_7369), .B (n_7322), .Y (n_7371));
NAND2X1 g20602(.A (n_7318), .B (n_7317), .Y (n_7369));
NAND2X1 g20603(.A (n_4843), .B (n_7323), .Y (n_7372));
NAND2X1 g20604(.A (n_5189), .B (n_7367), .Y (n_7373));
INVX2 g20605(.A (n_7367), .Y (n_7375));
NAND2X1 g20606(.A (n_7377), .B (n_7380), .Y (n_7381));
INVX1 g20607(.A (n_7376), .Y (n_7377));
NAND2X2 g20608(.A (n_7093), .B (n_3617), .Y (n_7376));
NAND2X1 g26_dup(.A (n_7378), .B (n_7379), .Y (n_7380));
NAND4X1 g20609(.A (n_7006), .B (n_6081), .C (n_3244), .D(desOut[61]), .Y (n_7378));
NAND2X2 g20610(.A (n_7004), .B (n_1893), .Y (n_7379));
NAND2X2 g20611(.A (n_7379), .B (n_7378), .Y (n_7382));
NAND3X1 g20626(.A (n_7401), .B (n_7403), .C (n_7405), .Y (n_7406));
NOR2X1 g20627(.A (n_7400), .B (n_3406), .Y (n_7401));
NAND2X1 g20628(.A (n_6488), .B (n_7399), .Y (n_7400));
NAND2X1 g20629(.A (n_7397), .B (n_2931), .Y (n_7399));
NAND2X1 g20630(.A (n_2806), .B (n_2541), .Y (n_7397));
NOR2X1 g20632(.A (n_6486), .B (n_7402), .Y (n_7403));
OR2X1 g20633(.A (n_2507), .B (n_6491), .Y (n_7402));
INVX1 g20634(.A (n_7404), .Y (n_7405));
NAND4X1 g20635(.A (n_3204), .B (n_3114), .C (n_3112), .D (n_1869), .Y(n_7404));
NAND4X1 g47(.A (n_7407), .B (n_7408), .C (n_7410), .D (n_7411), .Y(n_7412));
NOR2X1 g20636(.A (n_3340), .B (n_3339), .Y (n_7407));
AOI21X1 g20637(.A0 (n_1984), .A1 (n_2842), .B0 (n_7026), .Y (n_7408));
NOR2X1 g20638(.A (n_7409), .B (n_2837), .Y (n_7410));
NAND2X1 g20639(.A (n_2622), .B (n_2634), .Y (n_7409));
AOI21X1 g20640(.A0 (n_1626), .A1 (n_3054), .B0 (n_7028), .Y (n_7411));
NAND3X1 g20641(.A (n_7418), .B (n_7422), .C (n_7423), .Y (n_7424));
NAND2X1 g20642(.A (n_7415), .B (n_7417), .Y (n_7418));
NAND3X1 g20643(.A (n_4181), .B (n_4207), .C (n_7414), .Y (n_7415));
INVX1 g20644(.A (n_7413), .Y (n_7414));
AND2X1 g20645(.A (n_7612), .B (n_4060), .Y (n_7413));
CLKBUFX3 g20646(.A (n_7416), .Y (n_7417));
NAND2X2 g20647(.A (n_3774), .B (n_3747), .Y (n_7416));
INVX1 g20648(.A (n_7421), .Y (n_7422));
NAND3X1 g20649(.A (n_7420), .B (n_4883), .C (n_4838), .Y (n_7421));
NOR2X1 g20650(.A (n_7419), .B (n_4620), .Y (n_7420));
NAND2X1 g20651(.A (n_4754), .B (n_4714), .Y (n_7419));
NAND2X1 g20652(.A (n_5931), .B (n_4579), .Y (n_7423));
INVX2 g20654(.A (n_7416), .Y (n_7426));
MX2X1 g20655(.A (n_7428), .B (n_7427), .S0 (n_7432), .Y (desOut[18]));
INVX1 g20656(.A (n_7427), .Y (n_7428));
AOI22X1 g20657(.A0 (desIn[18]), .A1 (n_3668), .B0 (n_3564), .B1(n_3625), .Y (n_7427));
NAND3X1 g20658(.A (n_7429), .B (n_7430), .C (n_7431), .Y (n_7432));
NAND2X1 g20659(.A (n_5445), .B (n_5331), .Y (n_7429));
NOR2X1 g20660(.A (n_5311), .B (n_5221), .Y (n_7430));
NAND2X1 g20661(.A (n_5316), .B (n_5428), .Y (n_7431));
NAND2X1 g20662(.A (n_7435), .B (n_7449), .Y (n_7450));
AOI21X1 g20663(.A0 (n_1960), .A1 (n_7301), .B0 (n_7434), .Y (n_7435));
AOI21X1 g20664(.A0 (n_3104), .A1 (n_3117), .B0 (n_2907), .Y (n_7434));
AOI21X1 g20665(.A0 (n_1548), .A1 (n_3159), .B0 (n_7448), .Y (n_7449));
NOR2X1 g20666(.A (n_7437), .B (n_7447), .Y (n_7448));
INVX1 g20669(.A (n_7436), .Y (n_7437));
AND2X1 g20670(.A (n_132), .B (n_126), .Y (n_7436));
AND2X1 g20671(.A (n_7442), .B (n_7446), .Y (n_7447));
INVX1 g20673(.A (n_7442), .Y (n_7443));
INVX2 g20674(.A (n_7441), .Y (n_7442));
INVX2 g20675(.A (n_7440), .Y (n_7441));
NAND2X1 g20676(.A (n_767), .B (n_884), .Y (n_7440));
CLKBUFX3 g20677(.A (n_7445), .Y (n_7446));
NAND2X2 g20678(.A (n_779), .B (n_790), .Y (n_7445));
INVX1 g20679(.A (n_7443), .Y (n_7451));
MX2X1 g20681(.A (n_7453), .B (n_7454), .S0 (n_7455), .Y (desOut[4]));
OAI21X1 g20682(.A0 (n_3483), .A1 (n_3677), .B0 (n_7095), .Y (n_7453));
INVX1 g20683(.A (n_7453), .Y (n_7454));
NAND3X1 g20684(.A (n_7905), .B (n_7906), .C (n_6212), .Y (n_7455));
AOI21X1 g20685(.A0 (n_7465), .A1 (n_7466), .B0 (n_7469), .Y (n_7470));
INVX2 g20686(.A (n_7464), .Y (n_7465));
INVX4 g20687(.A (n_7463), .Y (n_7464));
INVX4 g20688(.A (n_7462), .Y (n_7463));
INVX2 g20689(.A (n_7461), .Y (n_7462));
MX2X1 g20690(.A (n_7458), .B (desOut[19]), .S0 (n_7460), .Y (n_7461));
OAI22X1 g20691(.A0 (n_1030), .A1 (n_701), .B0 (n_879), .B1(desIn[19]), .Y (n_7458));
NOR2X1 g20694(.A (n_3425), .B (n_7412), .Y (n_7460));
INVX1 g20696(.A (n_7466), .Y (n_7467));
NOR2X1 g20697(.A (n_7360), .B (n_7359), .Y (n_7466));
NAND2X1 g20698(.A (n_4957), .B (n_4858), .Y (n_7469));
NAND2X1 g20707(.A (n_7479), .B (n_7488), .Y (n_7489));
NOR2X1 g20708(.A (n_4055), .B (n_4044), .Y (n_7479));
CLKBUFX1 g20709(.A (n_7487), .Y (n_7488));
NAND2X2 g20710(.A (n_7483), .B (n_7486), .Y (n_7487));
OAI21X1 g20711(.A0 (n_7480), .A1 (n_7481), .B0 (desOut[15]), .Y(n_7483));
NAND2X1 g20712(.A (n_7290), .B (n_7807), .Y (n_7480));
INVX1 g20713(.A (n_7289), .Y (n_7481));
NAND2X1 g20714(.A (n_7284), .B (n_7285), .Y (desOut[15]));
NAND4X1 g20715(.A (n_7289), .B (n_7808), .C (n_7290), .D (n_7485), .Y(n_7486));
INVX1 g20717(.A (desOut[15]), .Y (n_7485));
INVX1 g20718(.A (n_7488), .Y (n_7490));
INVX1 g20719(.A (n_7488), .Y (n_7491));
INVX4 g20720(.A (n_7487), .Y (n_7492));
NAND4X1 g20721(.A (n_7493), .B (n_7495), .C (n_7497), .D (n_7500), .Y(n_7501));
NOR2X1 g20722(.A (n_2446), .B (n_3047), .Y (n_7493));
NOR2X1 g20723(.A (n_2997), .B (n_7494), .Y (n_7495));
INVX1 g20724(.A (n_2864), .Y (n_7494));
AOI21X1 g20725(.A0 (n_2800), .A1 (n_2402), .B0 (n_7496), .Y (n_7497));
NAND2X1 g20726(.A (n_2865), .B (n_2448), .Y (n_7496));
NOR2X1 g20727(.A (n_7498), .B (n_7499), .Y (n_7500));
NAND2X1 g20728(.A (n_2227), .B (n_1820), .Y (n_7498));
INVX1 g20729(.A (n_2447), .Y (n_7499));
AOI21X1 g20730(.A0 (n_7509), .A1 (kcy2[4]), .B0 (n_7510), .Y(n_7511));
NAND2X1 g20731(.A (n_7505), .B (n_7508), .Y (n_7509));
INVX2 g20732(.A (n_7504), .Y (n_7505));
INVX2 g20733(.A (n_7503), .Y (n_7504));
INVX4 g20734(.A (n_7502), .Y (n_7503));
NOR2X1 g20735(.A (n_7129), .B (n_6130), .Y (n_7502));
INVX1 g20736(.A (n_7507), .Y (n_7508));
INVX2 g20737(.A (n_7506), .Y (n_7507));
NAND3X1 g20738(.A (n_102), .B (n_7128), .C (roundSel[4]), .Y(n_7506));
NOR2X1 g20739(.A (n_81), .B (n_248), .Y (n_7510));
OAI22X1 g20741(.A0 (n_1776), .A1 (n_70), .B0 (n_3552), .B1 (n_3677),.Y (n_7512));
INVX1 g20742(.A (n_7512), .Y (n_7513));
NAND4X1 g20743(.A (n_7793), .B (n_7794), .C (n_7516), .D (n_7517), .Y(n_7518));
NOR2X1 g20744(.A (n_6192), .B (n_5039), .Y (n_7794));
NAND2X1 g20745(.A (n_6199), .B (n_7121), .Y (n_7793));
OAI21X1 g20746(.A0 (n_6136), .A1 (n_6137), .B0 (n_6195), .Y (n_7516));
NAND3X1 g20747(.A (n_5010), .B (n_4133), .C (n_4413), .Y (n_7517));
NAND2X2 g20748(.A (n_5532), .B (n_5543), .Y (desOut[36]));
NAND2X1 g13525_dup(.A (n_5532), .B (n_5543), .Y (n_7546));
INVX4 g20758(.A (n_7568), .Y (n_7559));
CLKBUFX2 g20761(.A (n_7559), .Y (n_7563));
INVX2 g20765(.A (n_859), .Y (n_7568));
INVX2 g20775(.A (n_7603), .Y (n_7604));
CLKBUFX3 g20776(.A (n_6935), .Y (n_7603));
INVX1 g20777(.A (n_7606), .Y (n_7605));
CLKBUFX1 g20778(.A (n_7607), .Y (n_7606));
INVX1 g20779(.A (n_7607), .Y (n_7608));
INVX1 g20780(.A (n_7615), .Y (n_7607));
INVX1 g20783(.A (n_7614), .Y (n_7612));
CLKBUFX1 g20784(.A (n_7615), .Y (n_7614));
MX2X1 g20794(.A (n_6481), .B (n_6480), .S0 (n_6972), .Y (desOut[62]));
MX2X1 g19756_dup(.A (n_6481), .B (n_6480), .S0 (n_6972), .Y (n_7627));
MX2X1 g20796(.A (n_6278), .B (n_6277), .S0 (n_6279), .Y (desOut[20]));
MX2X1 g19574_dup(.A (n_6278), .B (n_6277), .S0 (n_6279), .Y (n_7631));
NAND2X1 g20797(.A (n_742), .B (n_766), .Y (n_7632));
NAND2X1 g17738_dup(.A (n_742), .B (n_766), .Y (n_7633));
NAND2X1 g20798(.A (n_899), .B (n_887), .Y (n_7634));
NAND2X1 g17378_dup(.A (n_899), .B (n_887), .Y (n_7635));
NAND2X1 g20799(.A (n_793), .B (n_790), .Y (n_7636));
NAND2X1 g17444_dup(.A (n_793), .B (n_790), .Y (n_7637));
NAND2X1 g20809(.A (n_877), .B (n_815), .Y (n_7655));
NAND2X1 g17161_dup(.A (n_877), .B (n_815), .Y (n_7656));
CLKBUFX3 g17726_dup(.A (n_914), .Y (n_2068));
NAND2X1 g20811(.A (n_7158), .B (n_5480), .Y (desOut[10]));
NAND2X2 g13583_dup(.A (n_7158), .B (n_5480), .Y (n_7660));
NAND2X1 g20812(.A (n_7043), .B (n_5655), .Y (n_7661));
NAND2X1 g17939_dup(.A (n_7043), .B (n_5655), .Y (n_7662));
NAND2X1 g20813(.A (n_865), .B (n_864), .Y (n_7663));
NAND2X2 g17395_dup(.A (n_865), .B (n_864), .Y (n_7664));
NAND2X1 g20822(.A (n_2839), .B (n_1677), .Y (n_7683));
NAND2X1 g16939_dup(.A (n_2839), .B (n_1677), .Y (n_7684));
NAND2X1 g20823(.A (n_888), .B (n_887), .Y (n_7685));
NAND2X2 g17613_dup(.A (n_888), .B (n_887), .Y (n_7686));
MX2X1 g20824(.A (n_7512), .B (n_7513), .S0 (n_7518), .Y (desOut[58]));
MX2X1 g20740_dup(.A (n_7512), .B (n_7513), .S0 (n_7518), .Y (n_7688));
NAND2X1 g20834(.A (n_869), .B (n_7348), .Y (n_7700));
NAND2X1 g17341_dup(.A (n_869), .B (n_7348), .Y (n_7701));
NAND2X2 g20835(.A (n_6643), .B (n_6648), .Y (n_7702));
NAND2X2 g19914_dup(.A (n_6643), .B (n_6648), .Y (n_1495));
NAND2X1 g20836(.A (n_785), .B (n_784), .Y (n_7704));
NAND2X1 g17426_dup(.A (n_785), .B (n_784), .Y (n_7705));
NAND2X1 g20837(.A (n_6944), .B (n_6940), .Y (n_7706));
NAND2X1 g20183_dup(.A (n_6944), .B (n_6940), .Y (n_7707));
INVX2 g20838(.A (n_7714), .Y (n_7709));
INVX1 g20840(.A (n_7711), .Y (n_7712));
CLKBUFX3 g20842(.A (n_7711), .Y (n_7714));
INVX1 g20843(.A (n_7233), .Y (n_7711));
CLKBUFX1 g20854(.A (n_7733), .Y (n_7728));
CLKBUFX1 g20857(.A (n_7733), .Y (n_7732));
INVX1 g20860(.A (n_7735), .Y (n_7738));
INVX2 g20861(.A (n_4255), .Y (n_7735));
CLKBUFX1 g20862(.A (n_7741), .Y (n_7740));
NAND2X1 g20881(.A (n_7244), .B (n_7245), .Y (n_7803));
NAND2X1 g24_dup(.A (n_7244), .B (n_7245), .Y (n_7804));
INVX4 g20882(.A (n_6564), .Y (n_7805));
INVX4 g19840_dup(.A (n_6564), .Y (n_7806));
NOR2X1 g20883(.A (n_6930), .B (n_6352), .Y (n_7807));
NOR2X1 g20523_dup(.A (n_6930), .B (n_6352), .Y (n_7808));
INVX1 g20886(.A (n_7813), .Y (n_7812));
INVX4 g20888(.A (n_7816), .Y (n_7813));
INVX1 g20889(.A (n_7816), .Y (n_7815));
INVX2 g20890(.A (n_7820), .Y (n_7816));
CLKBUFX3 g20893(.A (n_7820), .Y (n_7819));
INVX2 g20894(.A (n_7857), .Y (n_7820));
INVX1 g20895(.A (n_7857), .Y (n_7821));
INVX4 g20898(.A (n_7854), .Y (n_7824));
INVX2 g20913(.A (n_7854), .Y (n_7846));
CLKBUFX3 g20921(.A (n_7857), .Y (n_7854));
INVX1 g20922(.A (n_7858), .Y (n_7859));
INVX4 g20924(.A (n_7857), .Y (n_7858));
INVX4 g20925(.A (n_7871), .Y (n_7857));
INVX1 g20931(.A (n_7869), .Y (n_7867));
CLKBUFX2 g20933(.A (n_7857), .Y (n_7869));
INVX2 g20935(.A (n_296), .Y (n_7871));
endmodule
