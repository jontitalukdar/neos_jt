module s15850(blif_clk_net, blif_reset_net, g18, g27, g109, g741,g742, g743, g744, g872, g873, g877, g881, g1712, g1960, g1961,g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608,g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172,g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181,g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926,g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313,g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349,g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977,g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986,g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461,g10463, g10465, g10628, g10801, g11163, g11206, g11489);
input blif_clk_net, blif_reset_net, g18, g27, g109, g741, g742, g743,g744, g872, g873, g877, g881, g1712, g1960, g1961;
output g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608,g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172,g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181,g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926,g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313,g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349,g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977,g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986,g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461,g10463, g10465, g10628, g10801, g11163, g11206, g11489;
wire blif_clk_net, blif_reset_net, g18, g27, g109, g741, g742, g743,g744, g872, g873, g877, g881, g1712, g1960, g1961;
wire g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608,g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172,g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181,g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926,g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313,g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349,g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977,g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986,g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461,g10463, g10465, g10628, g10801, g11163, g11206, g11489;
wire g253, g254, g255, g256, g257, g258, g259, g260;
wire g261, g262, g305, g309, g312, g315, g318, g321;
wire g324, g327, g330, g333, g369, g374, g378, g382;
wire g431, g590, g757, g869, g876, g882, g928, g932;
wire g936, g940, g971, g976, g981, g986, g1104, g1107;
wire g1110, g1113, g1117, g1121, g1125, g1129, g1133, g1137;
wire g1141, g1145, g1149, g1153, g1157, g1160, g1163, g1166;
wire g1212, g1216, g1218, g1223, g1227, g1231, g1235, g1240;
wire g1245, g1255, g1260, g1265, g1270, g1275, g1280, g1284;
wire g1289, g1292, g1296, g1300, g1304, g1336, g1341, g1346;
wire g1351, g1361, g1362, g1365, g1368, g1371, g1374, g1377;
wire g1380, g1383, g1386, g1389, g1397, g1400, g1512, g1615;
wire g1618, g1621, g1624, g1627, g1630, g1633, g1636, g1639;
wire g1710, g1713, g1718, g_1292, g_1295, g_1298, g_1301, g_1304;
wire g_1307, g_1325, g_1328, g_1331, g_1334, g_1340, g_1343, g_1346;
wire g_2336, g_2705, g_3128, g_3811, g_6600, g_7025, g_7375, g_7720;
wire g_8244, g_8484, g_8701, g_9187, g_9394, g_9514, g_9904, g_10008;
wire g_10087, g_10548, g_10572, g_10698, g_10714, g_10749, g_10855,g_10859;
wire gbuf5, gbuf6, gbuf12, gbuf13, n_1, n_5, n_6, n_9;
wire n_10, n_12, n_13, n_15, n_16, n_17, n_19, n_20;
wire n_22, n_24, n_25, n_26, n_27, n_28, n_29, n_30;
wire n_32, n_34, n_36, n_37, n_38, n_39, n_40, n_42;
wire n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51;
wire n_52, n_53, n_55, n_58, n_59, n_61, n_62, n_69;
wire n_70, n_76, n_77, n_78, n_79, n_80, n_81, n_83;
wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_98;
wire n_99, n_112, n_115, n_116, n_117, n_118, n_119, n_120;
wire n_122, n_123, n_124, n_127, n_128, n_129, n_130, n_131;
wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
wire n_140, n_141, n_143, n_144, n_145, n_146, n_148, n_149;
wire n_150, n_151, n_152, n_153, n_154, n_159, n_160, n_161;
wire n_162, n_165, n_167, n_168, n_169, n_170, n_171, n_172;
wire n_173, n_174, n_176, n_177, n_178, n_184, n_187, n_188;
wire n_189, n_193, n_194, n_196, n_197, n_198, n_199, n_200;
wire n_201, n_202, n_203, n_204, n_205, n_207, n_208, n_209;
wire n_210, n_211, n_212, n_213, n_214, n_215, n_217, n_218;
wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
wire n_235, n_238, n_243, n_244, n_246, n_247, n_248, n_249;
wire n_251, n_252, n_253, n_254, n_257, n_258, n_259, n_260;
wire n_261, n_262, n_263, n_264, n_265, n_266, n_268, n_269;
wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
wire n_278, n_279, n_280, n_281, n_282, n_284, n_285, n_286;
wire n_287, n_288, n_295, n_297, n_299, n_300, n_301, n_302;
wire n_303, n_304, n_305, n_306, n_307, n_309, n_310, n_311;
wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
wire n_337, n_338, n_339, n_340, n_342, n_343, n_344, n_345;
wire n_346, n_347, n_348, n_349, n_350, n_353, n_354, n_356;
wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_382;
wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
wire n_391, n_392, n_394, n_395, n_396, n_397, n_398, n_399;
wire n_400, n_401, n_402, n_405, n_406, n_409, n_410, n_411;
wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
wire n_420, n_421, n_422, n_423, n_425, n_426, n_427, n_429;
wire n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437;
wire n_438, n_439, n_440, n_441, n_442, n_445, n_446, n_447;
wire n_448, n_449, n_451, n_453, n_454, n_455, n_457, n_458;
wire n_459, n_461, n_463, n_464, n_465, n_466, n_469, n_470;
wire n_471, n_474, n_475, n_476, n_477, n_479, n_481, n_483;
wire n_485, n_486, n_500, n_503, n_518, n_520, n_523, n_526;
wire n_528, n_530, n_531, n_532, n_533, n_543, n_544, n_551;
wire n_576, n_584, n_585, n_586, n_587, n_588, n_589, n_593;
wire n_594, n_595, n_596, n_597, n_598, n_600, n_606, n_608;
wire n_641, n_642, n_660, n_661, n_664, n_665, n_671, n_676;
wire n_679, n_680, n_681, n_682, n_686, n_689, n_690, n_694;
wire n_695, n_697, n_700, n_710, n_711, n_712, n_713, n_718;
wire n_722, n_730, n_735, n_736, n_737, n_738, n_739, n_740;
wire n_741, n_742, n_744, n_747, n_748, n_749, n_750, n_751;
wire n_754, n_756, n_762, n_763, n_764, n_765, n_773, n_792;
wire n_793, n_797, n_798, n_799, n_800, n_802, n_803, n_804;
wire n_805, n_806, n_807, n_808, n_809, n_814, n_815, n_816;
wire n_818, n_819, n_820, n_823, n_826, n_827, n_828, n_829;
wire n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839;
wire n_840, n_841, n_846, n_849, n_850, n_852, n_853, n_854;
wire n_859, n_861, n_862, n_863, n_864, n_865, n_869, n_870;
wire n_885, n_891, n_892, n_893, n_900, n_912, n_913, n_915;
wire n_916, n_918, n_923, n_924, n_925, n_926, n_927, n_928;
wire n_929, n_930, n_931, n_932, n_933, n_934, n_935, n_936;
wire n_937, n_938, n_939, n_940, n_941, n_942, n_944, n_945;
wire n_946, n_947, n_948, n_949, n_950, n_951;
assign g11489 = 1'b0;
assign g11206 = 1'b1;
assign g10801 = 1'b1;
assign g10628 = 1'b1;
assign g10465 = 1'b1;
assign g10463 = 1'b1;
assign g10461 = 1'b1;
assign g10459 = 1'b1;
assign g10457 = 1'b1;
assign g10455 = 1'b1;
assign g10379 = 1'b1;
assign g10377 = 1'b1;
assign g9961 = 1'b0;
assign g9451 = 1'b0;
assign g8986 = 1'b0;
assign g8985 = 1'b0;
assign g8984 = 1'b0;
assign g8983 = 1'b0;
assign g8982 = 1'b0;
assign g8981 = 1'b0;
assign g8980 = 1'b0;
assign g8979 = 1'b0;
assign g8978 = 1'b0;
assign g8977 = 1'b0;
assign g8976 = 1'b0;
assign g8566 = 1'b0;
assign g8565 = 1'b0;
assign g8564 = 1'b0;
assign g8563 = 1'b0;
assign g8562 = 1'b0;
assign g8561 = 1'b0;
assign g8352 = 1'b0;
assign g8349 = 1'b0;
assign g8347 = 1'b0;
assign g8340 = 1'b0;
assign g8335 = 1'b0;
assign g8331 = 1'b0;
assign g8328 = 1'b0;
assign g8323 = 1'b0;
assign g8318 = 1'b0;
assign g8316 = 1'b0;
assign g8313 = 1'b0;
assign g8271 = 1'b1;
assign g8062 = g873;
assign g8061 = g872;
assign g7744 = g27;
assign g6955 = 1'b0;
assign g6949 = 1'b0;
assign g6942 = 1'b0;
assign g6932 = 1'b0;
assign g6926 = 1'b0;
assign g6920 = 1'b0;
assign g5816 = 1'b1;
assign g5105 = g873;
assign g5101 = g872;
assign g4888 = g1960;
assign g4887 = g1961;
assign g4172 = 1'b0;
assign g2612 = 1'b0;
assign g2611 = 1'b0;
assign g2610 = 1'b0;
assign g2609 = 1'b0;
assign g2608 = 1'b0;
assign g2607 = 1'b0;
assign g2606 = 1'b0;
assign g2605 = 1'b0;
assign g2604 = 1'b0;
assign g2603 = 1'b0;
assign g2602 = 1'b0;
assign g2601 = 1'b0;
assign g2355 = g18;
DFFSRX1 g976_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_532), .Q (), .QN (g976));
DFFSRX1 g981_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_531), .Q (), .QN (g981));
DFFSRX1 g986_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_530), .Q (), .QN (g986));
NAND2X2 g21280(.A (n_523), .B (n_589), .Y (n_532));
DFFSRX1 g971_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_840), .Q (g971), .QN ());
NAND2X2 g21281(.A (n_520), .B (n_765), .Y (n_531));
NAND2X2 g21282(.A (n_528), .B (n_526), .Y (n_530));
NAND3X1 g21287(.A (n_543), .B (n_773), .C (n_342), .Y (n_528));
NAND3X1 g21288(.A (n_344), .B (n_763), .C (n_773), .Y (n_526));
NAND3X1 g21289(.A (n_543), .B (n_773), .C (n_124), .Y (n_523));
NAND3X1 g21285(.A (n_543), .B (n_773), .C (n_235), .Y (n_520));
NAND3X1 g21293(.A (n_93), .B (g757), .C (g869), .Y (n_518));
DFFSRX1 g757_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_544), .Q (), .QN (g757));
DFFSRX1 g1341_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_939), .Q (), .QN (g1341));
DFFSRX1 g1346_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_503), .Q (), .QN (g1346));
DFFSRX1 g1351_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_500), .Q (), .QN (g1351));
DFFSRX1 g426_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_551), .Q (g_1325), .QN ());
OAI33X1 g21420(.A0 (n_937), .A1 (n_120), .A2 (n_160), .B0 (n_464),.B1 (n_927), .B2 (g1346), .Y (n_503));
OAI33X1 g21421(.A0 (n_937), .A1 (n_161), .A2 (n_224), .B0 (n_466),.B1 (n_927), .B2 (g1351), .Y (n_500));
DFFSRX1 g1336_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_865), .Q (), .QN (g1336));
DFFSRX1 g305_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g253), .Q (g305), .QN ());
DFFSRX1 g201_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_483), .Q (g_10749), .QN ());
DFFSRX1 g253_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_477), .Q (g253), .QN ());
AOI21X1 g21452(.A0 (g1361), .A1 (g3069), .B0 (n_476), .Y (n_486));
NOR2X1 g21326(.A (g321), .B (n_735), .Y (n_485));
AND2X1 g21307(.A (n_474), .B (n_232), .Y (n_483));
NOR2X1 g21311(.A (g318), .B (n_737), .Y (n_481));
NOR2X1 g21366(.A (g327), .B (n_944), .Y (n_479));
OAI21X1 g21333(.A0 (g_9904), .A1 (g18), .B0 (n_458), .Y (n_477));
DFFSRX1 g318_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g257), .Q (), .QN (g318));
NAND2X1 g21460(.A (g_3811), .B (g1212), .Y (n_476));
DFFSRX1 g321_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g258), .Q (), .QN (g321));
DFFSRX1 g330_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g261), .Q (), .QN (g330));
AOI21X1 g21335(.A0 (g315), .A1 (n_122), .B0 (n_471), .Y (n_475));
DFFSRX1 g333_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g262), .Q (), .QN (g333));
XOR2X1 g21312(.A (n_447), .B (n_470), .Y (n_474));
DFFSRX1 g309_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g254), .Q (), .QN (g309));
DFFSRX1 g327_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g260), .Q (), .QN (g327));
DFFSRX1 g324_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g259), .Q (), .QN (g324));
DFFSRX1 g257_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_469), .Q (g257), .QN ());
DFFSRX1 g108_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_465), .Q (), .QN (g_3811));
DFFSRX1 g258_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_461), .Q (g258), .QN ());
DFFSRX1 g261_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_463), .Q (g261), .QN ());
NOR2X1 g21337(.A (g315), .B (n_122), .Y (n_471));
DFFSRX1 g262_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_457), .Q (g262), .QN ());
DFFSRX1 g546_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_459), .Q (), .QN (g_9904));
DFFSRX1 g259_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_455), .Q (g259), .QN ());
NOR2X1 g21318(.A (n_197), .B (n_453), .Y (n_470));
DFFSRX1 g254_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_454), .Q (g254), .QN ());
DFFSRX1 g260_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_451), .Q (g260), .QN ());
OAI21X1 g21322(.A0 (g_10008), .A1 (g18), .B0 (n_438), .Y (n_469));
INVX1 g21472(.A (n_932), .Y (n_466));
INVX1 g21473(.A (n_932), .Y (n_465));
INVX1 g21474(.A (n_932), .Y (n_464));
DFFSRX1 g312_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g255), .Q (), .QN (g312));
OAI21X1 g21396(.A0 (g_9394), .A1 (g18), .B0 (n_434), .Y (n_463));
OAI21X1 g21338(.A0 (g_8244), .A1 (g18), .B0 (n_441), .Y (n_461));
DFFSRX1 g315_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g256), .Q (g315), .QN ());
AOI21X1 g21350(.A0 (n_449), .A1 (n_458), .B0 (g1718), .Y (n_459));
OAI21X1 g21424(.A0 (g_7375), .A1 (g18), .B0 (n_422), .Y (n_457));
OAI21X1 g21359(.A0 (g_3128), .A1 (g18), .B0 (n_431), .Y (n_455));
OAI21X1 g21459(.A0 (g_10855), .A1 (g18), .B0 (n_429), .Y (n_454));
OR4X1 g21323(.A (g1374), .B (n_446), .C (g_9187), .D (g1397), .Y(n_453));
OAI21X1 g21381(.A0 (g_2336), .A1 (g18), .B0 (n_426), .Y (n_451));
DFFSRX1 g865_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_681), .Q (g2648), .QN ());
DFFSRX1 g255_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_445), .Q (g255), .QN ());
DFFSRX1 g256_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_448), .Q (g256), .QN ());
DFFSRX1 g572_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_440), .Q (), .QN (g_7375));
DFFSRX1 g790_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_436), .Q (g4181), .QN ());
DFFSRX1 g1275_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_437), .Q (g1275), .QN ());
DFFSRX1 g557_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_439), .Q (), .QN (g_10008));
OR2X1 g21497(.A (g1618), .B (g18), .Y (n_449));
DFFSRX1 g569_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_435), .Q (), .QN (g_9394));
DFFSRX1 g560_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_442), .Q (), .QN (g_8244));
OAI21X1 g21355(.A0 (g_6600), .A1 (g18), .B0 (n_354), .Y (n_448));
DFFSRX1 g786_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_433), .Q (g4180), .QN ());
DFFSRX1 g563_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_432), .Q (), .QN (g_3128));
DFFSRX1 g575_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_430), .Q (), .QN (g_10855));
XOR2X1 g21327(.A (g_10749), .B (n_421), .Y (n_447));
NAND4X1 g21331(.A (g1400), .B (n_418), .C (n_22), .D (n_20), .Y(n_446));
DFFSRX1 g566_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_427), .Q (), .QN (g_2336));
OAI21X1 g21524(.A0 (g_8701), .A1 (g18), .B0 (n_345), .Y (n_445));
AOI21X1 g21356(.A0 (n_415), .A1 (n_441), .B0 (g1718), .Y (n_442));
OR2X1 g21450(.A (n_423), .B (g1718), .Y (n_440));
DFFSRX1 g1618_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_419), .Q (), .QN (g1618));
AOI21X1 g21334(.A0 (n_406), .A1 (n_438), .B0 (g1718), .Y (n_439));
NAND2X1 g21515(.A (n_420), .B (n_297), .Y (n_437));
NOR2X1 g21412(.A (n_425), .B (n_269), .Y (n_436));
AOI21X1 g21419(.A0 (n_417), .A1 (n_434), .B0 (g1718), .Y (n_435));
NOR2X1 g21437(.A (n_416), .B (n_269), .Y (n_433));
DFFSRX1 g1227_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_411), .Q (g1227), .QN ());
DFFSRX1 g1218_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_414), .Q (g1218), .QN ());
DFFSRX1 g1231_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_409), .Q (g1231), .QN ());
DFFSRX1 g1223_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_413), .Q (g1223), .QN ());
AOI21X1 g21378(.A0 (n_400), .A1 (n_431), .B0 (g1718), .Y (n_432));
NAND2X1 g21486(.A (n_412), .B (n_429), .Y (n_430));
AOI21X1 g21394(.A0 (n_395), .A1 (n_426), .B0 (g1718), .Y (n_427));
XOR2X1 g21428(.A (g4181), .B (n_682), .Y (n_425));
DFFSRX1 g554_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_401), .Q (), .QN (g_6600));
DFFSRX1 g782_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_402), .Q (g4179), .QN ());
DFFSRX1 g374_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_399), .Q (g374), .QN ());
DFFSRX1 g378_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_398), .Q (g378), .QN ());
DFFSRX1 g382_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_396), .Q (g382), .QN ());
OAI21X1 g21456(.A0 (g1633), .A1 (g18), .B0 (n_422), .Y (n_423));
DFFSRX1 g762_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_405), .Q (g4174), .QN ());
XOR2X1 g21336(.A (g_2705), .B (n_380), .Y (n_421));
NAND2X1 g21521(.A (n_394), .B (n_338), .Y (n_420));
XOR2X1 g21525(.A (n_99), .B (n_382), .Y (n_419));
NOR2X1 g21339(.A (n_392), .B (g1380), .Y (n_418));
DFFSRX1 g549_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_391), .Q (), .QN (g_8701));
OR2X1 g21436(.A (g1630), .B (g18), .Y (n_417));
XOR2X1 g21453(.A (g4180), .B (n_358), .Y (n_416));
OR2X1 g21365(.A (g1621), .B (g18), .Y (n_415));
DFFSRX1 g778_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_390), .Q (g4178), .QN ());
DFFSRX1 g928_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_378), .Q (), .QN (g928));
DFFSRX1 g932_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_376), .Q (), .QN (g932));
DFFSRX1 g936_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_379), .Q (), .QN (g936));
DFFSRX1 g940_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_375), .Q (), .QN (g940));
DFFSRX1 g369_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_389), .Q (g369), .QN ());
NOR2X1 g21499(.A (n_383), .B (n_225), .Y (n_414));
OAI21X1 g21500(.A0 (n_167), .A1 (n_410), .B0 (n_388), .Y (n_413));
AOI21X1 g21501(.A0 (g1636), .A1 (n_81), .B0 (g1718), .Y (n_412));
OAI21X1 g21502(.A0 (n_248), .A1 (n_410), .B0 (n_387), .Y (n_411));
OAI21X1 g21503(.A0 (n_280), .A1 (n_410), .B0 (n_384), .Y (n_409));
OR2X1 g21343(.A (g1615), .B (g18), .Y (n_406));
NAND2X1 g21593(.A (n_374), .B (n_310), .Y (n_405));
DFFSRX1 g1270_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_366), .Q (g1270), .QN ());
DFFSRX1 g1296_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_362), .Q (g1296), .QN ());
DFFSRX1 g774_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_350), .Q (g4177), .QN ());
DFFSRX1 g878_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_343), .Q (g3007), .QN ());
DFFSRX1 g770_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_349), .Q (g4176), .QN ());
DFFSRX1 g1235_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_373), .Q (g1235), .QN ());
DFFSRX1 g1245_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_371), .Q (g1245), .QN ());
DFFSRX1 g1255_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_369), .Q (g1255), .QN ());
DFFSRX1 g1265_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_367), .Q (g1265), .QN ());
DFFSRX1 g1280_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_365), .Q (g1280), .QN ());
DFFSRX1 g1284_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_364), .Q (g1284), .QN ());
DFFSRX1 g1292_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_363), .Q (g1292), .QN ());
NOR2X1 g21457(.A (n_353), .B (n_269), .Y (n_402));
DFFSRX1 g1300_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_361), .Q (g1300), .QN ());
DFFSRX1 g766_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_359), .Q (g4175), .QN ());
OR2X1 g21371(.A (n_356), .B (g1718), .Y (n_401));
DFFSRX1 g1260_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_368), .Q (g1260), .QN ());
DFFSRX1 g1250_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_370), .Q (n_330), .QN ());
OR2X1 g21386(.A (g1624), .B (g18), .Y (n_400));
AOI21X1 g21509(.A0 (n_287), .A1 (n_302), .B0 (n_397), .Y (n_399));
AOI21X1 g21510(.A0 (n_285), .A1 (n_301), .B0 (n_397), .Y (n_398));
AOI21X1 g21511(.A0 (n_284), .A1 (n_299), .B0 (n_397), .Y (n_396));
OR2X1 g21404(.A (g1627), .B (g18), .Y (n_395));
INVX1 g21539(.A (n_940), .Y (n_394));
DFFSRX1 g1304_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_360), .Q (g1304), .QN ());
DFFSRX1 g1240_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_372), .Q (g1240), .QN ());
NAND4X1 g21344(.A (n_347), .B (g1377), .C (n_15), .D (n_12), .Y(n_392));
OR2X1 g21563(.A (n_346), .B (g1718), .Y (n_391));
DFFSRX1 g1630_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_316), .Q (), .QN (g1630));
DFFSRX1 g1621_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_309), .Q (), .QN (g1621));
DFFSRX1 g1633_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_307), .Q (), .QN (g1633));
NOR2X1 g21487(.A (n_304), .B (n_269), .Y (n_390));
NOR2X1 g21508(.A (n_303), .B (n_397), .Y (n_389));
NAND3X1 g21512(.A (n_386), .B (n_385), .C (n_165), .Y (n_388));
NAND3X1 g21513(.A (n_386), .B (n_385), .C (n_247), .Y (n_387));
NAND3X1 g21514(.A (n_386), .B (n_385), .C (g1231), .Y (n_384));
XOR2X1 g21517(.A (n_596), .B (n_385), .Y (n_383));
XOR2X1 g21553(.A (n_140), .B (n_279), .Y (n_382));
XOR2X1 g21345(.A (g1386), .B (g1389), .Y (n_380));
DFFSRX1 g1615_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_340), .Q (), .QN (g1615));
NOR2X1 g21585(.A (n_377), .B (g936), .Y (n_379));
NOR2X1 g21586(.A (n_377), .B (g928), .Y (n_378));
NOR2X1 g21587(.A (n_377), .B (g932), .Y (n_376));
NOR2X1 g21588(.A (n_377), .B (g940), .Y (n_375));
NAND2X1 g21598(.A (n_348), .B (g4174), .Y (n_374));
INVX1 g21600(.A (n_339), .Y (n_373));
INVX1 g21602(.A (n_337), .Y (n_372));
INVX1 g21604(.A (n_334), .Y (n_371));
INVX1 g21606(.A (n_332), .Y (n_370));
INVX1 g21608(.A (n_331), .Y (n_369));
INVX1 g21610(.A (n_329), .Y (n_368));
INVX1 g21612(.A (n_327), .Y (n_367));
INVX1 g21614(.A (n_325), .Y (n_366));
INVX1 g21616(.A (n_323), .Y (n_365));
INVX1 g21618(.A (n_322), .Y (n_364));
INVX1 g21620(.A (n_320), .Y (n_363));
INVX1 g21622(.A (n_318), .Y (n_362));
INVX1 g21624(.A (n_315), .Y (n_361));
INVX1 g21626(.A (n_313), .Y (n_360));
NOR2X1 g21642(.A (n_152), .B (n_269), .Y (n_359));
INVX1 g21466(.A (n_711), .Y (n_358));
OAI21X1 g21376(.A0 (g1639), .A1 (g18), .B0 (n_354), .Y (n_356));
XOR2X1 g21478(.A (g4179), .B (n_713), .Y (n_353));
DFFSRX1 g1624_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_288), .Q (), .QN (g1624));
INVX1 g21734(.A (n_306), .Y (g5658));
INVX1 g21744(.A (n_305), .Y (g5659));
DFFSRX1 g1636_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_282), .Q (g1636), .QN ());
NOR2X1 g21520(.A (n_243), .B (n_269), .Y (n_350));
OR2X1 g21522(.A (n_225), .B (n_385), .Y (n_410));
DFFSRX1 g1627_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_281), .Q (), .QN (g1627));
NOR2X1 g21562(.A (n_234), .B (n_269), .Y (n_349));
DFFSRX1 g758_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_348), .Q (g4173), .QN ());
NOR2X1 g21351(.A (g1383), .B (g1386), .Y (n_347));
OAI21X1 g21590(.A0 (g1512), .A1 (g18), .B0 (n_345), .Y (n_346));
AND2X1 g21550(.A (n_606), .B (n_342), .Y (n_343));
XOR2X1 g21550_xor(.A (n_606), .B (n_342), .Y (n_344));
OAI21X1 g21354(.A0 (n_252), .A1 (g18), .B0 (n_458), .Y (n_340));
OAI21X1 g21599(.A0 (n_258), .A1 (g_9514), .B0 (n_232), .Y (n_377));
AOI22X1 g21601(.A0 (n_803), .A1 (n_335), .B0 (g1275), .B1 (n_338), .Y(n_339));
AOI22X1 g21603(.A0 (n_803), .A1 (n_333), .B0 (n_335), .B1 (n_338), .Y(n_337));
AOI22X1 g21605(.A0 (n_803), .A1 (g1245), .B0 (n_333), .B1 (n_338), .Y(n_334));
AOI22X1 g21607(.A0 (n_803), .A1 (n_330), .B0 (g1245), .B1 (n_338), .Y(n_332));
AOI22X1 g21609(.A0 (n_803), .A1 (n_328), .B0 (n_330), .B1 (n_338), .Y(n_331));
DFFSRX1 g1110_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_271), .Q (g1110), .QN ());
AOI22X1 g21611(.A0 (n_803), .A1 (n_326), .B0 (n_328), .B1 (n_338), .Y(n_329));
AOI22X1 g21613(.A0 (n_803), .A1 (n_324), .B0 (n_326), .B1 (n_338), .Y(n_327));
AOI22X1 g21615(.A0 (n_803), .A1 (n_311), .B0 (n_324), .B1 (n_338), .Y(n_325));
AOI22X1 g21617(.A0 (n_803), .A1 (n_131), .B0 (n_321), .B1 (n_338), .Y(n_323));
AOI22X1 g21619(.A0 (n_803), .A1 (n_321), .B0 (n_319), .B1 (n_338), .Y(n_322));
AOI22X1 g21621(.A0 (n_803), .A1 (n_319), .B0 (n_317), .B1 (n_338), .Y(n_320));
AOI22X1 g21623(.A0 (n_803), .A1 (n_317), .B0 (n_314), .B1 (n_338), .Y(n_318));
OAI21X1 g21451(.A0 (n_251), .A1 (g18), .B0 (n_431), .Y (n_316));
AOI22X1 g21625(.A0 (n_803), .A1 (n_314), .B0 (n_312), .B1 (n_338), .Y(n_315));
AOI22X1 g21627(.A0 (n_803), .A1 (n_312), .B0 (n_311), .B1 (n_338), .Y(n_313));
DFFSRX1 g1371_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_276), .Q (), .QN (g1371));
DFFSRX1 g1383_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_268), .Q (g1383), .QN ());
DFFSRX1 g213_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_264), .Q (g_8484), .QN ());
DFFSRX1 g1377_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_261), .Q (), .QN (g1377));
DFFSRX1 g219_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_277), .Q (g_10714), .QN ());
DFFSRX1 g231_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_265), .Q (g_10572), .QN ());
DFFSRX1 g1107_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_273), .Q (g1107), .QN ());
DFFSRX1 g1101_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_270), .Q (n_112), .QN ());
DFFSRX1 g1104_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_274), .Q (g1104), .QN ());
DFFSRX1 g243_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_266), .Q (), .QN (g_10087));
NAND3X1 g21646(.A (n_295), .B (n_13), .C (g4173), .Y (n_310));
OAI21X1 g21377(.A0 (n_253), .A1 (g18), .B0 (n_354), .Y (n_309));
OAI21X1 g21488(.A0 (n_254), .A1 (g18), .B0 (n_426), .Y (n_307));
NAND3X1 g21735(.A (g741), .B (n_232), .C (g742), .Y (n_306));
NAND3X1 g21745(.A (g743), .B (g744), .C (n_232), .Y (n_305));
XOR2X1 g21516(.A (g4178), .B (n_246), .Y (n_304));
XOR2X1 g21526(.A (n_127), .B (n_286), .Y (n_303));
NAND2X1 g21533(.A (n_129), .B (n_300), .Y (n_302));
NAND2X1 g21534(.A (n_189), .B (n_300), .Y (n_301));
NAND2X1 g21535(.A (n_193), .B (n_300), .Y (n_299));
DFFSRX1 g1362_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_278), .Q (), .QN (g1362));
DFFSRX1 g1386_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_260), .Q (g1386), .QN ());
DFFSRX1 g1380_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_249), .Q (g1380), .QN ());
DFFSRX1 g237_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_238), .Q (), .QN (g_10859));
NOR2X1 g21641(.A (n_269), .B (g4173), .Y (n_348));
NAND2X1 g21638(.A (n_803), .B (g1275), .Y (n_297));
OAI21X1 g21393(.A0 (n_228), .A1 (g18), .B0 (n_438), .Y (n_288));
NAND2X1 g21530(.A (n_286), .B (n_128), .Y (n_287));
NAND2X1 g21531(.A (n_286), .B (n_188), .Y (n_285));
NAND2X1 g21532(.A (n_286), .B (g382), .Y (n_284));
NAND2X1 g21537(.A (n_800), .B (n_262), .Y (n_385));
OAI21X1 g21538(.A0 (n_226), .A1 (g18), .B0 (n_434), .Y (n_282));
OAI21X1 g21417(.A0 (n_227), .A1 (g18), .B0 (n_441), .Y (n_281));
OAI21X1 g21564(.A0 (n_595), .A1 (g1231), .B0 (n_262), .Y (n_280));
DFFSRX1 g1365_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_244), .Q (), .QN (g1365));
AOI21X1 g21589(.A0 (n_221), .A1 (n_46), .B0 (n_96), .Y (n_279));
NOR2X1 g21640(.A (g_10087), .B (n_275), .Y (n_278));
DFFSRX1 g1400_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_203), .Q (), .QN (g1400));
NOR2X1 g21444(.A (g1371), .B (n_275), .Y (n_277));
DFFSRX1 g1145_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_217), .Q (g1145), .QN ());
DFFSRX1 g1157_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_220), .Q (g1157), .QN ());
DFFSRX1 g1639_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_230), .Q (), .QN (g1639));
DFFSRX1 g1512_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_229), .Q (), .QN (g1512));
DFFSRX1 g186_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_233), .Q (g_10698), .QN ());
DFFSRX1 g207_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_222), .Q (g_10548), .QN ());
DFFSRX1 g1149_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_214), .Q (g1149), .QN ());
NOR2X1 g21455(.A (n_10), .B (n_275), .Y (n_276));
DFFSRX1 g1141_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_212), .Q (g1141), .QN ());
DFFSRX1 g248_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_210), .Q (g_9187), .QN ());
DFFSRX1 g1166_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_213), .Q (g1166), .QN ());
DFFSRX1 g1389_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_218), .Q (g1389), .QN ());
DFFSRX1 g1397_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_208), .Q (g1397), .QN ());
DFFSRX1 g1163_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_199), .Q (g1163), .QN ());
DFFSRX1 g197_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_219), .Q (g_2705), .QN ());
DFFSRX1 g1121_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_204), .Q (g1121), .QN ());
DFFSRX1 g1129_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_205), .Q (g1129), .QN ());
DFFSRX1 g1137_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_207), .Q (g1137), .QN ());
DFFSRX1 g113_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_257), .Q (), .QN (gbuf6));
AND2X1 g21656(.A (n_272), .B (g1104), .Y (n_274));
AND2X1 g21658(.A (n_272), .B (g1107), .Y (n_273));
AND2X1 g21659(.A (n_272), .B (g1110), .Y (n_271));
AND2X1 g21660(.A (n_272), .B (n_112), .Y (n_270));
DFFSRX1 g1125_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_200), .Q (g1125), .QN ());
INVX1 g21669(.A (n_269), .Y (n_295));
NOR2X1 g21379(.A (n_22), .B (n_275), .Y (n_268));
NOR2X1 g21693(.A (g1400), .B (n_275), .Y (n_266));
DFFSRX1 g1113_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_201), .Q (g1113), .QN ());
NOR2X1 g21523(.A (g1365), .B (n_275), .Y (n_265));
DFFSRX1 g192_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_211), .Q (g_7720), .QN ());
DFFSRX1 g1153_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_196), .Q (g1153), .QN ());
NOR2X1 g21413(.A (g1377), .B (n_275), .Y (n_264));
INVX1 g21547(.A (n_286), .Y (n_300));
INVX1 g21551(.A (n_262), .Y (n_263));
DFFSRX1 g1117_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_198), .Q (g1117), .QN ());
DFFSRX1 g225_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_231), .Q (g_7025), .QN ());
DFFSRX1 g1160_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_202), .Q (g1160), .QN ());
DFFSRX1 g1368_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_223), .Q (g1368), .QN ());
DFFSRX1 g1374_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_215), .Q (g1374), .QN ());
DFFSRX1 g1133_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_209), .Q (g1133), .QN ());
NOR2X1 g21425(.A (n_15), .B (n_275), .Y (n_261));
NOR2X1 g21357(.A (n_20), .B (n_275), .Y (n_260));
NAND4X1 g21645(.A (n_145), .B (n_150), .C (n_34), .D (n_141), .Y(n_259));
INVX1 g21650(.A (n_257), .Y (n_258));
NAND2X1 g21670(.A (g590), .B (n_232), .Y (n_269));
XOR2X1 g21673(.A (g1141), .B (n_171), .Y (n_254));
XOR2X1 g21674(.A (g1125), .B (n_173), .Y (n_253));
XOR2X1 g21675(.A (g1121), .B (n_169), .Y (n_252));
XOR2X1 g21681(.A (g1137), .B (n_174), .Y (n_251));
NOR2X1 g21397(.A (n_12), .B (n_275), .Y (n_249));
OAI21X1 g21644(.A0 (n_151), .A1 (n_247), .B0 (n_187), .Y (n_248));
DFFSRX1 g1289_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_184), .Q (g1289), .QN ());
INVX1 g21541(.A (n_712), .Y (n_246));
NOR2X1 g21544(.A (g_10859), .B (n_275), .Y (n_244));
XOR2X1 g21546(.A (g4177), .B (n_194), .Y (n_243));
CLKBUFX1 g21548(.A (n_814), .Y (n_286));
INVX2 g21552(.A (n_661), .Y (n_262));
NOR2X1 g21591(.A (g1362), .B (n_275), .Y (n_238));
XOR2X1 g21628(.A (g4176), .B (n_154), .Y (n_234));
DFFSRX1 g883_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_162), .Q (g2986), .QN ());
AND2X1 g21370(.A (g1383), .B (n_232), .Y (n_233));
OR2X1 g21651(.A (n_176), .B (n_275), .Y (n_257));
AND2X1 g21470(.A (g1368), .B (n_232), .Y (n_231));
XOR2X1 g21672(.A (g1117), .B (n_144), .Y (n_230));
XOR2X1 g21676(.A (g1113), .B (n_137), .Y (n_229));
XOR2X1 g21677(.A (g1129), .B (n_139), .Y (n_228));
XOR2X1 g21678(.A (g1133), .B (n_133), .Y (n_227));
XOR2X1 g21679(.A (g1145), .B (n_134), .Y (n_226));
INVX1 g21686(.A (n_225), .Y (n_386));
CLKBUFX1 g21689(.A (n_800), .Y (n_338));
NOR2X1 g21691(.A (g1216), .B (n_275), .Y (n_272));
DFFSRX1 g1206_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_224), .Q (g3069), .QN ());
AND2X1 g21495(.A (g_10572), .B (n_232), .Y (n_223));
AND2X1 g21390(.A (g1380), .B (n_232), .Y (n_222));
NOR2X1 g21643(.A (n_177), .B (n_116), .Y (n_221));
AND2X1 g21791(.A (g1157), .B (n_232), .Y (n_220));
AND2X1 g21796(.A (g1374), .B (n_232), .Y (n_219));
AND2X1 g21799(.A (g_2705), .B (n_232), .Y (n_218));
AND2X1 g21800(.A (g1145), .B (n_232), .Y (n_217));
AND2X1 g21803(.A (g_10749), .B (n_232), .Y (n_215));
AND2X1 g21805(.A (g1149), .B (n_232), .Y (n_214));
AND2X1 g21810(.A (g1166), .B (n_232), .Y (n_213));
AND2X1 g21811(.A (g1141), .B (n_232), .Y (n_212));
AND2X1 g21812(.A (g1389), .B (n_232), .Y (n_211));
AND2X1 g21814(.A (g1397), .B (n_232), .Y (n_210));
AND2X1 g21815(.A (g1133), .B (n_232), .Y (n_209));
AND2X1 g21816(.A (g_7720), .B (n_232), .Y (n_208));
AND2X1 g21823(.A (g1137), .B (n_232), .Y (n_207));
AND2X1 g21824(.A (g1129), .B (n_232), .Y (n_205));
AND2X1 g21827(.A (g1121), .B (n_232), .Y (n_204));
AND2X1 g21828(.A (g_9187), .B (n_232), .Y (n_203));
AND2X1 g21829(.A (g1160), .B (n_232), .Y (n_202));
AND2X1 g21836(.A (g1113), .B (n_232), .Y (n_201));
AND2X1 g21841(.A (g1125), .B (n_232), .Y (n_200));
AND2X1 g21843(.A (g1163), .B (n_232), .Y (n_199));
AND2X1 g21844(.A (g1117), .B (n_232), .Y (n_198));
NAND4X1 g21414(.A (n_178), .B (n_69), .C (n_48), .D (n_78), .Y(n_197));
AND2X1 g21848(.A (g1153), .B (n_232), .Y (n_196));
XOR2X1 g21565(.A (g382), .B (n_832), .Y (n_193));
XOR2X1 g21647(.A (n_188), .B (n_826), .Y (n_189));
INVX1 g21653(.A (n_595), .Y (n_187));
DFFSRX1 g590_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g1713), .Q (), .QN (g590));
DFFSRX1 g1718_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g1713), .Q (g1718), .QN ());
OR2X1 g21687(.A (g1212), .B (n_275), .Y (n_225));
OR2X1 g21688(.A (g869), .B (n_275), .Y (n_397));
OR2X1 g21694(.A (g1212), .B (g1289), .Y (n_184));
NOR2X1 g21427(.A (n_123), .B (g1368), .Y (n_178));
NAND4X1 g21671(.A (n_118), .B (n_47), .C (n_51), .D (n_77), .Y(n_177));
AOI21X1 g21695(.A0 (g882), .A1 (g2986), .B0 (g881), .Y (n_176));
NAND2X1 g21637(.A (n_153), .B (g4176), .Y (n_194));
NAND2X1 g21740(.A (n_172), .B (n_168), .Y (n_174));
NAND2X1 g21741(.A (n_172), .B (n_170), .Y (n_173));
NAND2X1 g21743(.A (n_170), .B (n_136), .Y (n_171));
NAND2X1 g21747(.A (n_168), .B (n_143), .Y (n_169));
OAI21X1 g21749(.A0 (n_596), .A1 (n_165), .B0 (n_597), .Y (n_167));
INVX1 g21756(.A (n_130), .Y (n_162));
NOR2X1 g21581(.A (n_160), .B (n_159), .Y (n_161));
AND2X1 g21584(.A (n_160), .B (n_159), .Y (n_224));
INVX1 g21680(.A (n_153), .Y (n_154));
XOR2X1 g21696(.A (g4175), .B (n_117), .Y (n_152));
INVX1 g21698(.A (n_597), .Y (n_151));
DFFSRX1 g869_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(gbuf5), .Q (g869), .QN ());
DFFSRX1 g1212_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(gbuf13), .Q (g1212), .QN ());
DFFSRX1 g1216_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(gbuf12), .Q (g1216), .QN ());
DFFSRX1 g1713_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g1710), .Q (g1713), .QN ());
NOR2X1 g21728(.A (n_149), .B (g1245), .Y (n_150));
OR2X1 g21729(.A (g1275), .B (n_146), .Y (n_148));
AND2X1 g21736(.A (n_92), .B (n_83), .Y (n_145));
AND2X1 g21737(.A (n_135), .B (n_143), .Y (n_144));
NOR2X1 g21742(.A (n_90), .B (n_91), .Y (n_141));
NAND2X1 g21746(.A (n_138), .B (n_143), .Y (n_140));
NAND2X1 g21750(.A (n_172), .B (n_138), .Y (n_139));
AND2X1 g21751(.A (n_136), .B (n_135), .Y (n_137));
NAND2X1 g21752(.A (n_136), .B (n_138), .Y (n_134));
NAND2X1 g21753(.A (n_172), .B (n_135), .Y (n_133));
XOR2X1 g21755(.A (n_59), .B (n_131), .Y (n_132));
NAND4X1 g21757(.A (n_26), .B (n_1), .C (n_32), .D (n_55), .Y (n_130));
XOR2X1 g21758(.A (n_128), .B (n_127), .Y (n_129));
DFFSRX1 g431_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_98), .Q (g431), .QN ());
NAND4X1 g21438(.A (n_61), .B (g1362), .C (g_10087), .D (g_10859), .Y(n_123));
DFFSRX1 g444_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_58), .Q (g_1301), .QN ());
DFFSRX1 g386_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_122), .Q (g_1328), .QN ());
DFFSRX1 g448_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_36), .Q (g_1298), .QN ());
DFFSRX1 g440_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_39), .Q (g_1304), .QN ());
DFFSRX1 g396_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_735), .Q (g_1334), .QN ());
DFFSRX1 g406_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_944), .Q (g_1340), .QN ());
DFFSRX1 g435_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_53), .Q (g_1307), .QN ());
AND2X1 g21655(.A (n_934), .B (n_119), .Y (n_160));
NOR2X1 g21657(.A (n_934), .B (n_119), .Y (n_120));
DFFSRX1 g391_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_737), .Q (g_1331), .QN ());
NOR2X1 g21731(.A (n_79), .B (g1160), .Y (n_118));
NOR2X1 g21732(.A (n_117), .B (n_25), .Y (n_153));
NAND2X1 g21748(.A (n_50), .B (n_49), .Y (n_116));
OR2X1 g21792(.A (n_311), .B (n_324), .Y (n_115));
NOR2X1 g21802(.A (n_112), .B (g1104), .Y (n_170));
AND2X1 g21821(.A (n_112), .B (g1104), .Y (n_168));
DFFSRX1 g452_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_849), .Q (g_1295), .QN ());
DFFSRX1 g421_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_818), .Q (g_1292), .QN ());
DFFSRX1 g401_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_913), .Q (n_945), .QN ());
OR2X1 g21789(.A (g_10749), .B (n_81), .Y (n_99));
OR2X1 g21639(.A (g_10087), .B (n_81), .Y (n_422));
DFFSRX1 g114_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_24), .Q (g_9514), .QN ());
INVX1 g21876(.A (n_925), .Y (n_98));
DFFSRX1 g416_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_892), .Q (g_1346), .QN ());
XOR2X1 g21759(.A (g1149), .B (g1153), .Y (n_96));
DFFSRX1 g876_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g3007), .Q (g876), .QN ());
DFFSRX1 g1710_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(1'b1), .Q (g1710), .QN ());
DFFSRX1 g1360_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(1'b1), .Q (gbuf12), .QN ());
DFFSRX1 g1217_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(1'b1), .Q (gbuf13), .QN ());
DFFSRX1 g875_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(1'b1), .Q (gbuf5), .QN ());
DFFSRX1 g882_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g2986), .Q (), .QN (g882));
NAND2X1 g21809(.A (n_37), .B (n_80), .Y (n_146));
NOR2X1 g21785(.A (n_95), .B (g1110), .Y (n_172));
AND2X1 g21786(.A (n_95), .B (g1110), .Y (n_136));
NOR2X1 g21787(.A (n_94), .B (g1104), .Y (n_138));
AND2X1 g21788(.A (n_94), .B (g1104), .Y (n_135));
DFFSRX1 g32_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_16), .Q (), .QN (g11163));
NAND2X1 g21790(.A (n_6), .B (g3007), .Y (n_93));
AND2X1 g21797(.A (n_42), .B (n_30), .Y (n_92));
NAND2X1 g21804(.A (n_59), .B (n_27), .Y (n_91));
NAND2X1 g21808(.A (n_62), .B (n_76), .Y (n_90));
NAND2X1 g21818(.A (n_70), .B (n_45), .Y (n_149));
NAND2X1 g21830(.A (g_9187), .B (g18), .Y (n_429));
DFFSRX1 g1361_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(g3069), .Q (), .QN (g1361));
AND2X1 g21847(.A (n_29), .B (n_44), .Y (n_83));
OR2X1 g21545(.A (g_10859), .B (n_81), .Y (n_434));
DFFSRX1 g411_reg(.RN (n_533), .SN (1'b1), .CK (blif_clk_net), .D(n_854), .Q (g_1343), .QN ());
INVX4 g21948(.A (n_275), .Y (n_232));
NAND2X1 g21458(.A (g_7025), .B (g18), .Y (n_431));
NAND2X1 g21426(.A (g_10714), .B (g18), .Y (n_441));
INVX2 g21953(.A (n_40), .Y (n_122));
INVX1 g21963(.A (n_80), .Y (n_333));
OR2X1 g21839(.A (g1153), .B (g1145), .Y (n_79));
NOR2X1 g21838(.A (g_10749), .B (g_2705), .Y (n_78));
NOR2X1 g21833(.A (g1166), .B (g1113), .Y (n_77));
NAND2X1 g21358(.A (g_10698), .B (g18), .Y (n_458));
INVX1 g21898(.A (n_76), .Y (n_319));
INVX1 g21973(.A (n_641), .Y (n_127));
INVX1 g21929(.A (n_916), .Y (n_188));
INVX1 g21853(.A (n_70), .Y (n_328));
NOR2X1 g21461(.A (g_7025), .B (g_10572), .Y (n_69));
NAND2X1 g21398(.A (g_8484), .B (g18), .Y (n_438));
INVX1 g21886(.A (n_62), .Y (n_317));
AND2X1 g21445(.A (g1371), .B (g1365), .Y (n_61));
INVX1 g21879(.A (n_598), .Y (n_247));
NOR2X1 g21813(.A (g1107), .B (g1110), .Y (n_143));
NAND2X1 g21380(.A (g_10548), .B (g18), .Y (n_354));
INVX1 g21865(.A (n_59), .Y (n_321));
NAND2X1 g21498(.A (g_10572), .B (g18), .Y (n_426));
INVX1 g21927(.A (n_697), .Y (n_58));
INVX1 g21912(.A (n_52), .Y (n_53));
NOR2X1 g21801(.A (g1163), .B (g1149), .Y (n_51));
NOR2X1 g21806(.A (g1129), .B (g1133), .Y (n_50));
NOR2X1 g21842(.A (g1137), .B (g1141), .Y (n_49));
NOR2X1 g21807(.A (g1389), .B (g_7720), .Y (n_48));
NOR2X1 g21817(.A (g1121), .B (g1157), .Y (n_47));
NAND2X1 g21825(.A (g4174), .B (g4173), .Y (n_117));
NAND2X1 g21831(.A (g_7720), .B (g18), .Y (n_345));
NOR2X1 g21837(.A (g1125), .B (g1117), .Y (n_46));
INVX1 g21849(.A (n_45), .Y (n_326));
INVX1 g21857(.A (n_44), .Y (n_311));
INVX1 g21868(.A (n_642), .Y (n_128));
INVX1 g21881(.A (n_42), .Y (n_312));
INVX1 g21905(.A (n_38), .Y (n_39));
INVX1 g21969(.A (n_37), .Y (n_335));
INVX1 g21907(.A (n_700), .Y (n_36));
INVX1 g21959(.A (n_600), .Y (n_165));
INVX1 g21961(.A (n_30), .Y (n_314));
INVX1 g21965(.A (n_29), .Y (n_131));
INVX1 g21887(.A (g1296), .Y (n_62));
INVX1 g21972(.A (g1351), .Y (n_159));
INVX1 g21893(.A (blif_reset_net), .Y (n_533));
INVX1 g21917(.A (g986), .Y (n_342));
INVX1 g21871(.A (g936), .Y (n_55));
INVX1 g21976(.A (g_1334), .Y (n_28));
INVX1 g21955(.A (g_1325), .Y (n_40));
CLKBUFX1 g21862(.A (g1265), .Y (n_324));
INVX1 g21863(.A (g1265), .Y (n_27));
INVX1 g21851(.A (g928), .Y (n_26));
INVX1 g21904(.A (g1107), .Y (n_95));
INVX1 g21882(.A (g1304), .Y (n_42));
INVX1 g21858(.A (g1270), .Y (n_44));
INVX1 g21966(.A (g1280), .Y (n_29));
INVX1 g21958(.A (g940), .Y (n_32));
INVX1 g21875(.A (g4175), .Y (n_25));
INVX1 g21899(.A (g1292), .Y (n_76));
INVX1 g21911(.A (gbuf6), .Y (n_24));
INVX1 g21384(.A (g_10548), .Y (n_22));
INVX1 g21902(.A (g981), .Y (n_235));
INVX1 g21885(.A (g1346), .Y (n_119));
INVX1 g21964(.A (g1240), .Y (n_80));
INVX1 g21856(.A (n_112), .Y (n_94));
INVX1 g21970(.A (g1235), .Y (n_37));
INVX1 g21362(.A (g_10698), .Y (n_20));
INVX1 g21901(.A (g_1340), .Y (n_19));
INVX1 g21890(.A (g976), .Y (n_124));
INVX1 g21906(.A (g_1301), .Y (n_38));
INVX1 g21874(.A (g1341), .Y (n_17));
INVX1 g21861(.A (g11163), .Y (n_16));
INVX1 g21431(.A (g_10714), .Y (n_15));
INVX1 g21854(.A (g1255), .Y (n_70));
INVX1 g21883(.A (g4174), .Y (n_13));
INVX1 g21401(.A (g_8484), .Y (n_12));
INVX1 g21952(.A (n_330), .Y (n_34));
INVX1 g21464(.A (g_7025), .Y (n_10));
INVX1 g21852(.A (g4177), .Y (n_9));
INVX1 g21866(.A (g1284), .Y (n_59));
INVX1 g21968(.A (g876), .Y (n_6));
INVX1 g21910(.A (g_1343), .Y (n_5));
INVX1 g21850(.A (g1260), .Y (n_45));
INVX1 g21962(.A (g1300), .Y (n_30));
INVX1 g21913(.A (g_1304), .Y (n_52));
INVX1 g21864(.A (g932), .Y (n_1));
INVX1 g21921(.A (g18), .Y (n_81));
INVX1 g22142(.A (n_543), .Y (n_544));
INVX2 g22143(.A (n_763), .Y (n_543));
INVX1 g22148(.A (n_722), .Y (n_551));
INVX1 g22157(.A (n_797), .Y (n_576));
NAND3X1 g22159(.A (n_676), .B (n_841), .C (n_588), .Y (n_589));
INVX1 g43(.A (n_587), .Y (n_588));
NAND2X1 g44(.A (n_773), .B (n_586), .Y (n_587));
NOR2X1 g46(.A (n_584), .B (n_585), .Y (n_586));
NOR2X1 g58(.A (g971), .B (n_124), .Y (n_584));
AND2X1 g49(.A (n_124), .B (g971), .Y (n_585));
INVX1 g22(.A (n_593), .Y (n_594));
NAND3X1 g15(.A (g1223), .B (g1218), .C (g1227), .Y (n_593));
CLKBUFX1 g1(.A (n_594), .Y (n_595));
NAND2X1 g16(.A (g1223), .B (n_596), .Y (n_597));
CLKBUFX1 g21(.A (g1218), .Y (n_596));
INVX1 g17(.A (g1227), .Y (n_598));
INVX1 g22160(.A (g1223), .Y (n_600));
AND2X1 g22163(.A (n_585), .B (n_235), .Y (n_606));
OAI21X1 g40(.A0 (n_585), .A1 (n_235), .B0 (n_773), .Y (n_608));
INVX1 g22176(.A (g369), .Y (n_641));
INVX1 g14(.A (g374), .Y (n_642));
OAI21X1 g22187(.A0 (n_259), .A1 (n_148), .B0 (n_132), .Y (n_660));
AND2X1 g22188(.A (n_594), .B (g1231), .Y (n_661));
OR4X1 g22190(.A (g1275), .B (n_330), .C (n_146), .D (n_149), .Y(n_664));
OR2X1 g22192(.A (g1245), .B (n_115), .Y (n_665));
NOR2X1 g22196(.A (g971), .B (n_835), .Y (n_671));
OR2X1 g22200(.A (n_754), .B (n_576), .Y (n_676));
AOI21X1 g22203(.A0 (n_679), .A1 (g590), .B0 (n_680), .Y (n_681));
NAND3X1 g22204(.A (g4181), .B (g4180), .C (n_711), .Y (n_679));
NOR2X1 g19(.A (g590), .B (n_679), .Y (n_680));
NAND2X1 g22205(.A (g4180), .B (n_711), .Y (n_682));
NAND2X1 g22210(.A (n_28), .B (n_942), .Y (n_686));
NOR2X1 g22212(.A (g_1325), .B (g_1331), .Y (n_689));
INVX1 g22213(.A (g_1328), .Y (n_690));
NOR2X1 g22217(.A (g431), .B (g_1292), .Y (n_694));
NOR2X1 g22218(.A (g_1295), .B (g_1298), .Y (n_695));
INVX1 g22219(.A (g_1298), .Y (n_697));
INVX1 g22220(.A (g_1295), .Y (n_700));
NOR2X1 g22228(.A (n_194), .B (n_710), .Y (n_711));
NAND3X1 g22229(.A (g4177), .B (g4178), .C (g4179), .Y (n_710));
NAND2X1 g22231(.A (n_712), .B (g4178), .Y (n_713));
NOR2X1 g22232(.A (n_194), .B (n_9), .Y (n_712));
NAND2X1 g37(.A (n_850), .B (n_893), .Y (n_718));
INVX1 g22237(.A (n_747), .Y (n_722));
NAND2X1 g27_dup(.A (n_815), .B (n_829), .Y (n_730));
AOI21X1 g50(.A0 (g324), .A1 (n_913), .B0 (n_739), .Y (n_740));
NAND2X1 g52(.A (n_736), .B (n_738), .Y (n_739));
NAND2X1 g54(.A (n_735), .B (g321), .Y (n_736));
CLKBUFX1 g22249(.A (g_1331), .Y (n_735));
NAND2X1 g53(.A (n_737), .B (g318), .Y (n_738));
CLKBUFX1 g2(.A (g_1328), .Y (n_737));
INVX1 g57(.A (n_485), .Y (n_741));
NOR2X1 g56(.A (n_479), .B (n_481), .Y (n_742));
AOI21X1 g22250(.A0 (g327), .A1 (n_944), .B0 (n_912), .Y (n_744));
NAND3X1 g22251(.A (n_750), .B (n_805), .C (n_798), .Y (n_754));
NAND2X1 g22252(.A (n_747), .B (n_749), .Y (n_750));
NAND2X1 g31(.A (n_815), .B (n_829), .Y (n_747));
INVX1 g22253(.A (n_748), .Y (n_749));
CLKBUFX1 g22254(.A (g305), .Y (n_748));
AND2X1 g30(.A (g305), .B (n_828), .Y (n_751));
NAND2X2 g10(.A (g374), .B (g369), .Y (n_756));
NAND2X1 g22258(.A (n_763), .B (n_764), .Y (n_765));
INVX2 g22259(.A (n_762), .Y (n_763));
NAND2X2 g22260(.A (n_809), .B (n_841), .Y (n_762));
NOR2X1 g22264(.A (n_606), .B (n_608), .Y (n_764));
AND2X1 g22272(.A (n_518), .B (n_232), .Y (n_773));
NOR2X1 g22288(.A (n_475), .B (n_823), .Y (n_792));
INVX1 g36(.A (n_718), .Y (n_793));
NOR2X1 g22289(.A (n_475), .B (n_806), .Y (n_797));
NOR2X1 g22290(.A (n_823), .B (n_718), .Y (n_798));
INVX2 g12(.A (n_802), .Y (n_803));
OR2X1 g13(.A (n_800), .B (n_275), .Y (n_802));
NOR2X1 g22291(.A (g1713), .B (n_799), .Y (n_800));
INVX1 g22292(.A (g1289), .Y (n_799));
INVX4 g22293(.A (g109), .Y (n_275));
NAND3X1 g22294(.A (n_804), .B (n_805), .C (n_808), .Y (n_809));
NAND2X1 g39(.A (n_730), .B (n_749), .Y (n_804));
NAND2X1 g41(.A (n_751), .B (n_815), .Y (n_805));
NOR2X1 g22295(.A (n_806), .B (n_807), .Y (n_808));
NAND4X1 g22296(.A (n_740), .B (n_742), .C (n_744), .D (n_741), .Y(n_806));
NAND2X1 g22297(.A (n_793), .B (n_792), .Y (n_807));
NAND2X2 g29(.A (n_900), .B (n_814), .Y (n_815));
INVX1 g33(.A (n_834), .Y (n_814));
CLKBUFX1 g22302(.A (g_1346), .Y (n_816));
CLKBUFX1 g22303(.A (n_816), .Y (n_818));
INVX1 g22304(.A (g_1346), .Y (n_819));
NAND2X2 g22305(.A (n_820), .B (n_853), .Y (n_823));
XOR2X1 g22306(.A (g309), .B (n_816), .Y (n_820));
CLKBUFX1 g22309(.A (n_828), .Y (n_829));
NAND2X1 g22310(.A (n_827), .B (g305), .Y (n_828));
NAND2X1 g15_dup(.A (n_915), .B (n_826), .Y (n_827));
INVX2 g22313(.A (n_756), .Y (n_826));
NOR2X1 g22315(.A (n_916), .B (n_756), .Y (n_832));
NAND2X2 g22317(.A (n_837), .B (n_839), .Y (n_840));
OAI21X1 g22318(.A0 (n_833), .A1 (n_835), .B0 (n_836), .Y (n_837));
NOR2X1 g22319(.A (n_754), .B (n_576), .Y (n_833));
CLKBUFX1 g22320(.A (n_834), .Y (n_835));
NAND2X1 g34(.A (n_915), .B (n_826), .Y (n_834));
AND2X1 g35(.A (n_773), .B (g971), .Y (n_836));
OAI21X1 g22321(.A0 (n_576), .A1 (n_754), .B0 (n_838), .Y (n_839));
AND2X1 g22322(.A (n_671), .B (n_773), .Y (n_838));
INVX1 g22323(.A (n_835), .Y (n_841));
NAND2X1 g22329(.A (n_38), .B (n_52), .Y (n_846));
XOR2X1 g22330(.A (g312), .B (n_849), .Y (n_850));
CLKBUFX3 g22331(.A (g_1292), .Y (n_849));
XOR2X1 g22333(.A (g330), .B (n_852), .Y (n_853));
CLKBUFX1 g22334(.A (g_1340), .Y (n_852));
CLKBUFX1 g11(.A (n_852), .Y (n_854));
OAI21X1 g22339(.A0 (n_859), .A1 (n_863), .B0 (n_864), .Y (n_865));
AND2X1 g24(.A (n_931), .B (n_891), .Y (n_859));
NAND2X1 g23(.A (n_861), .B (n_862), .Y (n_863));
INVX1 g25(.A (n_927), .Y (n_861));
INVX1 g22340(.A (g1336), .Y (n_862));
NAND3X1 g22341(.A (n_859), .B (n_861), .C (g1336), .Y (n_864));
NAND2X1 g47(.A (n_19), .B (n_924), .Y (n_869));
NAND2X1 g22344(.A (n_819), .B (n_5), .Y (n_870));
CLKBUFX1 g22358(.A (n_661), .Y (n_885));
NAND2X1 g22361(.A (n_918), .B (n_940), .Y (n_891));
XOR2X1 g22362(.A (g333), .B (n_892), .Y (n_893));
CLKBUFX2 g22363(.A (g_1343), .Y (n_892));
NAND2X2 g22365(.A (n_951), .B (n_926), .Y (n_900));
NOR2X1 g4(.A (g_1334), .B (g324), .Y (n_912));
CLKBUFX1 g22381(.A (g_1334), .Y (n_913));
AND2X1 g8(.A (g378), .B (g382), .Y (n_915));
INVX1 g9(.A (g378), .Y (n_916));
NOR2X1 g22385(.A (n_664), .B (n_665), .Y (n_918));
XOR2X1 g22388(.A (n_923), .B (n_925), .Y (n_926));
CLKBUFX1 g22389(.A (g431), .Y (n_923));
CLKBUFX3 g22390(.A (n_924), .Y (n_925));
INVX1 g22391(.A (g_1307), .Y (n_924));
NAND2X1 g22392(.A (n_933), .B (n_938), .Y (n_939));
NAND2X1 g51(.A (n_928), .B (n_932), .Y (n_933));
NOR2X1 g22393(.A (g1341), .B (n_927), .Y (n_928));
OR2X1 g22394(.A (n_275), .B (n_486), .Y (n_927));
NAND2X2 g22395(.A (n_929), .B (n_931), .Y (n_932));
NAND2X1 g22396(.A (n_941), .B (n_918), .Y (n_929));
INVX1 g59(.A (n_930), .Y (n_931));
NAND2X1 g60(.A (n_263), .B (n_800), .Y (n_930));
OR2X1 g22397(.A (n_936), .B (n_937), .Y (n_938));
OR2X1 g55(.A (n_934), .B (n_935), .Y (n_936));
NOR2X1 g22398(.A (g1336), .B (g1341), .Y (n_934));
NOR2X1 g61(.A (n_17), .B (n_862), .Y (n_935));
NAND3X1 g22399(.A (n_891), .B (n_931), .C (n_861), .Y (n_937));
NAND2X1 g22400(.A (n_660), .B (n_885), .Y (n_940));
NAND2X1 g22384_dup(.A (n_660), .B (n_885), .Y (n_941));
INVX1 g22401(.A (n_945), .Y (n_942));
CLKBUFX1 g22403(.A (n_945), .Y (n_944));
NAND3X1 g22404(.A (n_948), .B (n_949), .C (n_950), .Y (n_951));
NOR2X1 g22405(.A (n_946), .B (n_947), .Y (n_948));
NAND2X1 g22406(.A (n_690), .B (n_695), .Y (n_946));
NAND2X1 g38(.A (n_694), .B (n_689), .Y (n_947));
NOR2X1 g22407(.A (n_846), .B (n_686), .Y (n_949));
NOR2X1 g22408(.A (n_869), .B (n_870), .Y (n_950));
endmodule
