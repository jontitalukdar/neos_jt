module s38584(blif_clk_net, blif_reset_net, g35, g36, g6744,g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753,g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178,g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353,g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785,g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917,g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306,g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770,g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832,g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259,g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096,g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451,g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738,g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659,g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874,g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423,g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649,g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739,g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845,g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099,g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652,g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292,g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759,g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584,g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875,g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210,g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218,g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332,g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863,g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636,g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948,g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234,g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425,g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915,g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972);
input blif_clk_net, blif_reset_net, g35, g36, g6744, g6745, g6746,g6747, g6748, g6749, g6750, g6751, g6752, g6753;
output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178,g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353,g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785,g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917,g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306,g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770,g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832,g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259,g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096,g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451,g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738,g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659,g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874,g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423,g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649,g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739,g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845,g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099,g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652,g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292,g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759,g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584,g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875,g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210,g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218,g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332,g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863,g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636,g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948,g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234,g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425,g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915,g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972;
wire blif_clk_net, blif_reset_net, g35, g36, g6744, g6745, g6746,g6747, g6748, g6749, g6750, g6751, g6752, g6753;
wire g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178,g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353,g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785,g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917,g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306,g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770,g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832,g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259,g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096,g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451,g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738,g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659,g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874,g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423,g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649,g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739,g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845,g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099,g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652,g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292,g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759,g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584,g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875,g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210,g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218,g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332,g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863,g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636,g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948,g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234,g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425,g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915,g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972;
wire g55, g1171, g1178, g1183, g1189, g1199, g1221, g1236;
wire g1242, g1246, g1291, g1300, g1306, g1312, g1319, g1322;
wire g1333, g1339, g1345, g1351, g1361, g1367, g1373, g1379;
wire g1384, g1389, g1395, g1404, g1413, g1430, g1437, g1442;
wire g1448, g1454, g1467, g1472, g1478, g1484, g1489, g1521;
wire g1526, g1532, g1536, g1542, g1548, g1554, g1564, g1579;
wire g1585, g1589, g1592, g1600, g1604, g1608, g1612, g1616;
wire g1620, g1624, g1632, g1636, g1644, g1657, g1664, g1677;
wire g1682, g1687, g1691, g1696, g1700, g1706, g1710, g1714;
wire g1720, g1724, g1728, g1736, g1740, g1744, g1748, g1752;
wire g1756, g1760, g1768, g1772, g1779, g1792, g1798, g1811;
wire g1816, g1821, g1825, g1830, g1834, g1840, g1844, g1848;
wire g1854, g1858, g1862, g1870, g1874, g1878, g1882, g1886;
wire g1890, g1894, g1902, g1906, g1913, g1926, g1932, g1936;
wire g1945, g1950, g1955, g1959, g1964, g1968, g1974, g1978;
wire g1982, g1988, g1992, g1996, g2004, g2008, g2012, g2016;
wire g2020, g2024, g2028, g2036, g2040, g2047, g2060, g2066;
wire g2070, g2079, g2084, g2089, g2093, g2098, g2102, g2108;
wire g2112, g2116, g2122, g2126, g2130, g2138, g2145, g2153;
wire g2161, g2165, g2169, g2173, g2177, g2181, g2185, g2193;
wire g2197, g2204, g2217, g2223, g2227, g2236, g2241, g2246;
wire g2250, g2255, g2259, g2265, g2269, g2273, g2279, g2283;
wire g2287, g2295, g2299, g2303, g2307, g2311, g2315, g2319;
wire g2327, g2331, g2338, g2351, g2357, g2361, g2370, g2375;
wire g2380, g2384, g2389, g2393, g2399, g2403, g2407, g2413;
wire g2417, g2421, g2429, g2433, g2437, g2441, g2445, g2449;
wire g2453, g2461, g2465, g2472, g2485, g2491, g2504, g2509;
wire g2514, g2518, g2523, g2527, g2533, g2537, g2541, g2547;
wire g2551, g2555, g2563, g2567, g2571, g2575, g2579, g2583;
wire g2587, g2595, g2599, g2606, g2619, g2625, g2629, g2638;
wire g2643, g2648, g2652, g2657, g2661, g2667, g2671, g2675;
wire g2681, g2685, g2697, g2704, g2715, g2724, g2735, g2748;
wire g2756, g2759, g2763, g2767, g2771, g2775, g2779, g2783;
wire g2787, g2791, g2795, g2799, g2803, g2807, g2811, g2815;
wire g2819, g2823, g2827, g2844, g2848, g2852, g2856, g2860;
wire g2864, g2868, g2873, g2878, g2882, g2886, g2890, g2894;
wire g2898, g2902, g2907, g2912, g2917, g2922, g2927, g2932;
wire g2936, g2941, g2946, g2950, g2955, g2960, g2965, g2970;
wire g2975, g2980, g2984, g2988, g2994, g2999, g3003, g3050;
wire g3100, g3106, g3111, g3115, g3119, g3125, g3129, g3133;
wire g3139, g3143, g3147, g3155, g3161, g3171, g3179, g3187;
wire g3191, g3195, g3199, g3203, g3207, g3211, g3215, g3219;
wire g3223, g3227, g3231, g3235, g3239, g3243, g3247, g3251;
wire g3255, g3259, g3263, g3288, g3329, g3333, g3338, g3343;
wire g3347, g3401, g3451, g3457, g3462, g3466, g3470, g3476;
wire g3480, g3484, g3490, g3494, g3498, g3506, g3512, g3522;
wire g3530, g3538, g3542, g3546, g3550, g3554, g3558, g3562;
wire g3566, g3570, g3574, g3578, g3582, g3586, g3590, g3594;
wire g3598, g3602, g3606, g3610, g3614, g3639, g3680, g3684;
wire g3689, g3694, g3698, g3752, g3802, g3808, g3813, g3817;
wire g3821, g3827, g3831, g3835, g3841, g3845, g3849, g3857;
wire g3863, g3873, g3881, g3889, g3893, g3897, g3901, g3905;
wire g3909, g3913, g3917, g3921, g3925, g3929, g3933, g3937;
wire g3941, g3945, g3949, g3953, g3957, g3961, g3965, g3990;
wire g4031, g4035, g4040, g4045, g4049, g4054, g4057, g4064;
wire g4072, g4076, g4082, g4087, g4093, g4098, g4104, g4108;
wire g4112, g4116, g4119, g4122, g4141, g4145, g4146, g4153;
wire g4157, g4164, g4172, g4176, g4235, g4239, g4242, g4245;
wire g4249, g4253, g4258, g4264, g4269, g4273, g4281, g4284;
wire g4291, g4297, g4300, g4308, g4311, g4332, g4349, g4366;
wire g4369, g4372, g4375, g4382, g4388, g4392, g4401, g4405;
wire g4411, g4417, g4420, g4423, g4427, g4430, g4434, g4438;
wire g4443, g4452, g4455, g4456, g4459, g4462, g4467, g4473;
wire g4474, g4477, g4480, g4483, g4486, g4489, g4492, g4495;
wire g4498, g4501, g4504, g4512, g4515, g4519, g4521, g4527;
wire g4531, g4534, g4540, g4543, g4546, g4549, g4552, g4555;
wire g4558, g4561, g4564, g4567, g4570, g4572, g4575, g4578;
wire g4581, g4584, g4593, g4601, g4608, g4616, g4621, g4628;
wire g4633, g4653, g4659, g4664, g4669, g4688, g4698, g4704;
wire g4709, g4717, g4722, g4727, g4732, g4737, g4743, g4749;
wire g4754, g4760, g4765, g4771, g4776, g4785, g4793, g4821;
wire g4826, g4831, g4843, g4849, g4854, g4878, g4888, g4894;
wire g4899, g4907, g4912, g4917, g4922, g4927, g4933, g4939;
wire g4944, g4950, g4955, g4961, g4966, g4983, g4991, g5011;
wire g5016, g5029, g5033, g5037, g5041, g5046, g5052, g5057;
wire g5069, g5073, g5077, g5080, g5084, g5092, g5097, g5109;
wire g5112, g5120, g5124, g5128, g5134, g5138, g5142, g5148;
wire g5152, g5156, g5164, g5170, g5180, g5188, g5196, g5200;
wire g5204, g5208, g5212, g5216, g5220, g5224, g5228, g5232;
wire g5236, g5240, g5244, g5248, g5252, g5256, g5260, g5264;
wire g5268, g5272, g5297, g5339, g5343, g5348, g5352, g5406;
wire g5456, g5467, g5471, g5475, g5481, g5485, g5489, g5495;
wire g5499, g5503, g5511, g5517, g5527, g5535, g5543, g5547;
wire g5551, g5555, g5559, g5563, g5567, g5571, g5575, g5579;
wire g5583, g5587, g5591, g5595, g5599, g5603, g5607, g5611;
wire g5615, g5619, g5644, g5685, g5689, g5694, g5698, g5752;
wire g5802, g5813, g5817, g5821, g5827, g5831, g5835, g5841;
wire g5845, g5849, g5857, g5863, g5873, g5881, g5889, g5893;
wire g5897, g5901, g5905, g5909, g5913, g5917, g5921, g5925;
wire g5929, g5933, g5937, g5941, g5945, g5949, g5953, g5957;
wire g5961, g5965, g5990, g6031, g6035, g6040, g6044, g6098;
wire g6148, g6159, g6163, g6167, g6173, g6177, g6181, g6187;
wire g6191, g6195, g6203, g6209, g6219, g6227, g6235, g6239;
wire g6243, g6247, g6251, g6255, g6259, g6263, g6267, g6271;
wire g6275, g6279, g6283, g6287, g6291, g6295, g6299, g6303;
wire g6307, g6311, g6336, g6377, g6381, g6386, g6390, g6395;
wire g6444, g6494, g6505, g6509, g6513, g6519, g6523, g6527;
wire g6533, g6537, g6541, g6549, g6555, g6565, g6573, g6581;
wire g6585, g6589, g6593, g6597, g6601, g6605, g6609, g6613;
wire g6617, g6621, g6625, g6629, g6633, g6637, g6641, g6645;
wire g6649, g6653, g6657, g6723, g6732, g6736, g6741, g34026;
wire g34027, g34028, g34034, g34035, g34036, g_3381, g_3861, g_3974;
wire g_4050, g_4409, g_4449, g_5029, g_5156, g_5313, g_5342, g_5450;
wire g_5508, g_6131, g_6165, g_6192, g_6283, g_6579, g_6701, g_7062;
wire g_7220, g_7563, g_8657, g_8864, g_8896, g_9174, g_9176, g_9298;
wire g_9338, g_9584, g_10092, g_10233, g_10278, g_10556, g_10715,g_10903;
wire g_11037, g_11293, g_11413, g_12275, g_12276, g_12433, g_12465,g_12791;
wire g_12922, g_13091, g_13255, g_13278, g_13758, g_13838, g_13871,g_13901;
wire g_14265, g_14342, g_14535, g_14587, g_14843, g_14965, g_15016,g_15127;
wire g_15287, g_15380, g_15381, g_15691, g_15740, g_15758, g_15801,g_15838;
wire g_15879, g_16063, g_16296, g_16311, g_16404, g_16456, g_16464,g_16475;
wire g_16571, g_16677, g_16769, g_16792, g_16958, g_16983, g_17065,g_17086;
wire g_17426, g_17653, g_17934, g_18015, g_18112, g_18200, g_18220,g_18238;
wire g_18308, g_18330, g_18488, g_18590, g_18635, g_18739, g_18793,g_18795;
wire g_18869, g_18902, g_18980, g_18996, g_19113, g_19136, g_19172,g_19187;
wire g_19233, g_19241, g_19289, g_19304, g_19414, g_19459, g_19492,g_19515;
wire g_19659, g_19789, g_19911, g_19913, g_20073, g_20159, g_20208,g_20244;
wire g_20268, g_20563, g_20614, g_20837, g_20839, g_20909, g_20951,g_20952;
wire g_21318, g_21447, g_21576, g_21651, g_21720, g_21778, g_21792,g_21799;
wire g_21806, g_21813, g_22021, g_22034, g_22038, g_22070, g_22236,g_22306;
wire g_22328, g_22349, g_22371, g_22379, g_22464, g_22552, g_22600,g_22605;
wire g_22639, gbuf1, gbuf3, n_0, n_1, n_2, n_5, n_11;
wire n_12, n_13, n_16, n_17, n_19, n_20, n_21, n_22;
wire n_23, n_26, n_27, n_28, n_29, n_30, n_32, n_35;
wire n_38, n_39, n_40, n_43, n_46, n_50, n_52, n_54;
wire n_57, n_59, n_60, n_64, n_65, n_67, n_69, n_70;
wire n_74, n_75, n_79, n_83, n_85, n_86, n_87, n_89;
wire n_92, n_93, n_94, n_95, n_96, n_98, n_101, n_103;
wire n_105, n_107, n_110, n_117, n_118, n_125, n_126, n_127;
wire n_128, n_129, n_134, n_136, n_143, n_144, n_150, n_151;
wire n_153, n_157, n_158, n_162, n_165, n_168, n_169, n_172;
wire n_187, n_188, n_191, n_194, n_196, n_202, n_204, n_205;
wire n_209, n_213, n_215, n_218, n_220, n_221, n_223, n_224;
wire n_227, n_234, n_235, n_238, n_240, n_241, n_242, n_243;
wire n_245, n_247, n_248, n_251, n_259, n_261, n_262, n_263;
wire n_268, n_269, n_271, n_273, n_276, n_278, n_281, n_282;
wire n_284, n_286, n_287, n_290, n_291, n_294, n_295, n_297;
wire n_298, n_302, n_303, n_307, n_308, n_309, n_311, n_316;
wire n_317, n_322, n_323, n_325, n_326, n_327, n_328, n_330;
wire n_332, n_334, n_335, n_336, n_338, n_339, n_340, n_342;
wire n_343, n_344, n_347, n_351, n_353, n_356, n_360, n_362;
wire n_364, n_365, n_367, n_368, n_370, n_371, n_374, n_376;
wire n_377, n_379, n_380, n_382, n_383, n_386, n_388, n_389;
wire n_392, n_397, n_399, n_401, n_404, n_406, n_408, n_409;
wire n_411, n_412, n_413, n_415, n_416, n_417, n_418, n_423;
wire n_424, n_425, n_428, n_429, n_433, n_436, n_437, n_441;
wire n_442, n_444, n_446, n_447, n_448, n_450, n_453, n_455;
wire n_456, n_458, n_459, n_460, n_461, n_463, n_464, n_465;
wire n_469, n_470, n_471, n_474, n_477, n_479, n_482, n_486;
wire n_487, n_488, n_490, n_491, n_493, n_496, n_503, n_504;
wire n_511, n_512, n_515, n_518, n_519, n_521, n_522, n_523;
wire n_524, n_527, n_538, n_540, n_546, n_549, n_551, n_552;
wire n_553, n_556, n_557, n_558, n_561, n_562, n_563, n_564;
wire n_565, n_566, n_568, n_571, n_572, n_575, n_578, n_579;
wire n_580, n_581, n_584, n_585, n_587, n_588, n_589, n_590;
wire n_591, n_592, n_594, n_595, n_596, n_597, n_598, n_599;
wire n_600, n_603, n_607, n_608, n_609, n_610, n_611, n_612;
wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_623;
wire n_624, n_626, n_627, n_628, n_629, n_635, n_636, n_637;
wire n_638, n_639, n_640, n_643, n_644, n_647, n_648, n_649;
wire n_650, n_652, n_653, n_659, n_660, n_661, n_662, n_663;
wire n_664, n_667, n_669, n_670, n_673, n_674, n_675, n_676;
wire n_677, n_678, n_680, n_684, n_685, n_686, n_688, n_690;
wire n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
wire n_702, n_704, n_705, n_707, n_708, n_709, n_714, n_715;
wire n_716, n_717, n_718, n_719, n_720, n_722, n_723, n_724;
wire n_730, n_739, n_740, n_741, n_744, n_745, n_746, n_747;
wire n_748, n_765, n_769, n_771, n_772, n_775, n_776, n_777;
wire n_778, n_779, n_780, n_782, n_783, n_784, n_786, n_789;
wire n_790, n_791, n_793, n_794, n_795, n_797, n_798, n_799;
wire n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807;
wire n_808, n_810, n_812, n_814, n_816, n_817, n_818, n_819;
wire n_820, n_821, n_822, n_823, n_824, n_826, n_827, n_828;
wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
wire n_845, n_846, n_847, n_848, n_849, n_851, n_852, n_854;
wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
wire n_863, n_864, n_866, n_867, n_868, n_871, n_872, n_876;
wire n_877, n_878, n_880, n_881, n_882, n_883, n_884, n_885;
wire n_886, n_887, n_888, n_890, n_891, n_893, n_894, n_895;
wire n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903;
wire n_904, n_905, n_906, n_908, n_909, n_910, n_911, n_912;
wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
wire n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_931;
wire n_932, n_933, n_934, n_937, n_938, n_940, n_942, n_943;
wire n_946, n_947, n_948, n_950, n_952, n_954, n_955, n_956;
wire n_957, n_958, n_961, n_963, n_965, n_967, n_969, n_970;
wire n_971, n_973, n_974, n_975, n_976, n_977, n_978, n_980;
wire n_981, n_982, n_983, n_986, n_987, n_988, n_989, n_991;
wire n_992, n_993, n_994, n_995, n_998, n_999, n_1002, n_1011;
wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1021, n_1023, n_1024;
wire n_1040, n_1043, n_1044, n_1046, n_1052, n_1053, n_1054, n_1055;
wire n_1058, n_1059, n_1060, n_1062, n_1063, n_1064, n_1065, n_1069;
wire n_1071, n_1072, n_1074, n_1075, n_1077, n_1079, n_1081, n_1082;
wire n_1083, n_1084, n_1085, n_1090, n_1093, n_1094, n_1095, n_1096;
wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104;
wire n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112;
wire n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120;
wire n_1121, n_1122, n_1123, n_1124, n_1127, n_1128, n_1130, n_1131;
wire n_1133, n_1135, n_1136, n_1137, n_1138, n_1139, n_1143, n_1144;
wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1152, n_1153;
wire n_1154, n_1155, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1173;
wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189;
wire n_1191, n_1192, n_1193, n_1194, n_1195, n_1198, n_1199, n_1200;
wire n_1201, n_1202, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210;
wire n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1219;
wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227;
wire n_1228, n_1230, n_1231, n_1232, n_1234, n_1235, n_1236, n_1237;
wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
wire n_1246, n_1247, n_1248, n_1250, n_1251, n_1252, n_1255, n_1257;
wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267, n_1268;
wire n_1269, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
wire n_1278, n_1279, n_1282, n_1283, n_1285, n_1286, n_1290, n_1291;
wire n_1292, n_1293, n_1295, n_1296, n_1298, n_1299, n_1300, n_1304;
wire n_1307, n_1308, n_1310, n_1311, n_1312, n_1313, n_1315, n_1321;
wire n_1322, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
wire n_1349, n_1351, n_1352, n_1353, n_1354, n_1356, n_1363, n_1364;
wire n_1366, n_1367, n_1369, n_1370, n_1373, n_1375, n_1377, n_1380;
wire n_1381, n_1382, n_1384, n_1388, n_1390, n_1391, n_1392, n_1393;
wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
wire n_1402, n_1403, n_1404, n_1405, n_1407, n_1408, n_1409, n_1411;
wire n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419;
wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
wire n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446;
wire n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
wire n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462;
wire n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470;
wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478;
wire n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1486, n_1487;
wire n_1488, n_1491, n_1493, n_1494, n_1499, n_1500, n_1502, n_1503;
wire n_1505, n_1506, n_1507, n_1509, n_1510, n_1511, n_1514, n_1515;
wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523;
wire n_1524, n_1525, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532;
wire n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540;
wire n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548;
wire n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556;
wire n_1557, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1567;
wire n_1568, n_1569, n_1570, n_1571, n_1574, n_1575, n_1576, n_1578;
wire n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587;
wire n_1590, n_1591, n_1592, n_1597, n_1599, n_1605, n_1625, n_1626;
wire n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1636;
wire n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647;
wire n_1649, n_1650, n_1652, n_1655, n_1656, n_1657, n_1658, n_1662;
wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672;
wire n_1674, n_1675, n_1676, n_1677, n_1678, n_1680, n_1681, n_1682;
wire n_1686, n_1687, n_1688, n_1689, n_1691, n_1694, n_1695, n_1696;
wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705;
wire n_1706, n_1707, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714;
wire n_1715, n_1716, n_1717, n_1718, n_1719, n_1721, n_1722, n_1723;
wire n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731;
wire n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1740;
wire n_1741, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
wire n_1758, n_1759, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766;
wire n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1775;
wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1783, n_1785, n_1786;
wire n_1787, n_1788, n_1789, n_1791, n_1792, n_1793, n_1794, n_1795;
wire n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803;
wire n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811;
wire n_1812, n_1813, n_1814, n_1817, n_1818, n_1819, n_1820, n_1821;
wire n_1822, n_1826, n_1827, n_1830, n_1831, n_1832, n_1833, n_1838;
wire n_1839, n_1840, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847;
wire n_1848, n_1849, n_1850, n_1851, n_1854, n_1855, n_1857, n_1858;
wire n_1859, n_1860, n_1861, n_1862, n_1863, n_1865, n_1869, n_1875;
wire n_1882, n_1883, n_1884, n_1885, n_1887, n_1968, n_1969, n_1971;
wire n_1972, n_1975, n_1976, n_1977, n_1979, n_1980, n_1982, n_1985;
wire n_1986, n_1989, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996;
wire n_1997, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
wire n_2007, n_2008, n_2009, n_2011, n_2014, n_2015, n_2016, n_2017;
wire n_2018, n_2019, n_2020, n_2023, n_2024, n_2025, n_2027, n_2029;
wire n_2030, n_2031, n_2032, n_2034, n_2038, n_2039, n_2042, n_2043;
wire n_2044, n_2045, n_2046, n_2048, n_2049, n_2051, n_2053, n_2054;
wire n_2055, n_2056, n_2057, n_2060, n_2061, n_2062, n_2063, n_2064;
wire n_2065, n_2067, n_2068, n_2069, n_2070, n_2072, n_2077, n_2078;
wire n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086;
wire n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094;
wire n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2103;
wire n_2106, n_2107, n_2108, n_2110, n_2111, n_2113, n_2114, n_2115;
wire n_2116, n_2118, n_2119, n_2120, n_2121, n_2122, n_2126, n_2127;
wire n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135;
wire n_2137, n_2138, n_2140, n_2141, n_2143, n_2144, n_2145, n_2146;
wire n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155;
wire n_2156, n_2157, n_2159, n_2160, n_2161, n_2163, n_2165, n_2166;
wire n_2167, n_2168, n_2172, n_2173, n_2174, n_2176, n_2177, n_2178;
wire n_2180, n_2181, n_2182, n_2192, n_2203, n_2204, n_2205, n_2206;
wire n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2215, n_2216;
wire n_2218, n_2219, n_2221, n_2223, n_2224, n_2225, n_2227, n_2228;
wire n_2229, n_2230, n_2231, n_2233, n_2234, n_2237, n_2239, n_2241;
wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249;
wire n_2250, n_2252, n_2253, n_2254, n_2255, n_2256, n_2258, n_2259;
wire n_2260, n_2263, n_2264, n_2265, n_2266, n_2268, n_2269, n_2270;
wire n_2271, n_2272, n_2274, n_2276, n_2277, n_2278, n_2280, n_2281;
wire n_2283, n_2284, n_2285, n_2286, n_2288, n_2289, n_2290, n_2291;
wire n_2293, n_2294, n_2296, n_2298, n_2301, n_2302, n_2303, n_2304;
wire n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312;
wire n_2316, n_2319, n_2320, n_2321, n_2323, n_2324, n_2325, n_2326;
wire n_2327, n_2329, n_2331, n_2332, n_2334, n_2336, n_2338, n_2339;
wire n_2340, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2356, n_2361;
wire n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2370, n_2372;
wire n_2373, n_2374, n_2375, n_2376, n_2378, n_2379, n_2382, n_2385;
wire n_2387, n_2388, n_2389, n_2391, n_2392, n_2397, n_2398, n_2400;
wire n_2403, n_2406, n_2408, n_2409, n_2410, n_2413, n_2414, n_2415;
wire n_2416, n_2419, n_2421, n_2423, n_2425, n_2426, n_2427, n_2428;
wire n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436;
wire n_2437, n_2438, n_2439, n_2441, n_2442, n_2443, n_2444, n_2447;
wire n_2448, n_2449, n_2451, n_2452, n_2453, n_2454, n_2456, n_2457;
wire n_2458, n_2459, n_2460, n_2461, n_2463, n_2464, n_2465, n_2466;
wire n_2468, n_2469, n_2471, n_2472, n_2474, n_2475, n_2479, n_2480;
wire n_2481, n_2483, n_2484, n_2485, n_2486, n_2488, n_2491, n_2492;
wire n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500;
wire n_2501, n_2502, n_2503, n_2504, n_2506, n_2507, n_2509, n_2510;
wire n_2512, n_2514, n_2515, n_2517, n_2518, n_2519, n_2520, n_2521;
wire n_2522, n_2523, n_2524, n_2526, n_2528, n_2529, n_2530, n_2531;
wire n_2533, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2543;
wire n_2545, n_2546, n_2548, n_2550, n_2551, n_2554, n_2555, n_2556;
wire n_2557, n_2558, n_2559, n_2560, n_2562, n_2563, n_2564, n_2566;
wire n_2567, n_2572, n_2573, n_2574, n_2575, n_2577, n_2578, n_2579;
wire n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587;
wire n_2588, n_2589, n_2590, n_2592, n_2593, n_2594, n_2595, n_2597;
wire n_2598, n_2600, n_2601, n_2602, n_2603, n_2604, n_2606, n_2607;
wire n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615;
wire n_2616, n_2619, n_2624, n_2625, n_2628, n_2629, n_2630, n_2632;
wire n_2634, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2644;
wire n_2645, n_2646, n_2647, n_2648, n_2651, n_2652, n_2653, n_2654;
wire n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662;
wire n_2663, n_2664, n_2665, n_2666, n_2668, n_2669, n_2670, n_2671;
wire n_2672, n_2673, n_2675, n_2677, n_2678, n_2679, n_2680, n_2682;
wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2699, n_2700;
wire n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2709, n_2710;
wire n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2718, n_2719;
wire n_2720, n_2722, n_2723, n_2725, n_2727, n_2729, n_2730, n_2732;
wire n_2733, n_2734, n_2735, n_2736, n_2738, n_2739, n_2740, n_2741;
wire n_2742, n_2743, n_2744, n_2746, n_2747, n_2748, n_2749, n_2751;
wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
wire n_2761, n_2762, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769;
wire n_2770, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778;
wire n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2787;
wire n_2788, n_2789, n_2790, n_2791, n_2793, n_2794, n_2795, n_2796;
wire n_2797, n_2798, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805;
wire n_2806, n_2807, n_2808, n_2809, n_2810, n_2812, n_2813, n_2814;
wire n_2815, n_2816, n_2817, n_2819, n_2820, n_2821, n_2822, n_2823;
wire n_2824, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832;
wire n_2833, n_2834, n_2835, n_2837, n_2838, n_2839, n_2840, n_2841;
wire n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849;
wire n_2850, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858;
wire n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2866, n_2867;
wire n_2868, n_2869, n_2870, n_2871, n_2872, n_2875, n_2878, n_2879;
wire n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887;
wire n_2888, n_2889, n_2890, n_2891, n_2892, n_2894, n_2895, n_2896;
wire n_2897, n_2898, n_2900, n_2902, n_2903, n_2904, n_2905, n_2906;
wire n_2907, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915;
wire n_2917, n_2918, n_2920, n_2923, n_2924, n_2925, n_2926, n_2928;
wire n_2929, n_2930, n_2931, n_2933, n_2934, n_2936, n_2937, n_2938;
wire n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946;
wire n_2947, n_2948, n_2949, n_2951, n_2953, n_2954, n_2955, n_2956;
wire n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964;
wire n_2965, n_2966, n_2967, n_2968, n_2969, n_2971, n_2972, n_2973;
wire n_2974, n_2975, n_2977, n_2979, n_2980, n_2981, n_2983, n_2985;
wire n_2986, n_2987, n_2988, n_2989, n_2996, n_3001, n_3003, n_3004;
wire n_3005, n_3007, n_3008, n_3010, n_3011, n_3012, n_3013, n_3014;
wire n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022;
wire n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032;
wire n_3033, n_3034, n_3035, n_3036, n_3038, n_3040, n_3041, n_3042;
wire n_3043, n_3044, n_3047, n_3048, n_3049, n_3050, n_3052, n_3053;
wire n_3055, n_3056, n_3057, n_3058, n_3059, n_3062, n_3063, n_3065;
wire n_3066, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3077;
wire n_3079, n_3080, n_3081, n_3082, n_3084, n_3085, n_3086, n_3087;
wire n_3088, n_3090, n_3091, n_3092, n_3094, n_3095, n_3096, n_3097;
wire n_3098, n_3099, n_3100, n_3102, n_3103, n_3104, n_3105, n_3106;
wire n_3108, n_3109, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116;
wire n_3117, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3127;
wire n_3130, n_3131, n_3132, n_3133, n_3135, n_3136, n_3137, n_3138;
wire n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146;
wire n_3147, n_3148, n_3149, n_3152, n_3153, n_3154, n_3156, n_3157;
wire n_3158, n_3160, n_3161, n_3162, n_3164, n_3165, n_3167, n_3170;
wire n_3171, n_3172, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179;
wire n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3189;
wire n_3191, n_3192, n_3193, n_3194, n_3196, n_3197, n_3200, n_3201;
wire n_3202, n_3204, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211;
wire n_3212, n_3213, n_3214, n_3216, n_3217, n_3218, n_3219, n_3221;
wire n_3222, n_3223, n_3224, n_3225, n_3226, n_3228, n_3229, n_3233;
wire n_3234, n_3236, n_3239, n_3241, n_3242, n_3243, n_3244, n_3247;
wire n_3249, n_3253, n_3254, n_3255, n_3257, n_3258, n_3259, n_3260;
wire n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268;
wire n_3269, n_3270, n_3271, n_3273, n_3274, n_3275, n_3276, n_3277;
wire n_3278, n_3279, n_3281, n_3282, n_3283, n_3285, n_3286, n_3287;
wire n_3288, n_3289, n_3290, n_3291, n_3292, n_3296, n_3298, n_3299;
wire n_3300, n_3301, n_3302, n_3303, n_3305, n_3307, n_3308, n_3309;
wire n_3310, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3319;
wire n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327;
wire n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335;
wire n_3336, n_3337, n_3339, n_3340, n_3341, n_3343, n_3344, n_3345;
wire n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353;
wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362;
wire n_3363, n_3364, n_3365, n_3366, n_3368, n_3369, n_3370, n_3371;
wire n_3372, n_3373, n_3376, n_3377, n_3381, n_3382, n_3383, n_3384;
wire n_3385, n_3387, n_3388, n_3389, n_3390, n_3391, n_3394, n_3395;
wire n_3398, n_3399, n_3400, n_3402, n_3403, n_3404, n_3406, n_3407;
wire n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415;
wire n_3416, n_3417, n_3418, n_3420, n_3422, n_3423, n_3424, n_3425;
wire n_3426, n_3427, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434;
wire n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442;
wire n_3447, n_3448, n_3449, n_3454, n_3455, n_3458, n_3459, n_3460;
wire n_3461, n_3463, n_3464, n_3465, n_3466, n_3468, n_3469, n_3470;
wire n_3471, n_3473, n_3475, n_3477, n_3478, n_3479, n_3480, n_3481;
wire n_3482, n_3483, n_3484, n_3486, n_3487, n_3488, n_3489, n_3490;
wire n_3491, n_3492, n_3493, n_3494, n_3496, n_3497, n_3498, n_3499;
wire n_3500, n_3501, n_3502, n_3503, n_3505, n_3506, n_3507, n_3508;
wire n_3510, n_3511, n_3512, n_3514, n_3516, n_3517, n_3518, n_3519;
wire n_3520, n_3521, n_3522, n_3523, n_3529, n_3530, n_3531, n_3532;
wire n_3533, n_3534, n_3535, n_3537, n_3538, n_3540, n_3541, n_3542;
wire n_3543, n_3546, n_3547, n_3549, n_3550, n_3551, n_3552, n_3554;
wire n_3555, n_3557, n_3559, n_3560, n_3561, n_3563, n_3564, n_3566;
wire n_3567, n_3569, n_3570, n_3571, n_3572, n_3574, n_3577, n_3578;
wire n_3580, n_3581, n_3582, n_3585, n_3588, n_3589, n_3590, n_3591;
wire n_3592, n_3593, n_3596, n_3598, n_3599, n_3601, n_3603, n_3604;
wire n_3605, n_3606, n_3609, n_3611, n_3612, n_3613, n_3614, n_3615;
wire n_3616, n_3618, n_3620, n_3621, n_3622, n_3624, n_3625, n_3626;
wire n_3627, n_3628, n_3629, n_3631, n_3633, n_3634, n_3636, n_3637;
wire n_3638, n_3639, n_3640, n_3641, n_3642, n_3645, n_3646, n_3647;
wire n_3648, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3658;
wire n_3659, n_3660, n_3661, n_3662, n_3666, n_3670, n_3671, n_3672;
wire n_3673, n_3674, n_3675, n_3677, n_3679, n_3680, n_3681, n_3683;
wire n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692;
wire n_3693, n_3695, n_3697, n_3700, n_3701, n_3702, n_3703, n_3706;
wire n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3715;
wire n_3716, n_3717, n_3718, n_3720, n_3721, n_3722, n_3723, n_3724;
wire n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732;
wire n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3740, n_3742;
wire n_3744, n_3745, n_3746, n_3752, n_3753, n_3755, n_3758, n_3761;
wire n_3764, n_3765, n_3766, n_3767, n_3769, n_3770, n_3771, n_3774;
wire n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782;
wire n_3784, n_3785, n_3786, n_3788, n_3789, n_3792, n_3793, n_3795;
wire n_3797, n_3798, n_3800, n_3801, n_3802, n_3803, n_3807, n_3808;
wire n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816;
wire n_3817, n_3819, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826;
wire n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835;
wire n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3843, n_3844;
wire n_3845, n_3846, n_3847, n_3848, n_3849, n_3851, n_3852, n_3854;
wire n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3863;
wire n_3866, n_3868, n_3869, n_3870, n_3873, n_3877, n_3878, n_3879;
wire n_3881, n_3882, n_3883, n_3885, n_3886, n_3891, n_3893, n_3894;
wire n_3895, n_3896, n_3897, n_3898, n_3900, n_3902, n_3903, n_3904;
wire n_3905, n_3906, n_3907, n_3910, n_3911, n_3913, n_3914, n_3915;
wire n_3916, n_3922, n_3925, n_3929, n_3932, n_3933, n_3934, n_3936;
wire n_3937, n_3938, n_3939, n_3941, n_3942, n_3943, n_3944, n_3945;
wire n_3946, n_3947, n_3948, n_3949, n_3951, n_3952, n_3953, n_3955;
wire n_3956, n_3957, n_3958, n_3959, n_3960, n_3962, n_3963, n_3964;
wire n_3966, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974;
wire n_3977, n_3978, n_3979, n_3981, n_3982, n_3983, n_3984, n_3985;
wire n_3990, n_3991, n_3992, n_3993, n_3995, n_3996, n_3997, n_3998;
wire n_4000, n_4002, n_4005, n_4006, n_4008, n_4009, n_4010, n_4011;
wire n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019;
wire n_4020, n_4021, n_4022, n_4024, n_4025, n_4028, n_4029, n_4030;
wire n_4031, n_4032, n_4033, n_4034, n_4035, n_4037, n_4038, n_4040;
wire n_4042, n_4043, n_4044, n_4045, n_4046, n_4048, n_4049, n_4050;
wire n_4053, n_4054, n_4055, n_4056, n_4059, n_4060, n_4062, n_4065;
wire n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073;
wire n_4074, n_4076, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085;
wire n_4086, n_4087, n_4088, n_4090, n_4091, n_4092, n_4096, n_4098;
wire n_4101, n_4102, n_4103, n_4105, n_4107, n_4108, n_4109, n_4110;
wire n_4111, n_4113, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122;
wire n_4123, n_4124, n_4125, n_4126, n_4131, n_4133, n_4134, n_4135;
wire n_4136, n_4137, n_4139, n_4140, n_4142, n_4145, n_4147, n_4148;
wire n_4149, n_4150, n_4151, n_4152, n_4154, n_4155, n_4156, n_4157;
wire n_4159, n_4160, n_4161, n_4163, n_4165, n_4167, n_4168, n_4169;
wire n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177;
wire n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185;
wire n_4186, n_4187, n_4188, n_4189, n_4190, n_4192, n_4193, n_4194;
wire n_4196, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204;
wire n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212;
wire n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220;
wire n_4221, n_4223, n_4224, n_4225, n_4226, n_4227, n_4230, n_4231;
wire n_4232, n_4233, n_4235, n_4237, n_4238, n_4239, n_4241, n_4242;
wire n_4243, n_4246, n_4247, n_4248, n_4250, n_4251, n_4252, n_4253;
wire n_4254, n_4255, n_4257, n_4260, n_4262, n_4263, n_4264, n_4265;
wire n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273;
wire n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281;
wire n_4282, n_4283, n_4284, n_4285, n_4286, n_4288, n_4290, n_4291;
wire n_4293, n_4296, n_4297, n_4298, n_4299, n_4301, n_4302, n_4303;
wire n_4304, n_4305, n_4306, n_4308, n_4313, n_4314, n_4315, n_4316;
wire n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324;
wire n_4325, n_4327, n_4328, n_4329, n_4330, n_4331, n_4333, n_4336;
wire n_4338, n_4339, n_4340, n_4343, n_4344, n_4345, n_4346, n_4347;
wire n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355;
wire n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363;
wire n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371;
wire n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379;
wire n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387;
wire n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395;
wire n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403;
wire n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411;
wire n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419;
wire n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427;
wire n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4436;
wire n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4444, n_4445;
wire n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453;
wire n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461;
wire n_4462, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470;
wire n_4471, n_4472, n_4473, n_4474, n_4475, n_4477, n_4478, n_4479;
wire n_4481, n_4482, n_4483, n_4485, n_4486, n_4487, n_4488, n_4489;
wire n_4490, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498;
wire n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4506, n_4507;
wire n_4508, n_4510, n_4512, n_4513, n_4514, n_4515, n_4516, n_4518;
wire n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526;
wire n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534;
wire n_4535, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4545;
wire n_4546, n_4547, n_4550, n_4553, n_4554, n_4555, n_4556, n_4557;
wire n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565;
wire n_4566, n_4567, n_4568, n_4569, n_4570, n_4572, n_4573, n_4574;
wire n_4575, n_4576, n_4577, n_4578, n_4579, n_4581, n_4582, n_4583;
wire n_4584, n_4585, n_4586, n_4587, n_4589, n_4590, n_4591, n_4592;
wire n_4593, n_4594, n_4597, n_4598, n_4600, n_4603, n_4605, n_4607;
wire n_4611, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620;
wire n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628;
wire n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4636, n_4637;
wire n_4638, n_4639, n_4640, n_4642, n_4645, n_4647, n_4649, n_4650;
wire n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658;
wire n_4659, n_4660, n_4661, n_4662, n_4663, n_4665, n_4666, n_4667;
wire n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4676, n_4677;
wire n_4678, n_4679, n_4680, n_4682, n_4683, n_4684, n_4688, n_4689;
wire n_4690, n_4693, n_4695, n_4699, n_4700, n_4704, n_4705, n_4706;
wire n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714;
wire n_4715, n_4716, n_4717, n_4719, n_4721, n_4723, n_4725, n_4726;
wire n_4727, n_4730, n_4731, n_4732, n_4734, n_4735, n_4736, n_4737;
wire n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4746;
wire n_4747, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756;
wire n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764;
wire n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4772, n_4773;
wire n_4774, n_4775, n_4776, n_4777, n_4779, n_4780, n_4781, n_4782;
wire n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790;
wire n_4791, n_4792, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799;
wire n_4800, n_4803, n_4804, n_4805, n_4806, n_4809, n_4810, n_4811;
wire n_4812, n_4813, n_4815, n_4820, n_4821, n_4822, n_4823, n_4824;
wire n_4827, n_4828, n_4829, n_4830, n_4832, n_4833, n_4834, n_4835;
wire n_4836, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844;
wire n_4845, n_4846, n_4847, n_4849, n_4850, n_4851, n_4852, n_4853;
wire n_4854, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4864;
wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4874, n_4875;
wire n_4876, n_4877, n_4878, n_4879, n_4881, n_4884, n_4885, n_4886;
wire n_4887, n_4888, n_4889, n_4891, n_4893, n_4896, n_4897, n_4898;
wire n_4899, n_4900, n_4904, n_4905, n_4906, n_4907, n_4911, n_4912;
wire n_4913, n_4915, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922;
wire n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930;
wire n_4931, n_4934, n_4935, n_4936, n_4939, n_4940, n_4942, n_4943;
wire n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951;
wire n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4959, n_4960;
wire n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968;
wire n_4969, n_4970, n_4971, n_4972, n_4974, n_4975, n_4976, n_4977;
wire n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985;
wire n_4986, n_4987, n_4988, n_4990, n_4991, n_4996, n_4999, n_5000;
wire n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008;
wire n_5009, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018;
wire n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026;
wire n_5028, n_5029, n_5030, n_5032, n_5033, n_5034, n_5035, n_5037;
wire n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045;
wire n_5046, n_5047, n_5048, n_5050, n_5051, n_5052, n_5053, n_5055;
wire n_5056, n_5057, n_5058, n_5059, n_5060, n_5062, n_5063, n_5064;
wire n_5065, n_5067, n_5068, n_5069, n_5071, n_5072, n_5073, n_5075;
wire n_5076, n_5077, n_5079, n_5081, n_5082, n_5083, n_5084, n_5085;
wire n_5086, n_5087, n_5088, n_5090, n_5091, n_5092, n_5093, n_5094;
wire n_5095, n_5097, n_5098, n_5100, n_5101, n_5103, n_5104, n_5106;
wire n_5107, n_5109, n_5110, n_5111, n_5112, n_5113, n_5115, n_5116;
wire n_5118, n_5119, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126;
wire n_5127, n_5128, n_5129, n_5130, n_5131, n_5133, n_5134, n_5135;
wire n_5136, n_5137, n_5139, n_5141, n_5143, n_5144, n_5146, n_5148;
wire n_5149, n_5150, n_5151, n_5152, n_5154, n_5155, n_5156, n_5158;
wire n_5159, n_5160, n_5161, n_5163, n_5164, n_5165, n_5167, n_5168;
wire n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5177, n_5179;
wire n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5189;
wire n_5190, n_5192, n_5193, n_5195, n_5197, n_5199, n_5200, n_5201;
wire n_5202, n_5204, n_5205, n_5206, n_5207, n_5209, n_5210, n_5212;
wire n_5213, n_5214, n_5215, n_5218, n_5219, n_5221, n_5222, n_5223;
wire n_5224, n_5225, n_5226, n_5227, n_5229, n_5230, n_5231, n_5232;
wire n_5233, n_5235, n_5236, n_5238, n_5239, n_5240, n_5241, n_5242;
wire n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5251, n_5252;
wire n_5253, n_5254, n_5258, n_5259, n_5265, n_5266, n_5267, n_5268;
wire n_5270, n_5271, n_5272, n_5273, n_5275, n_5276, n_5278, n_5279;
wire n_5282, n_5283, n_5284, n_5287, n_5288, n_5289, n_5290, n_5291;
wire n_5293, n_5294, n_5296, n_5297, n_5299, n_5300, n_5302, n_5304;
wire n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313;
wire n_5315, n_5317, n_5318, n_5319, n_5321, n_5323, n_5324, n_5325;
wire n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5333, n_5335;
wire n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5344;
wire n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5352, n_5353;
wire n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5361, n_5362;
wire n_5363, n_5364, n_5365, n_5369, n_5370, n_5372, n_5373, n_5374;
wire n_5375, n_5377, n_5378, n_5379, n_5380, n_5382, n_5383, n_5384;
wire n_5385, n_5386, n_5387, n_5388, n_5391, n_5392, n_5393, n_5394;
wire n_5395, n_5396, n_5397, n_5398, n_5400, n_5402, n_5403, n_5404;
wire n_5405, n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412;
wire n_5414, n_5415, n_5420, n_5422, n_5423, n_5424, n_5425, n_5428;
wire n_5430, n_5431, n_5432, n_5436, n_5437, n_5440, n_5442, n_5444;
wire n_5445, n_5447, n_5448, n_5449, n_5450, n_5451, n_5453, n_5454;
wire n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462;
wire n_5464, n_5465, n_5466, n_5467, n_5468, n_5471, n_5474, n_5476;
wire n_5481, n_5483, n_5485, n_5486, n_5487, n_5489, n_5490, n_5492;
wire n_5495, n_5497, n_5499, n_5500, n_5501, n_5502, n_5504, n_5505;
wire n_5506, n_5508, n_5513, n_5514, n_5515, n_5517, n_5518, n_5519;
wire n_5520, n_5521, n_5522, n_5524, n_5526, n_5527, n_5529, n_5530;
wire n_5531, n_5532, n_5534, n_5536, n_5537, n_5538, n_5539, n_5540;
wire n_5541, n_5542, n_5543, n_5544, n_5547, n_5549, n_5553, n_5556;
wire n_5557, n_5559, n_5560, n_5562, n_5563, n_5564, n_5565, n_5566;
wire n_5567, n_5568, n_5569, n_5570, n_5571, n_5573, n_5574, n_5575;
wire n_5576, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584;
wire n_5587, n_5590, n_5591, n_5592, n_5593, n_5596, n_5599, n_5600;
wire n_5602, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613;
wire n_5614, n_5615, n_5617, n_5619, n_5622, n_5624, n_5625, n_5626;
wire n_5627, n_5629, n_5630, n_5631, n_5633, n_5634, n_5637, n_5639;
wire n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5650;
wire n_5652, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660;
wire n_5661, n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668;
wire n_5669, n_5671, n_5672, n_5674, n_5675, n_5676, n_5677, n_5678;
wire n_5680, n_5681, n_5683, n_5686, n_5688, n_5689, n_5690, n_5692;
wire n_5693, n_5694, n_5695, n_5700, n_5701, n_5702, n_5703, n_5704;
wire n_5705, n_5707, n_5709, n_5711, n_5712, n_5714, n_5715, n_5716;
wire n_5718, n_5719, n_5720, n_5723, n_5724, n_5725, n_5726, n_5727;
wire n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735;
wire n_5736, n_5737, n_5738, n_5740, n_5741, n_5742, n_5743, n_5744;
wire n_5745, n_5746, n_5749, n_5755, n_5756, n_5757, n_5758, n_5759;
wire n_5760, n_5761, n_5762, n_5765, n_5767, n_5768, n_5769, n_5772;
wire n_5774, n_5775, n_5776, n_5777, n_5779, n_5780, n_5781, n_5782;
wire n_5784, n_5786, n_5788, n_5790, n_5792, n_5794, n_5795, n_5796;
wire n_5797, n_5798, n_5799, n_5800, n_5801, n_5803, n_5804, n_5805;
wire n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5813, n_5814;
wire n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822;
wire n_5824, n_5825, n_5828, n_5830, n_5831, n_5833, n_5837, n_5839;
wire n_5844, n_5849, n_5852, n_5854, n_5857, n_5859, n_5860, n_5862;
wire n_5863, n_5865, n_5866, n_5868, n_5869, n_5870, n_5871, n_5872;
wire n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880;
wire n_5881, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888;
wire n_5889, n_5891, n_5896, n_5899, n_5901, n_5904, n_5905, n_5906;
wire n_5907, n_5908, n_5909, n_5910, n_5913, n_5914, n_5916, n_5917;
wire n_5918, n_5920, n_5921, n_5922, n_5924, n_5925, n_5926, n_5927;
wire n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935;
wire n_5936, n_5937, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944;
wire n_5945, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953;
wire n_5954, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962;
wire n_5964, n_5965, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972;
wire n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5981;
wire n_5982, n_5983, n_5984, n_5985, n_5986, n_5988, n_5991, n_5992;
wire n_5993, n_5994, n_5995, n_5996, n_5997, n_5999, n_6000, n_6001;
wire n_6002, n_6003, n_6004, n_6005, n_6006, n_6008, n_6009, n_6010;
wire n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018;
wire n_6019, n_6020, n_6021, n_6024, n_6025, n_6026, n_6027, n_6028;
wire n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036;
wire n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044;
wire n_6045, n_6046, n_6048, n_6049, n_6050, n_6051, n_6052, n_6054;
wire n_6055, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6064;
wire n_6065, n_6066, n_6067, n_6068, n_6070, n_6071, n_6072, n_6073;
wire n_6074, n_6076, n_6078, n_6079, n_6080, n_6081, n_6082, n_6084;
wire n_6086, n_6087, n_6089, n_6091, n_6092, n_6093, n_6094, n_6095;
wire n_6096, n_6098, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105;
wire n_6107, n_6108, n_6109, n_6110, n_6111, n_6112, n_6114, n_6116;
wire n_6117, n_6118, n_6120, n_6121, n_6123, n_6125, n_6126, n_6128;
wire n_6129, n_6130, n_6132, n_6133, n_6134, n_6136, n_6137, n_6138;
wire n_6140, n_6141, n_6142, n_6143, n_6145, n_6146, n_6149, n_6150;
wire n_6153, n_6154, n_6155, n_6156, n_6157, n_6160, n_6161, n_6162;
wire n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6171, n_6174;
wire n_6176, n_6178, n_6180, n_6182, n_6183, n_6184, n_6185, n_6186;
wire n_6188, n_6189, n_6190, n_6192, n_6194, n_6197, n_6198, n_6199;
wire n_6201, n_6202, n_6203, n_6204, n_6206, n_6207, n_6208, n_6209;
wire n_6210, n_6211, n_6214, n_6216, n_6217, n_6218, n_6220, n_6221;
wire n_6222, n_6223, n_6224, n_6225, n_6226, n_6228, n_6229, n_6230;
wire n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239;
wire n_6240, n_6241, n_6243, n_6246, n_6247, n_6248, n_6250, n_6252;
wire n_6253, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259, n_6260;
wire n_6262, n_6264, n_6265, n_6266, n_6267, n_6271, n_6274, n_6275;
wire n_6279, n_6280, n_6281, n_6282, n_6283, n_6285, n_6286, n_6287;
wire n_6288, n_6290, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300;
wire n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6308, n_6309;
wire n_6310, n_6311, n_6312, n_6313, n_6315, n_6316, n_6317, n_6318;
wire n_6320, n_6321, n_6323, n_6324, n_6326, n_6327, n_6328, n_6330;
wire n_6331, n_6332, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339;
wire n_6342, n_6345, n_6346, n_6347, n_6348, n_6351, n_6352, n_6353;
wire n_6355, n_6356, n_6357, n_6359, n_6360, n_6361, n_6362, n_6363;
wire n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371;
wire n_6372, n_6373, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380;
wire n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6388, n_6389;
wire n_6390, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398;
wire n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, n_6406;
wire n_6407, n_6408, n_6409, n_6410, n_6411, n_6412, n_6413, n_6414;
wire n_6415, n_6416, n_6417, n_6418, n_6419, n_6421, n_6422, n_6454;
wire n_6457, n_6460, n_6464, n_6468, n_6479, n_6488, n_6490, n_6501;
wire n_6503, n_6504, n_6506, n_6507, n_6508, n_6517, n_6522, n_6523;
wire n_6524, n_6527, n_6539, n_6545, n_6547, n_6548, n_6549, n_6551;
wire n_6552, n_6553, n_6562, n_6564, n_6565, n_6570, n_6572, n_6574;
wire n_6577, n_6578, n_6582, n_6584, n_6610, n_6612, n_6618, n_6620;
wire n_6621, n_6631, n_6639, n_6655, n_6663, n_6664, n_6666, n_6668;
wire n_6669, n_6670, n_6673, n_6676, n_6677, n_6679, n_6680, n_6683;
wire n_6684, n_6685, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692;
wire n_6693, n_6694, n_6695, n_6696, n_6697, n_6705, n_6707, n_6714;
wire n_6715, n_6716, n_6734, n_6735, n_6742, n_6746, n_6752, n_6754;
wire n_6755, n_6756, n_6757, n_6758, n_6759, n_6760, n_6762, n_6764;
wire n_6765, n_6766, n_6767, n_6781, n_6782, n_6785, n_6786, n_6787;
wire n_6788, n_6789, n_6790, n_6791, n_6794, n_6796, n_6798, n_6799;
wire n_6800, n_6801, n_6806, n_6807, n_6808, n_6809, n_6821, n_6822;
wire n_6823, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853, n_6854;
wire n_6856, n_6857, n_6858, n_6864, n_6865, n_6866, n_6872, n_6876;
wire n_6877, n_6878, n_6880, n_6891, n_6892, n_6893, n_6895, n_6896;
wire n_6897, n_6898, n_6899, n_6903, n_6906, n_6907, n_6922, n_6923;
wire n_6925, n_6926, n_6927, n_6928, n_6937, n_6938, n_6940, n_6941;
wire n_6948, n_6951, n_6953, n_6954, n_6956, n_6958, n_6967, n_6970;
wire n_6972, n_6973, n_6978, n_6979, n_7003, n_7004, n_7010, n_7018;
wire n_7022, n_7023, n_7024, n_7025, n_7032, n_7039, n_7040, n_7042;
wire n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049, n_7085;
wire n_7086, n_7087, n_7088, n_7089, n_7090, n_7093, n_7094, n_7097;
wire n_7099, n_7101, n_7102, n_7103, n_7105, n_7116, n_7118, n_7119;
wire n_7120, n_7121, n_7122, n_7123, n_7124, n_7127, n_7128, n_7130;
wire n_7131, n_7132, n_7133, n_7140, n_7141, n_7142, n_7143, n_7144;
wire n_7145, n_7146, n_7150, n_7164, n_7165, n_7167, n_7168, n_7208;
wire n_7213, n_7214, n_7217, n_7218, n_7219, n_7229, n_7235, n_7242;
wire n_7243, n_7245, n_7247, n_7260, n_7268, n_7275, n_7320, n_7321;
wire n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328, n_7329;
wire n_7330, n_7331, n_7332, n_7333, n_7343, n_7344, n_7348, n_7352;
wire n_7353, n_7354, n_7383, n_7395, n_7402, n_8508, n_8509, n_8532;
wire n_8534, n_8537, n_8540, n_8546, n_8547, n_8548, n_8552, n_8555;
wire n_8556, n_8557, n_8571, n_8572, n_8582, n_8583, n_8584, n_8585;
wire n_8586, n_8587, n_8588, n_8589, n_8591, n_8594, n_8599, n_8600;
wire n_8601, n_8603, n_8604, n_8605, n_8609, n_8610, n_8611, n_8615;
wire n_8616, n_8618, n_8619, n_8620, n_8627, n_8628, n_8629, n_8632;
wire n_8633, n_8634, n_8637, n_8638, n_8639, n_8675, n_8676, n_8677;
wire n_8678, n_8679, n_8680, n_8681, n_8682, n_8686, n_8687, n_8690;
wire n_8691, n_8693, n_8694, n_8697, n_8702, n_8703, n_8704, n_8705;
wire n_8706, n_8707, n_8730, n_8731, n_8733, n_8734, n_8735, n_8736;
wire n_8755, n_8756, n_8757, n_8758, n_8759, n_8761, n_8762, n_8763;
wire n_8764, n_8768, n_8769, n_8770, n_8776, n_8777, n_8778, n_8792;
wire n_8793, n_8796, n_8799, n_8800, n_8806, n_8807, n_8809, n_8810;
wire n_8816, n_8817, n_8818, n_8819, n_8820, n_8821, n_8831, n_8832;
wire n_8833, n_8834, n_8835, n_8836, n_8837, n_8839, n_8840, n_8846;
wire n_8848, n_8850, n_8855, n_8864, n_8879, n_8880, n_8882, n_8883;
wire n_8885, n_8886, n_8895, n_8898, n_8906, n_8908, n_8909, n_8913;
wire n_8915, n_8917, n_8921, n_8955, n_9000, n_9019, n_9091, n_9107;
wire n_9129, n_9139, n_9141, n_9156, n_9167, n_9172, n_9176, n_9193;
wire n_9209, n_9218, n_9234, n_9240, n_9256, n_9269, n_9279, n_9297;
wire n_9300, n_9311, n_9333, n_9351, n_9353, n_9358, n_9359, n_9371;
wire n_9398, n_9404, n_9419, n_9422, n_9425, n_9431, n_9443, n_9448;
wire n_9453, n_9454, n_9461, n_9466, n_9469, n_9491, n_9493, n_9501;
wire n_9505, n_9521, n_9526, n_9553, n_9558, n_9599, n_9627, n_9628;
wire n_9630, n_9651, n_9664, n_9672, n_9681, n_9693, n_9697, n_9698;
wire n_9717, n_9750, n_9772, n_9775, n_9797, n_9811, n_9830, n_9834;
wire n_9836, n_9856, n_9862, n_9871, n_9874, n_9883, n_9884, n_9894;
wire n_9903, n_9928, n_9940, n_9952, n_9976, n_9978, n_9992, n_10005;
wire n_10013, n_10063, n_10078, n_10097, n_10099, n_10100, n_10101,n_10103;
wire n_10107, n_10108, n_10112, n_10113, n_10115, n_10119, n_10120,n_10123;
wire n_10125, n_10128, n_10129, n_10134, n_10139, n_10142, n_10173,n_10175;
wire n_10176, n_10177, n_10180, n_10181, n_10184, n_10185, n_10188,n_10192;
wire n_10196, n_10197, n_10199, n_10200, n_10201, n_10202, n_10203,n_10205;
wire n_10206, n_10213, n_10214, n_10216, n_10217, n_10224, n_10225,n_10226;
wire n_10227, n_10228, n_10229, n_10238, n_10239, n_10240, n_10241,n_10242;
wire n_10243, n_10245, n_10247, n_10257, n_10259, n_10260, n_10261,n_10262;
wire n_10263, n_10264, n_10268, n_10270, n_10271, n_10280, n_10281,n_10282;
wire n_10283, n_10285, n_10286, n_10287, n_10288, n_10289, n_10290,n_10296;
wire n_10303, n_10304, n_10306, n_10307, n_10308, n_10309, n_10310,n_10311;
wire n_10312, n_10313, n_10314, n_10315, n_10316, n_10317, n_10318,n_10319;
wire n_10320, n_10321, n_10322, n_10323, n_10325, n_10327, n_10328,n_10329;
wire n_10330, n_10341, n_10342, n_10343, n_10344, n_10345, n_10346,n_10347;
wire n_10357, n_10361, n_10362, n_10363, n_10368, n_10369, n_10371,n_10372;
wire n_10373, n_10374, n_10376, n_10377, n_10378, n_10379, n_10380,n_10381;
wire n_10382, n_10383, n_10385, n_10386, n_10387, n_10388, n_10390,n_10391;
wire n_10392, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399,n_10400;
wire n_10401, n_10402, n_10404, n_10411, n_10412, n_10413, n_10414,n_10415;
wire n_10416, n_10422, n_10423, n_10424, n_10425, n_10426, n_10427,n_10428;
wire n_10429, n_10430, n_10431, n_10443, n_10444, n_10445, n_10446,n_10447;
wire n_10448, n_10460, n_10461, n_10462, n_10463, n_10464, n_10466,n_10467;
wire n_10470, n_10472, n_10473, n_10475, n_10494, n_10495, n_10496,n_10499;
wire n_10503, n_10504, n_10505, n_10506, n_10508, n_10512, n_10513,n_10514;
wire n_10515, n_10516, n_10517, n_10518, n_10519, n_10520, n_10522,n_10524;
wire n_10525, n_10526, n_10527, n_10528, n_10529, n_10532, n_10534,n_10535;
wire n_10548, n_10549, n_10550, n_10551, n_10552, n_10553, n_10554,n_10557;
wire n_10558, n_10560, n_10563, n_10564, n_10565, n_10566, n_10567,n_10568;
wire n_10569, n_10573, n_10576, n_10577, n_10578, n_10579, n_10580,n_10581;
wire n_10582, n_10587, n_10588, n_10589, n_10590, n_10595, n_10596,n_10597;
wire n_10598, n_10599, n_10600, n_10601, n_10607, n_10609, n_10613,n_10614;
wire n_10616, n_10617, n_10618, n_10620, n_10621, n_10622, n_10623,n_10624;
wire n_10625, n_10626, n_10628, n_10630, n_10631, n_10632, n_10633,n_10634;
wire n_10637, n_10638, n_10639, n_10644, n_10647, n_10649, n_10650,n_10656;
wire n_10657, n_10660, n_10664, n_10667, n_10669, n_10670, n_10671,n_10672;
wire n_10674, n_10675, n_10678, n_10682, n_10683, n_10684, n_10685,n_10686;
wire n_10687, n_10689, n_10690, n_10693, n_10694, n_10695, n_10696,n_10697;
wire n_10698, n_10699, n_10700, n_10708, n_10709, n_10710, n_10713,n_10714;
wire n_10715, n_10716, n_10717, n_10718, n_10720, n_10723, n_10724,n_10725;
wire n_10745, n_10746, n_10747, n_10748, n_10749, n_10750, n_10751,n_10752;
wire n_10753, n_10754, n_10755, n_10756, n_10758, n_10759, n_10760,n_10761;
wire n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768,n_10769;
wire n_10770, n_10771, n_10772, n_10773, n_10781, n_10782, n_10785,n_10787;
wire n_10789, n_10790, n_10801, n_10802, n_10803, n_10804, n_10805,n_10806;
wire n_10808, n_10809, n_10813, n_10814, n_10818, n_10823, n_10826,n_10827;
wire n_10829, n_10830, n_10831, n_10833, n_10834, n_10839, n_10841,n_10846;
wire n_10852, n_10853, n_10854, n_10856, n_10857, n_10861, n_10863,n_10867;
wire n_10871, n_10873, n_10874, n_10877, n_10879, n_10883, n_10889,n_10893;
wire n_10894, n_10895, n_10897, n_10898, n_10899, n_10901, n_10903,n_10905;
wire n_10906, n_10907, n_10910, n_10911, n_10912, n_10913, n_10915,n_10916;
wire n_10917, n_10920, n_10921, n_10932, n_10934, n_10936, n_10937,n_10939;
wire n_10940, n_10941, n_10942, n_10943, n_10944, n_10947, n_10948,n_10949;
wire n_10950, n_10951, n_10952, n_10953, n_10954, n_10955, n_10956,n_10959;
wire n_10960, n_10961, n_10962, n_10963, n_10964, n_10965, n_10966,n_10967;
wire n_10968, n_10969, n_10970, n_10971, n_10972, n_10973, n_10974,n_10975;
wire n_10976, n_10978, n_10980, n_10981, n_10982, n_10983, n_10984,n_10986;
wire n_10987, n_10988, n_10989, n_10991, n_10992, n_10993, n_10994,n_10995;
wire n_10996, n_10997, n_10998, n_11012, n_11013, n_11025, n_11026,n_11027;
wire n_11028, n_11029, n_11030, n_11031, n_11032, n_11033, n_11034,n_11035;
wire n_11036, n_11037, n_11038, n_11039, n_11040, n_11041, n_11042,n_11045;
wire n_11050, n_11051, n_11055, n_11056, n_11064, n_11065, n_11070,n_11071;
wire n_11073, n_11076, n_11077, n_11079, n_11080, n_11081, n_11088,n_11091;
wire n_11094, n_11095, n_11097, n_11099, n_11101, n_11104, n_11105,n_11106;
wire n_11110, n_11113, n_11116, n_11118, n_11119, n_11120, n_11121,n_11122;
wire n_11124, n_11126, n_11128, n_11129, n_11133, n_11134, n_11138,n_11150;
wire n_11157, n_11160, n_11162, n_11163, n_11165, n_11171, n_11173,n_11177;
wire n_11178, n_11184, n_11185, n_11186, n_11187, n_11188, n_11189,n_11190;
wire n_11191, n_11192, n_11193, n_11194, n_11195, n_11196, n_11197,n_11198;
wire n_11201, n_11203, n_11205, n_11206, n_11207, n_11208, n_11209,n_11210;
wire n_11211, n_11212, n_11216, n_11217, n_11218, n_11219, n_11220,n_11221;
assign g34972 = 1'b1;
assign g34956 = g34839;
assign g34927 = 1'b1;
assign g34925 = 1'b1;
assign g34923 = 1'b1;
assign g34921 = 1'b1;
assign g34919 = 1'b1;
assign g34917 = 1'b1;
assign g34915 = 1'b1;
assign g34913 = 1'b1;
assign g34788 = g33894;
assign g34597 = 1'b0;
assign g34437 = 1'b1;
assign g34436 = 1'b1;
assign g34435 = g31521;
assign g34425 = 1'b1;
assign g34383 = 1'b1;
assign g34240 = 1'b1;
assign g34239 = 1'b1;
assign g34238 = 1'b1;
assign g34237 = 1'b1;
assign g34236 = 1'b1;
assign g34235 = 1'b1;
assign g34234 = 1'b1;
assign g34233 = 1'b1;
assign g34232 = 1'b1;
assign g34221 = 1'b1;
assign g34201 = 1'b1;
assign g33959 = g28753;
assign g33950 = 1'b1;
assign g33949 = 1'b1;
assign g33948 = 1'b1;
assign g33947 = 1'b1;
assign g33946 = 1'b1;
assign g33945 = 1'b1;
assign g33935 = 1'b1;
assign g33874 = 1'b1;
assign g33659 = 1'b1;
assign g33636 = 1'b1;
assign g33533 = g27831;
assign g32975 = g26801;
assign g32454 = 1'b1;
assign g32429 = 1'b1;
assign g31863 = g25167;
assign g31862 = g25259;
assign g31861 = g25219;
assign g31860 = g25114;
assign g31665 = 1'b1;
assign g31656 = 1'b1;
assign g30332 = g23683;
assign g30331 = g23759;
assign g30330 = g23652;
assign g30329 = g23612;
assign g30327 = g23002;
assign g29221 = g21292;
assign g29220 = g21245;
assign g29219 = g20654;
assign g29218 = g18881;
assign g29217 = g21270;
assign g29216 = g21176;
assign g29215 = g20901;
assign g29214 = g20652;
assign g29213 = g20557;
assign g29212 = g20899;
assign g29211 = g20763;
assign g29210 = g20049;
assign g25590 = 1'b1;
assign g25589 = 1'b1;
assign g25588 = 1'b1;
assign g25587 = 1'b1;
assign g25586 = 1'b1;
assign g25585 = 1'b1;
assign g25584 = 1'b1;
assign g25583 = 1'b1;
assign g25582 = 1'b1;
assign g24151 = 1'b1;
assign g23190 = 1'b1;
assign g21698 = g36;
assign g18101 = g6746;
assign g18100 = g6751;
assign g18099 = g6745;
assign g18098 = g6744;
assign g18097 = g6747;
assign g18096 = g6750;
assign g18095 = g6749;
assign g18094 = g6748;
assign g18092 = g6753;
assign g12368 = 1'b0;
assign g9048 = 1'b0;
assign g8403 = 1'b0;
assign g8353 = 1'b0;
assign g8283 = 1'b0;
assign g8235 = 1'b0;
assign g8178 = 1'b0;
assign g8132 = 1'b0;
DFFSRX1 g2955_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6422), .Q (g2955), .QN ());
MX2X1 g60853(.A (g2941), .B (n_6417), .S0 (n_8955), .Y (n_6422));
DFFSRX1 g2864_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6419), .Q (), .QN (g2864));
NAND3X1 g60850(.A (n_6418), .B (n_6408), .C (n_6416), .Y (g31793));
MX2X1 g60856(.A (n_3499), .B (n_6415), .S0 (n_9000), .Y (n_6419));
NOR2X1 g60852(.A (n_6411), .B (n_6412), .Y (n_6418));
NAND4X1 g60857(.A (n_6414), .B (n_2449), .C (n_3614), .D (n_3498), .Y(n_6417));
AOI21X1 g60855(.A0 (n_6394), .A1 (n_6401), .B0 (n_6410), .Y (n_6416));
OR2X1 g60860(.A (n_6413), .B (n_271), .Y (n_6415));
NOR2X1 g60861(.A (n_3502), .B (n_6413), .Y (n_6414));
OAI33X1 g60854(.A0 (n_1414), .A1 (n_6409), .A2 (n_901), .B0 (n_1454),.B1 (n_6397), .B2 (n_3812), .Y (n_6412));
NAND3X1 g60858(.A (n_6405), .B (n_6386), .C (n_6403), .Y (n_6411));
OAI33X1 g60859(.A0 (n_3376), .A1 (n_1537), .A2 (n_6390), .B0(n_6409), .B1 (n_6402), .B2 (n_6406), .Y (n_6410));
NAND3X1 g60863(.A (n_6407), .B (n_6404), .C (n_2019), .Y (n_6408));
NAND4X1 g60864(.A (n_6407), .B (n_6406), .C (n_1321), .D (n_6398), .Y(n_6413));
NAND4X1 g60865(.A (n_6393), .B (n_1543), .C (n_1321), .D (n_6404), .Y(n_6405));
OR4X1 g60866(.A (n_6390), .B (n_6402), .C (n_6400), .D (n_6399), .Y(n_6403));
OAI21X1 g60862(.A0 (n_6388), .A1 (n_6400), .B0 (n_6389), .Y (n_6401));
NAND4X1 g60867(.A (n_6396), .B (n_6399), .C (n_6395), .D (n_6398), .Y(n_6409));
NAND4X1 g60868(.A (n_6396), .B (n_1212), .C (n_6395), .D (n_6406), .Y(n_6397));
AND2X1 g60869(.A (n_6394), .B (n_6392), .Y (n_6407));
AND2X1 g60871(.A (n_1213), .B (n_6392), .Y (n_6393));
INVX1 g60875(.A (n_6396), .Y (n_6390));
NAND4X1 g60872(.A (n_6388), .B (n_6404), .C (n_4878), .D (n_1321), .Y(n_6389));
AND2X1 g60873(.A (n_6388), .B (n_1055), .Y (n_6392));
AND2X1 g60876(.A (n_6388), .B (n_3641), .Y (n_6396));
NAND4X1 g60870(.A (n_6388), .B (n_1536), .C (n_6399), .D (n_3211), .Y(n_6386));
OAI21X1 g60877(.A0 (g4420), .A1 (g4427), .B0 (g35), .Y (n_6388));
DFFSRX1 g4420_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6385), .Q (g4420), .QN ());
MX2X1 g60879(.A (g4534), .B (n_6384), .S0 (n_10005), .Y (n_6385));
XOR2X1 g60880(.A (g4534), .B (g10306), .Y (n_6384));
DFFSRX1 g4534_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6383), .Q (g4534), .QN ());
OAI21X1 g60882(.A0 (n_6379), .A1 (n_9627), .B0 (n_6382), .Y (n_6383));
OAI21X1 g60883(.A0 (n_6381), .A1 (g2988), .B0 (n_9091), .Y (n_6382));
INVX1 g60884(.A (n_6380), .Y (n_6381));
NAND4X1 g60885(.A (g4564), .B (g4555), .C (g4561), .D (g4558), .Y(n_6380));
INVX1 g60886(.A (g4564), .Y (n_6379));
DFFSRX1 g4564_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6378), .Q (g4564), .QN ());
NAND2X1 g60888(.A (n_6377), .B (n_3113), .Y (n_6378));
NAND2X1 g60889(.A (g4561), .B (n_10078), .Y (n_6377));
DFFSRX1 g4561_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6376), .Q (g4561), .QN ());
NAND2X1 g60891(.A (n_6375), .B (n_3115), .Y (n_6376));
NAND2X1 g60892(.A (g4558), .B (n_10078), .Y (n_6375));
DFFSRX1 g4558_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6373), .Q (g4558), .QN ());
NAND2X1 g60896(.A (n_6372), .B (n_3117), .Y (n_6373));
NAND2X1 g60898(.A (g4555), .B (n_10078), .Y (n_6372));
DFFSRX1 g4555_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(gbuf3), .Q (g4555), .QN ());
DFFSRX1 g4571_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g4570), .Q (gbuf3), .QN ());
DFFSRX1 g74_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6370), .Q (g20763), .QN ());
DFFSRX1 g4570_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6371), .Q (g4570), .QN ());
DFFSRX1 g355_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6369), .Q (g_12276), .QN ());
OAI21X1 g60911(.A0 (n_6364), .A1 (g4552), .B0 (n_6060), .Y (n_6371));
MX2X1 g60962(.A (g_12276), .B (n_6367), .S0 (n_8955), .Y (n_6370));
OAI21X1 g60984(.A0 (g_21792), .A1 (n_9422), .B0 (n_6368), .Y(n_6369));
DFFSRX1 g4552_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6365), .Q (), .QN (g4552));
NAND3X1 g61012(.A (n_6366), .B (g_21792), .C (n_9681), .Y (n_6368));
MX2X1 g61019(.A (n_6366), .B (g20763), .S0 (g_21792), .Y (n_6367));
OAI21X1 g60929(.A0 (g4549), .A1 (n_6364), .B0 (n_6055), .Y (n_6365));
DFFSRX1 g351_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6363), .Q (), .QN (g_21792));
DFFSRX1 g4512_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6362), .Q (), .QN (g4512));
MX2X1 g61142(.A (n_6359), .B (n_9772), .S0 (g_8657), .Y (n_6363));
DFFSRX1 g4549_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6361), .Q (), .QN (g4549));
DFFSRX1 g4300_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6360), .Q (g4300), .QN ());
OAI21X1 g60944(.A0 (g4504), .A1 (n_6364), .B0 (n_5821), .Y (n_6362));
OAI21X1 g60986(.A0 (g4546), .A1 (n_6364), .B0 (n_6320), .Y (n_6361));
MX2X1 g61143(.A (g4297), .B (n_6357), .S0 (n_9750), .Y (n_6360));
DFFSRX1 g554_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6508), .Q (g_9338), .QN ());
AND2X1 g61205(.A (n_9553), .B (g7540), .Y (n_6359));
DFFSRX1 g347_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7540), .Q (g_8657), .QN ());
DFFSRX1 g4504_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6356), .Q (), .QN (g4504));
DFFSRX1 g807_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6355), .Q (g_10233), .QN ());
DFFSRX1 g4546_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6351), .Q (), .QN (g4546));
OR2X1 g61211(.A (g4242), .B (g4300), .Y (n_6357));
DFFSRX1 g344_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6348), .Q (g7540), .QN ());
DFFSRX1 g194_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6353), .Q (g8358), .QN ());
DFFSRX1 g2902_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6352), .Q (g2902), .QN ());
OAI21X1 g61017(.A0 (g4501), .A1 (n_6334), .B0 (n_6299), .Y (n_6356));
DFFSRX1 g794_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6347), .Q (), .QN (g_5342));
NAND2X1 g61308(.A (n_6345), .B (n_6346), .Y (n_6355));
MX2X1 g61137(.A (g_10092), .B (n_2648), .S0 (n_9000), .Y (n_6353));
MX2X1 g61168(.A (g2970), .B (n_6336), .S0 (n_9359), .Y (n_6352));
DFFSRX1 g4242_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6342), .Q (g4242), .QN ());
OAI21X1 g61078(.A0 (g4567), .A1 (n_6364), .B0 (n_6297), .Y (n_6351));
OAI22X1 g61330(.A0 (g_8657), .A1 (n_9269), .B0 (g_12275), .B1(n_9830), .Y (n_6348));
NAND2X1 g61367(.A (n_6338), .B (n_6332), .Y (n_6347));
NAND2X1 g61368(.A (g_12275), .B (n_30), .Y (n_6366));
NAND3X1 g61384(.A (n_2221), .B (n_6454), .C (n_10310), .Y (n_6346));
DFFSRX1 g534_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6337), .Q (g_15801), .QN ());
DFFSRX1 g790_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6339), .Q (), .QN (g_20909));
AOI22X1 g61383(.A0 (n_2554), .A1 (n_10306), .B0 (n_6331), .B1(n_9526), .Y (n_6345));
DFFSRX1 g4501_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6335), .Q (), .QN (g4501));
OAI22X1 g61329(.A0 (n_6330), .A1 (n_9599), .B0 (g4235), .B1 (n_9862),.Y (n_6342));
DFFSRX1 g333_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6323), .Q (), .QN (g_12275));
NAND2X1 g61400(.A (n_6317), .B (n_6326), .Y (n_6339));
DFFSRX1 g4567_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6321), .Q (), .QN (g4567));
AOI21X1 g61432(.A0 (n_6324), .A1 (n_9856), .B0 (n_6328), .Y (n_6338));
DFFSRX1 g222_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10715), .Q (g_10092), .QN ());
MX2X1 g61224(.A (g_19459), .B (n_6316), .S0 (n_9834), .Y (n_6337));
NAND3X1 g61259(.A (n_6318), .B (n_11055), .C (n_3765), .Y (n_6336));
DFFSRX1 g785_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6327), .Q (), .QN (g_17086));
OAI21X1 g61131(.A0 (g4498), .A1 (n_6334), .B0 (n_6254), .Y (n_6335));
NAND4X1 g61431(.A (n_10315), .B (n_10310), .C (n_9651), .D (n_6331),.Y (n_6332));
XOR2X1 g61434(.A (n_4247), .B (n_6310), .Y (n_6330));
NOR2X1 g61465(.A (n_1865), .B (n_10315), .Y (n_6328));
NAND2X1 g61475(.A (n_6312), .B (n_6309), .Y (n_6327));
NAND3X1 g61477(.A (n_7395), .B (n_6468), .C (n_6324), .Y (n_6326));
OAI22X1 g61483(.A0 (n_6306), .A1 (n_9193), .B0 (g_18980), .B1(n_9698), .Y (n_6323));
OAI21X1 g61221(.A0 (g4543), .A1 (n_6364), .B0 (n_6320), .Y (n_6321));
DFFSRX1 g781_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6313), .Q (g_16464), .QN ());
NOR2X1 g61306(.A (n_6315), .B (n_6958), .Y (n_6318));
AOI22X1 g61481(.A0 (n_2311), .A1 (n_6621), .B0 (n_6308), .B1(n_9697), .Y (n_6317));
DFFSRX1 g160_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6311), .Q (), .QN (g_16769));
NAND2X1 g61305(.A (g_19913), .B (n_32), .Y (n_6316));
INVX1 g61363(.A (g_19913), .Y (n_6315));
NAND2X1 g61497(.A (n_6290), .B (n_6302), .Y (n_6313));
AOI21X1 g61518(.A0 (g_16464), .A1 (n_9019), .B0 (n_6305), .Y(n_6312));
DFFSRX1 g4498_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6300), .Q (), .QN (g4498));
DFFSRX1 g776_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6303), .Q (g_21799), .QN ());
DFFSRX1 g106_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6301), .Q (g21176), .QN ());
DFFSRX1 g301_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6295), .Q (), .QN (g_19913));
NAND2X2 g61373(.A (n_6285), .B (n_6296), .Y (n_6311));
NAND2X1 g61504(.A (n_6258), .B (n_6288), .Y (n_6310));
NAND3X1 g61512(.A (n_7402), .B (n_6304), .C (n_6308), .Y (n_6309));
AOI21X1 g61547(.A0 (n_6208), .A1 (n_6280), .B0 (n_6286), .Y (n_6306));
DFFSRX1 g3106_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_8605), .Q (), .QN (g3106));
DFFSRX1 g3457_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_7133), .Q (), .QN (g3457));
DFFSRX1 g3808_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6878), .Q (), .QN (g3808));
DFFSRX1 g2799_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6287), .Q (g2799), .QN ());
DFFSRX1 g4543_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6298), .Q (), .QN (g4543));
NOR3X1 g61536(.A (n_6304), .B (n_6308), .C (n_10078), .Y (n_6305));
NAND2X1 g61544(.A (n_6282), .B (n_6271), .Y (n_6303));
NAND3X1 g61546(.A (n_7395), .B (n_8819), .C (g_16464), .Y (n_6302));
OAI21X1 g61587(.A0 (n_9501), .A1 (n_101), .B0 (n_6281), .Y (n_6301));
OAI21X1 g61261(.A0 (g4495), .A1 (n_6334), .B0 (n_6299), .Y (n_6300));
DFFSRX1 g772_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6283), .Q (g_15879), .QN ());
OAI21X1 g61382(.A0 (g4540), .A1 (n_6364), .B0 (n_6297), .Y (n_6298));
NAND3X1 g61401(.A (n_6274), .B (n_2290), .C (n_9398), .Y (n_6296));
AOI21X1 g61402(.A0 (n_6264), .A1 (n_10005), .B0 (g_16769), .Y(n_6295));
AOI22X1 g61549(.A0 (n_2248), .A1 (n_11138), .B0 (g_21799), .B1(n_9193), .Y (n_6290));
OR4X1 g61552(.A (n_6267), .B (g8917), .C (g8915), .D (g8916), .Y(n_6288));
OAI21X1 g61567(.A0 (n_5610), .A1 (n_5761), .B0 (n_6266), .Y (n_6287));
NAND2X1 g61573(.A (n_5520), .B (n_6265), .Y (n_6286));
DFFSRX1 g157_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6275), .Q (), .QN (g_18590));
DFFSRX1 g732_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6279), .Q (g_18793), .QN ());
AOI22X1 g61427(.A0 (n_2291), .A1 (n_6798), .B0 (n_6252), .B1(n_9193), .Y (n_6285));
INVX1 g61569(.A (n_6620), .Y (n_6304));
NAND2X1 g61574(.A (n_6240), .B (n_6259), .Y (n_6283));
AOI21X1 g61591(.A0 (g_15879), .A1 (n_9431), .B0 (n_6262), .Y(n_6282));
OR4X1 g61649(.A (n_6280), .B (g_6192), .C (n_9599), .D (g_18980), .Y(n_6281));
DFFSRX1 g767_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6260), .Q (g_10903), .QN ());
DFFSRX1 g4495_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6255), .Q (), .QN (g4495));
NAND3X1 g61449(.A (n_4252), .B (n_6218), .C (n_4025), .Y (n_6279));
NAND2X1 g61468(.A (n_6220), .B (n_6253), .Y (n_6275));
NOR2X1 g61471(.A (n_6153), .B (n_6798), .Y (n_6274));
NAND3X1 g61585(.A (n_7395), .B (n_8821), .C (g_21799), .Y (n_6271));
OR2X1 g61642(.A (n_6239), .B (n_6093), .Y (n_6267));
AOI22X1 g61645(.A0 (g2799), .A1 (n_5675), .B0 (n_9599), .B1 (g20654),.Y (n_6266));
NAND4X1 g61648(.A (g_19187), .B (g_18980), .C (g_16983), .D (n_3519),.Y (n_6265));
DFFSRX1 g142_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6257), .Q (), .QN (g_22605));
DFFSRX1 g3333_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6247), .Q (), .QN (g3333));
DFFSRX1 g3684_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6246), .Q (), .QN (g3684));
DFFSRX1 g4035_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6241), .Q (), .QN (g4035));
DFFSRX1 g1768_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6256), .Q (), .QN (g1768));
DFFSRX1 g4540_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6221), .Q (), .QN (g4540));
INVX1 g61506(.A (n_6798), .Y (n_6264));
NOR3X1 g61627(.A (n_8821), .B (g_21799), .C (n_9772), .Y (n_6262));
NAND2X1 g61639(.A (n_6214), .B (n_6149), .Y (n_6260));
NAND3X1 g61641(.A (n_7402), .B (n_8820), .C (g_15879), .Y (n_6259));
XOR2X1 g61651(.A (g8870), .B (g4235), .Y (n_6258));
DFFSRX1 g4483_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(gbuf1), .Q (g4483), .QN ());
DFFSRX1 g1570_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6217), .Q (g12923), .QN ());
DFFSRX1 g2661_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6235), .Q (), .QN (g2661));
DFFSRX1 g2685_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6234), .Q (g2685), .QN ());
DFFSRX1 g1724_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6232), .Q (g1724), .QN ());
DFFSRX1 g1830_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6230), .Q (g1830), .QN ());
DFFSRX1 g1902_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6238), .Q (), .QN (g1902));
DFFSRX1 g1964_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6229), .Q (g1964), .QN ());
DFFSRX1 g2102_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6228), .Q (), .QN (g2102));
DFFSRX1 g2126_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6226), .Q (g2126), .QN ());
DFFSRX1 g2259_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6225), .Q (), .QN (g2259));
DFFSRX1 g2283_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6224), .Q (g2283), .QN ());
DFFSRX1 g2327_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6237), .Q (), .QN (g2327));
DFFSRX1 g2389_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6223), .Q (g2389), .QN ());
DFFSRX1 g1700_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6233), .Q (), .QN (g1700));
DFFSRX1 g2523_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6222), .Q (g2523), .QN ());
DFFSRX1 g2461_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6236), .Q (), .QN (g2461));
NAND2X2 g61375(.A (n_6091), .B (n_6927), .Y (n_6257));
NAND3X1 g61922(.A (n_6156), .B (n_2551), .C (n_6066), .Y (n_6256));
OAI21X1 g61405(.A0 (g4480), .A1 (n_6364), .B0 (n_6254), .Y (n_6255));
NAND3X1 g61505(.A (n_6154), .B (n_6252), .C (n_9425), .Y (n_6253));
MX2X1 g61519(.A (g3263), .B (n_6100), .S0 (n_9218), .Y (n_6247));
MX2X1 g61520(.A (g3614), .B (n_6098), .S0 (n_9000), .Y (n_6246));
MX2X1 g61556(.A (g3965), .B (n_6096), .S0 (n_9000), .Y (n_6241));
AOI22X1 g61647(.A0 (n_2250), .A1 (n_6211), .B0 (g_10903), .B1(n_9491), .Y (n_6240));
DFFSRX1 g153_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6155), .Q (), .QN (g_9176));
DFFSRX1 g763_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6150), .Q (g_18112), .QN ());
DFFSRX1 g2657_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6206), .Q (g2657), .QN ());
DFFSRX1 g2681_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6203), .Q (), .QN (g2681));
DFFSRX1 g1696_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6204), .Q (g1696), .QN ());
DFFSRX1 g1720_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6202), .Q (), .QN (g1720));
DFFSRX1 g1760_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6201), .Q (g1760), .QN ());
DFFSRX1 g1834_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6199), .Q (), .QN (g1834));
DFFSRX1 g1858_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6198), .Q (g1858), .QN ());
DFFSRX1 g1894_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6197), .Q (g1894), .QN ());
DFFSRX1 g1968_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6194), .Q (), .QN (g1968));
DFFSRX1 g2028_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6176), .Q (g2028), .QN ());
DFFSRX1 g2098_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6190), .Q (g2098), .QN ());
DFFSRX1 g1992_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6192), .Q (g1992), .QN ());
DFFSRX1 g2122_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6189), .Q (), .QN (g2122));
DFFSRX1 g2185_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6174), .Q (g2185), .QN ());
DFFSRX1 g2193_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6210), .Q (), .QN (g2193));
DFFSRX1 g2255_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6188), .Q (g2255), .QN ());
DFFSRX1 g2279_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6186), .Q (), .QN (g2279));
DFFSRX1 g2319_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6185), .Q (g2319), .QN ());
DFFSRX1 g2393_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6184), .Q (), .QN (g2393));
DFFSRX1 g2417_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6183), .Q (g2417), .QN ());
DFFSRX1 g2453_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6182), .Q (g2453), .QN ());
DFFSRX1 g2527_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6180), .Q (), .QN (g2527));
DFFSRX1 g2551_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6178), .Q (g2551), .QN ());
DFFSRX1 g1624_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6171), .Q (g1624), .QN ());
DFFSRX1 g1632_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6209), .Q (), .QN (g1632));
DFFSRX1 g2587_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6169), .Q (g2587), .QN ());
DFFSRX1 g1783_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6165), .Q (n_5996), .QN ());
DFFSRX1 g1792_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6166), .Q (g1792), .QN ());
DFFSRX1 g1811_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6164), .Q (g1811), .QN ());
DFFSRX1 g1917_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6162), .Q (n_5925), .QN ());
DFFSRX1 g2036_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6168), .Q (), .QN (g2036));
DFFSRX1 g2342_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6161), .Q (n_5917), .QN ());
DFFSRX1 g2476_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6160), .Q (n_5921), .QN ());
DFFSRX1 g2595_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6167), .Q (), .QN (g2595));
DFFSRX1 g1825_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6157), .Q (), .QN (g1825));
NAND2X1 g61732(.A (n_6207), .B (g4235), .Y (n_6239));
NAND3X1 g61802(.A (n_6065), .B (n_2307), .C (n_6092), .Y (n_6238));
NAND3X1 g61811(.A (n_6064), .B (n_2294), .C (n_6087), .Y (n_6237));
NAND3X1 g61818(.A (n_6062), .B (n_2781), .C (n_6086), .Y (n_6236));
MX2X1 g61845(.A (g2657), .B (n_6078), .S0 (n_8955), .Y (n_6235));
OAI22X1 g61848(.A0 (n_6082), .A1 (n_9976), .B0 (g2681), .B1 (n_9992),.Y (n_6234));
MX2X1 g61849(.A (g1696), .B (n_6070), .S0 (n_9172), .Y (n_6233));
OAI22X1 g61850(.A0 (n_6080), .A1 (n_9976), .B0 (g1720), .B1 (n_9992),.Y (n_6232));
MX2X1 g61853(.A (n_827), .B (n_6074), .S0 (n_8955), .Y (n_6230));
MX2X1 g61858(.A (n_836), .B (n_6073), .S0 (n_9240), .Y (n_6229));
MX2X1 g61863(.A (g2098), .B (n_6076), .S0 (n_9240), .Y (n_6228));
OAI22X1 g61865(.A0 (n_6081), .A1 (n_9269), .B0 (g2122), .B1 (n_9209),.Y (n_6226));
MX2X1 g61867(.A (g2255), .B (n_6068), .S0 (n_9750), .Y (n_6225));
OAI22X1 g61869(.A0 (n_6079), .A1 (n_9193), .B0 (g2279), .B1 (n_9830),.Y (n_6224));
MX2X1 g61871(.A (n_831), .B (n_6072), .S0 (n_9256), .Y (n_6223));
MX2X1 g61877(.A (n_839), .B (n_6071), .S0 (n_9359), .Y (n_6222));
NAND3X1 g61514(.A (n_6320), .B (n_3996), .C (n_6011), .Y (n_6221));
AOI22X1 g61516(.A0 (n_2308), .A1 (n_6562), .B0 (n_6057), .B1(n_9193), .Y (n_6220));
OR2X1 g61535(.A (n_6216), .B (n_10687), .Y (n_6218));
OAI21X1 g61551(.A0 (n_392), .A1 (n_9425), .B0 (n_6216), .Y (n_6217));
DFFSRX1 g1854_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6142), .Q (), .QN (g1854));
DFFSRX1 g758_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6143), .Q (g_13871), .QN ());
DFFSRX1 g1988_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6141), .Q (), .QN (g1988));
DFFSRX1 g2413_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6140), .Q (), .QN (g2413));
DFFSRX1 g2547_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6138), .Q (), .QN (g2547));
DFFSRX1 g1926_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6133), .Q (g1926), .QN ());
DFFSRX1 g1945_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6132), .Q (g1945), .QN ());
DFFSRX1 g117_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6134), .Q (g21270), .QN ());
DFFSRX1 g2051_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6130), .Q (n_5932), .QN ());
DFFSRX1 g2208_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6126), .Q (n_5941), .QN ());
DFFSRX1 g2217_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6125), .Q (g2217), .QN ());
DFFSRX1 g2236_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6123), .Q (g2236), .QN ());
DFFSRX1 g2060_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6129), .Q (g2060), .QN ());
DFFSRX1 g2351_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6121), .Q (g2351), .QN ());
DFFSRX1 g2370_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6120), .Q (g2370), .QN ());
DFFSRX1 g2079_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6128), .Q (g2079), .QN ());
DFFSRX1 g2485_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6118), .Q (g2485), .QN ());
DFFSRX1 g2504_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6117), .Q (g2504), .QN ());
DFFSRX1 g1648_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6116), .Q (n_5936), .QN ());
DFFSRX1 g1657_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6114), .Q (g1657), .QN ());
DFFSRX1 g2610_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6112), .Q (n_5928), .QN ());
DFFSRX1 g2619_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6110), .Q (g2619), .QN ());
DFFSRX1 g2638_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6109), .Q (g2638), .QN ());
DFFSRX1 g1677_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6111), .Q (g1677), .QN ());
DFFSRX1 g2652_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6101), .Q (g2652), .QN ());
DFFSRX1 g1691_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6108), .Q (g1691), .QN ());
DFFSRX1 g1959_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6107), .Q (), .QN (g1959));
DFFSRX1 g2093_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6102), .Q (g2093), .QN ());
DFFSRX1 g2250_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6105), .Q (g2250), .QN ());
DFFSRX1 g2384_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6104), .Q (), .QN (g2384));
DFFSRX1 g2518_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6103), .Q (), .QN (g2518));
DFFSRX1 g4520_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g4519), .Q (gbuf1), .QN ());
AOI21X1 g61743(.A0 (g_18112), .A1 (n_9419), .B0 (n_6146), .Y(n_6214));
DFFSRX1 g121_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6136), .Q (g20654), .QN ());
DFFSRX1 g329_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6137), .Q (), .QN (g_18980));
NAND3X1 g61808(.A (n_6010), .B (n_2259), .C (n_6044), .Y (n_6210));
NAND3X1 g61820(.A (n_6009), .B (n_2522), .C (n_6043), .Y (n_6209));
OAI21X1 g61832(.A0 (g_19304), .A1 (g_16983), .B0 (g_19187), .Y(n_6208));
NOR2X1 g61835(.A (g11770), .B (g8920), .Y (n_6207));
MX2X1 g61844(.A (g2652), .B (n_6024), .S0 (n_9311), .Y (n_6206));
MX2X1 g61846(.A (g1691), .B (n_6030), .S0 (n_9156), .Y (n_6204));
MX2X1 g61847(.A (n_6020), .B (n_6021), .S0 (n_9172), .Y (n_6203));
MX2X1 g61851(.A (n_6027), .B (n_6028), .S0 (n_9000), .Y (n_6202));
OAI22X1 g61852(.A0 (n_6042), .A1 (n_9269), .B0 (g1768), .B1 (n_9627),.Y (n_6201));
MX2X1 g61854(.A (g1830), .B (n_6016), .S0 (n_9234), .Y (n_6199));
OAI22X1 g61855(.A0 (n_6038), .A1 (n_10952), .B0 (g1854), .B1(n_9311), .Y (n_6198));
OAI22X1 g61857(.A0 (n_6041), .A1 (n_9599), .B0 (g1902), .B1(n_10063), .Y (n_6197));
MX2X1 g61859(.A (g1964), .B (n_6015), .S0 (n_9834), .Y (n_6194));
OAI22X1 g61861(.A0 (n_6037), .A1 (n_9976), .B0 (g1988), .B1 (n_9862),.Y (n_6192));
MX2X1 g61862(.A (g2093), .B (n_6019), .S0 (n_9172), .Y (n_6190));
MX2X1 g61864(.A (n_6017), .B (n_6018), .S0 (n_9091), .Y (n_6189));
MX2X1 g61866(.A (g2250), .B (n_6029), .S0 (n_9256), .Y (n_6188));
MX2X1 g61868(.A (n_6025), .B (n_6026), .S0 (n_9000), .Y (n_6186));
OAI22X1 g61870(.A0 (n_6040), .A1 (n_9884), .B0 (g2327), .B1 (n_9830),.Y (n_6185));
MX2X1 g61872(.A (g2389), .B (n_6014), .S0 (n_9156), .Y (n_6184));
OAI22X1 g61874(.A0 (n_6034), .A1 (n_9461), .B0 (g2413), .B1(n_10063), .Y (n_6183));
OAI22X1 g61875(.A0 (n_6039), .A1 (n_9772), .B0 (g2461), .B1(n_10005), .Y (n_6182));
MX2X1 g61878(.A (g2523), .B (n_6013), .S0 (n_9797), .Y (n_6180));
OAI22X1 g61880(.A0 (n_6033), .A1 (n_9431), .B0 (g2547), .B1 (n_9811),.Y (n_6178));
OAI22X1 g61881(.A0 (n_6036), .A1 (n_9976), .B0 (g2036), .B1 (n_9627),.Y (n_6176));
OAI22X1 g61882(.A0 (n_6035), .A1 (n_9976), .B0 (g2193), .B1 (n_9651),.Y (n_6174));
OAI22X1 g61883(.A0 (n_6032), .A1 (n_9772), .B0 (g1632), .B1 (n_9862),.Y (n_6171));
OAI22X1 g61884(.A0 (n_6031), .A1 (n_9772), .B0 (g2595), .B1 (n_9811),.Y (n_6169));
NAND3X1 g61924(.A (n_6089), .B (n_2795), .C (n_5956), .Y (n_6168));
NAND3X1 g61936(.A (n_6084), .B (n_2254), .C (n_5951), .Y (n_6167));
MX2X1 g61973(.A (g1798), .B (n_5997), .S0 (n_9894), .Y (n_6166));
MX2X1 g61974(.A (g1760), .B (n_5999), .S0 (n_9469), .Y (n_6165));
MX2X1 g61975(.A (g1792), .B (n_6000), .S0 (n_9425), .Y (n_6164));
MX2X1 g61976(.A (g1894), .B (n_6002), .S0 (n_9091), .Y (n_6162));
MX2X1 g61986(.A (g2319), .B (n_5995), .S0 (n_9469), .Y (n_6161));
MX2X1 g61989(.A (g2453), .B (n_6001), .S0 (n_9091), .Y (n_6160));
OAI21X1 g62028(.A0 (n_2464), .A1 (n_5849), .B0 (n_6061), .Y (n_6157));
NAND3X1 g62054(.A (n_3948), .B (n_5993), .C (n_9501), .Y (n_6156));
NAND2X1 g61541(.A (n_6003), .B (n_6058), .Y (n_6155));
NOR2X1 g61542(.A (n_6153), .B (n_6562), .Y (n_6154));
DFFSRX1 g4527_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6050), .Q (g4527), .QN ());
NAND2X1 g61720(.A (n_6094), .B (n_6048), .Y (n_6150));
NAND3X1 g61731(.A (n_7395), .B (n_6145), .C (g_10903), .Y (n_6149));
DFFSRX1 g4235_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8920), .Q (), .QN (g4235));
INVX1 g61798(.A (n_8820), .Y (n_6211));
NOR3X1 g61803(.A (n_6145), .B (g_10903), .C (n_9772), .Y (n_6146));
NAND2X1 g61824(.A (n_6045), .B (n_5988), .Y (n_6143));
MX2X1 g61856(.A (n_5978), .B (n_5979), .S0 (n_8955), .Y (n_6142));
MX2X1 g61860(.A (n_5975), .B (n_5976), .S0 (n_8955), .Y (n_6141));
MX2X1 g61873(.A (n_5972), .B (n_5973), .S0 (n_9091), .Y (n_6140));
MX2X1 g61879(.A (n_5969), .B (n_5970), .S0 (n_9000), .Y (n_6138));
INVX1 g61904(.A (g_19187), .Y (n_6137));
OAI21X1 g61917(.A0 (g23759), .A1 (n_9425), .B0 (n_5795), .Y (n_6136));
OAI21X1 g61932(.A0 (g23652), .A1 (n_9681), .B0 (n_5792), .Y (n_6134));
MX2X1 g61977(.A (g1932), .B (n_5926), .S0 (n_9797), .Y (n_6133));
MX2X1 g61978(.A (g1926), .B (n_5924), .S0 (n_9558), .Y (n_6132));
MX2X1 g61979(.A (g2028), .B (n_5934), .S0 (n_9681), .Y (n_6130));
MX2X1 g61980(.A (g2066), .B (n_5933), .S0 (n_8955), .Y (n_6129));
MX2X1 g61981(.A (g2060), .B (n_5931), .S0 (n_9425), .Y (n_6128));
MX2X1 g61983(.A (g2185), .B (n_5943), .S0 (n_9558), .Y (n_6126));
MX2X1 g61984(.A (g2223), .B (n_5942), .S0 (n_9234), .Y (n_6125));
MX2X1 g61985(.A (g2217), .B (n_5940), .S0 (n_9139), .Y (n_6123));
MX2X1 g61987(.A (g2357), .B (n_5918), .S0 (n_8955), .Y (n_6121));
MX2X1 g61988(.A (g2351), .B (n_5916), .S0 (n_9558), .Y (n_6120));
MX2X1 g61990(.A (g2491), .B (n_5922), .S0 (n_9091), .Y (n_6118));
MX2X1 g61991(.A (g2485), .B (n_5920), .S0 (n_9558), .Y (n_6117));
MX2X1 g61992(.A (g1624), .B (n_5939), .S0 (n_9558), .Y (n_6116));
MX2X1 g61993(.A (g1664), .B (n_5937), .S0 (n_9091), .Y (n_6114));
MX2X1 g61994(.A (g2587), .B (n_5930), .S0 (n_10063), .Y (n_6112));
MX2X1 g61995(.A (g1657), .B (n_5935), .S0 (n_9558), .Y (n_6111));
MX2X1 g61996(.A (g2625), .B (n_5929), .S0 (n_9992), .Y (n_6110));
MX2X1 g61997(.A (g2619), .B (n_5927), .S0 (n_10063), .Y (n_6109));
NAND3X1 g62022(.A (n_5875), .B (n_2523), .C (n_5904), .Y (n_6108));
OAI21X1 g62033(.A0 (n_2463), .A1 (n_5839), .B0 (n_6008), .Y (n_6107));
NAND3X1 g62038(.A (n_5948), .B (n_2537), .C (n_5899), .Y (n_6105));
OAI21X1 g62042(.A0 (n_2461), .A1 (n_5844), .B0 (n_6006), .Y (n_6104));
OAI21X1 g62046(.A0 (n_2460), .A1 (n_5833), .B0 (n_6004), .Y (n_6103));
NAND3X1 g62049(.A (n_5950), .B (n_2419), .C (n_5901), .Y (n_6102));
NAND3X1 g62051(.A (n_5945), .B (n_2524), .C (n_5896), .Y (n_6101));
DFFSRX1 g4480_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6012), .Q (), .QN (g4480));
NOR2X1 g61539(.A (n_6059), .B (n_6005), .Y (n_6320));
NOR2X1 g61540(.A (n_6054), .B (n_6334), .Y (n_6297));
NAND2X1 g61581(.A (g_19492), .B (n_9894), .Y (n_6216));
OAI21X1 g61593(.A0 (n_3775), .A1 (n_7235), .B0 (n_3603), .Y (n_6100));
OAI21X1 g61594(.A0 (n_3779), .A1 (n_8908), .B0 (n_3599), .Y (n_6098));
OAI21X1 g61650(.A0 (n_6243), .A1 (n_6095), .B0 (n_3593), .Y (n_6096));
DFFSRX1 g4515_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5994), .Q (g4515), .QN ());
DFFSRX1 g749_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6046), .Q (n_8793), .QN ());
DFFSRX1 g4519_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5991), .Q (g4519), .QN ());
AOI22X1 g61840(.A0 (n_2546), .A1 (n_6457), .B0 (g_13871), .B1(n_9193), .Y (n_6094));
DFFSRX1 g4232_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8919), .Q (g8920), .QN ());
DFFSRX1 g319_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5986), .Q (), .QN (g_19187));
OR2X1 g61944(.A (n_5984), .B (g8919), .Y (n_6093));
NAND3X1 g62055(.A (n_3945), .B (n_5909), .C (n_9811), .Y (n_6092));
NAND3X1 g61466(.A (n_5981), .B (n_10713), .C (n_10063), .Y (n_6091));
NAND3X1 g62057(.A (n_4318), .B (n_5882), .C (n_9425), .Y (n_6089));
NAND3X1 g62067(.A (n_4124), .B (n_5907), .C (n_9698), .Y (n_6087));
NAND3X1 g62070(.A (n_4122), .B (n_5905), .C (n_9698), .Y (n_6086));
NAND3X1 g62072(.A (n_4118), .B (n_5877), .C (n_9359), .Y (n_6084));
AOI21X1 g62081(.A0 (n_10790), .A1 (g2685), .B0 (n_5957), .Y (n_6082));
AOI21X1 g62087(.A0 (n_10995), .A1 (g2126), .B0 (n_5952), .Y (n_6081));
AOI21X1 g62090(.A0 (n_10617), .A1 (g1724), .B0 (n_10618), .Y(n_6080));
AOI21X1 g62091(.A0 (n_6067), .A1 (g2283), .B0 (n_5960), .Y (n_6079));
OAI21X1 g62106(.A0 (n_5958), .A1 (n_10790), .B0 (n_5959), .Y(n_6078));
OAI21X1 g62109(.A0 (n_5953), .A1 (n_10995), .B0 (n_5954), .Y(n_6076));
MX2X1 g62119(.A (g1830), .B (n_828), .S0 (n_5884), .Y (n_6074));
MX2X1 g62121(.A (g1964), .B (n_837), .S0 (n_5883), .Y (n_6073));
MX2X1 g62125(.A (g2389), .B (n_832), .S0 (n_5880), .Y (n_6072));
MX2X1 g62128(.A (g2523), .B (n_840), .S0 (n_5878), .Y (n_6071));
OAI21X1 g62130(.A0 (n_5964), .A1 (n_10617), .B0 (n_5965), .Y(n_6070));
OAI21X1 g62131(.A0 (n_5961), .A1 (n_6067), .B0 (n_5962), .Y (n_6068));
NAND3X1 g62255(.A (n_5992), .B (n_136), .C (n_9750), .Y (n_6066));
NAND3X1 g62256(.A (n_5910), .B (n_67), .C (n_9139), .Y (n_6065));
NAND3X1 g62264(.A (n_5908), .B (n_57), .C (n_9139), .Y (n_6064));
NAND3X1 g62265(.A (n_5906), .B (n_12), .C (n_10063), .Y (n_6062));
AOI22X1 g62270(.A0 (n_2168), .A1 (n_5849), .B0 (g1811), .B1(n_10376), .Y (n_6061));
INVX1 g61576(.A (n_6059), .Y (n_6060));
NAND3X1 g61580(.A (n_5913), .B (n_6057), .C (n_10063), .Y (n_6058));
INVX1 g61578(.A (n_6054), .Y (n_6055));
NOR2X1 g61622(.A (n_6052), .B (n_8908), .Y (n_6248));
NOR2X1 g61621(.A (n_6051), .B (n_6956), .Y (n_6250));
OAI22X1 g60899(.A0 (n_5869), .A1 (n_9976), .B0 (g4521), .B1 (n_9830),.Y (n_6050));
DFFSRX1 g298_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5982), .Q (), .QN (g_22070));
DFFSRX1 g150_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5914), .Q (g_16311), .QN ());
DFFSRX1 g739_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5983), .Q (g_10556), .QN ());
DFFSRX1 g744_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5985), .Q (g_16296), .QN ());
DFFSRX1 g542_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5967), .Q (g_19459), .QN ());
NOR2X1 g61707(.A (n_6049), .B (n_6095), .Y (n_8883));
NAND3X1 g61833(.A (n_7402), .B (n_6715), .C (g_18112), .Y (n_6048));
INVX1 g61919(.A (n_6716), .Y (n_6145));
NAND2X1 g61923(.A (n_5830), .B (n_5889), .Y (n_6046));
AOI21X1 g61961(.A0 (n_8793), .A1 (n_9141), .B0 (n_5891), .Y (n_6045));
NAND3X1 g62059(.A (n_4109), .B (n_5872), .C (n_9091), .Y (n_6044));
NAND3X1 g62071(.A (n_3938), .B (n_5870), .C (n_9811), .Y (n_6043));
AOI22X1 g62083(.A0 (n_1040), .A1 (n_5788), .B0 (n_5818), .B1 (g1760),.Y (n_6042));
AOI22X1 g62084(.A0 (n_1044), .A1 (n_5784), .B0 (n_5816), .B1 (g1894),.Y (n_6041));
AOI22X1 g62088(.A0 (n_1053), .A1 (n_5786), .B0 (n_5817), .B1 (g2319),.Y (n_6040));
AOI22X1 g62089(.A0 (n_1052), .A1 (n_5782), .B0 (n_5815), .B1 (g2453),.Y (n_6039));
AOI21X1 g62092(.A0 (n_5977), .A1 (g1858), .B0 (n_5888), .Y (n_6038));
AOI21X1 g62093(.A0 (n_5974), .A1 (g1992), .B0 (n_5887), .Y (n_6037));
AOI22X1 g62094(.A0 (n_765), .A1 (n_5949), .B0 (n_5809), .B1 (g2028),.Y (n_6036));
AOI22X1 g62095(.A0 (n_775), .A1 (n_5947), .B0 (n_5806), .B1 (g2185),.Y (n_6035));
AOI21X1 g62096(.A0 (n_5971), .A1 (g2417), .B0 (n_5886), .Y (n_6034));
AOI21X1 g62098(.A0 (n_5968), .A1 (g2551), .B0 (n_5885), .Y (n_6033));
AOI22X1 g62099(.A0 (n_769), .A1 (n_5799), .B0 (n_5801), .B1 (g1624),.Y (n_6032));
AOI22X1 g62100(.A0 (n_782), .A1 (n_5944), .B0 (n_5803), .B1 (g2587),.Y (n_6031));
MX2X1 g62107(.A (n_841), .B (g1696), .S0 (n_5800), .Y (n_6030));
MX2X1 g62110(.A (n_833), .B (g2255), .S0 (n_5797), .Y (n_6029));
MX2X1 g62115(.A (n_6027), .B (n_878), .S0 (n_10617), .Y (n_6028));
MX2X1 g62116(.A (n_6025), .B (n_975), .S0 (n_6067), .Y (n_6026));
MX2X1 g62117(.A (n_829), .B (g2657), .S0 (n_5814), .Y (n_6024));
MX2X1 g62118(.A (n_6020), .B (n_852), .S0 (n_10790), .Y (n_6021));
MX2X1 g62123(.A (n_834), .B (g2098), .S0 (n_5807), .Y (n_6019));
MX2X1 g62124(.A (n_6017), .B (n_860), .S0 (n_10995), .Y (n_6018));
XOR2X1 g62133(.A (n_4948), .B (n_5811), .Y (n_6016));
XOR2X1 g62134(.A (n_4946), .B (n_5810), .Y (n_6015));
XOR2X1 g62135(.A (n_4942), .B (n_5805), .Y (n_6014));
XOR2X1 g62136(.A (n_5229), .B (n_5804), .Y (n_6013));
NAND3X1 g61527(.A (n_6011), .B (n_2356), .C (n_6299), .Y (n_6012));
NAND3X1 g62250(.A (n_5873), .B (n_96), .C (n_9139), .Y (n_6010));
NAND3X1 g62252(.A (n_5871), .B (n_105), .C (n_10063), .Y (n_6009));
AOI22X1 g62271(.A0 (n_2212), .A1 (n_5839), .B0 (g1945), .B1 (n_9193),.Y (n_6008));
AOI22X1 g62275(.A0 (n_2229), .A1 (n_5844), .B0 (g2370), .B1 (n_9404),.Y (n_6006));
AND2X1 g61577(.A (g4575), .B (n_6005), .Y (n_6059));
AOI22X1 g62276(.A0 (n_2230), .A1 (n_5833), .B0 (g2504), .B1 (n_9599),.Y (n_6004));
AND2X1 g61579(.A (g4578), .B (n_6005), .Y (n_6054));
AOI22X1 g61589(.A0 (n_2270), .A1 (n_10261), .B0 (g_16311), .B1(n_10376), .Y (n_6003));
MX2X1 g62310(.A (n_5925), .B (g1894), .S0 (n_5784), .Y (n_6002));
DFFSRX1 g496_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5879), .Q (g_19492), .QN ());
MX2X1 g62313(.A (n_5921), .B (g2453), .S0 (n_5782), .Y (n_6001));
MX2X1 g62316(.A (g1811), .B (n_2975), .S0 (n_5788), .Y (n_6000));
MX2X1 g62317(.A (n_5996), .B (g1760), .S0 (n_5788), .Y (n_5999));
MX2X1 g62318(.A (g1792), .B (n_5996), .S0 (n_5788), .Y (n_5997));
MX2X1 g62319(.A (n_5917), .B (g2319), .S0 (n_5786), .Y (n_5995));
DFFSRX1 g1227_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5874), .Q (g12919), .QN ());
DFFSRX1 g2771_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5868), .Q (g2771), .QN ());
DFFSRX1 g2775_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5866), .Q (g2775), .QN ());
DFFSRX1 g2783_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5865), .Q (g2783), .QN ());
DFFSRX1 g2787_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5863), .Q (g2787), .QN ());
DFFSRX1 g2803_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5862), .Q (g2803), .QN ());
DFFSRX1 g2807_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5860), .Q (g2807), .QN ());
DFFSRX1 g2815_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5859), .Q (g2815), .QN ());
DFFSRX1 g2819_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5857), .Q (g2819), .QN ());
MX2X1 g60900(.A (g4527), .B (n_5813), .S0 (n_9000), .Y (n_5994));
INVX1 g62591(.A (n_5992), .Y (n_5993));
MX2X1 g60909(.A (g4515), .B (n_5837), .S0 (n_8955), .Y (n_5991));
AND2X1 g61806(.A (n_5781), .B (n_5831), .Y (n_6095));
NAND3X1 g61942(.A (n_7395), .B (n_6524), .C (g_13871), .Y (n_5988));
DFFSRX1 g4229_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8918), .Q (g8919), .QN ());
NAND2X1 g62029(.A (n_5822), .B (n_5573), .Y (n_5986));
NAND2X1 g62048(.A (n_5775), .B (n_5824), .Y (n_5985));
OR2X1 g62060(.A (g8918), .B (g8870), .Y (n_5984));
OAI21X1 g62085(.A0 (n_7094), .A1 (n_9797), .B0 (n_5825), .Y (n_5983));
NAND2X1 g61496(.A (n_5779), .B (n_5828), .Y (n_5982));
NOR2X1 g61501(.A (n_5723), .B (n_7144), .Y (n_5981));
MX2X1 g62120(.A (n_5978), .B (n_883), .S0 (n_5977), .Y (n_5979));
MX2X1 g62122(.A (n_5975), .B (n_885), .S0 (n_5974), .Y (n_5976));
MX2X1 g62126(.A (n_5972), .B (n_866), .S0 (n_5971), .Y (n_5973));
MX2X1 g62129(.A (n_5969), .B (n_858), .S0 (n_5968), .Y (n_5970));
DFFSRX1 g2834_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5794), .Q (), .QN (g23652));
DFFSRX1 g2831_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5796), .Q (), .QN (g23759));
OAI21X1 g63520(.A0 (n_35), .A1 (n_9493), .B0 (n_5820), .Y (n_5967));
NAND2X1 g62218(.A (n_5964), .B (n_10617), .Y (n_5965));
NAND2X1 g62220(.A (n_5961), .B (n_6067), .Y (n_5962));
NOR2X1 g62221(.A (n_976), .B (n_6067), .Y (n_5960));
NAND2X1 g62223(.A (n_5958), .B (n_10790), .Y (n_5959));
NOR2X1 g62224(.A (n_10790), .B (n_10554), .Y (n_5957));
NAND3X1 g62231(.A (n_5881), .B (n_54), .C (n_9425), .Y (n_5956));
NAND2X1 g62232(.A (n_5953), .B (n_10995), .Y (n_5954));
NOR2X1 g62233(.A (n_861), .B (n_10995), .Y (n_5952));
NAND3X1 g62249(.A (n_5876), .B (n_52), .C (n_9811), .Y (n_5951));
NAND3X1 g62258(.A (n_2080), .B (n_5949), .C (n_9501), .Y (n_5950));
NAND3X1 g62261(.A (n_2079), .B (n_5947), .C (n_9698), .Y (n_5948));
NAND3X1 g62266(.A (n_2081), .B (n_5944), .C (n_9425), .Y (n_5945));
MX2X1 g62295(.A (n_5941), .B (g2185), .S0 (n_5947), .Y (n_5943));
MX2X1 g62296(.A (g2217), .B (n_5941), .S0 (n_5947), .Y (n_5942));
MX2X1 g62297(.A (g2236), .B (n_2651), .S0 (n_5947), .Y (n_5940));
MX2X1 g62299(.A (n_5936), .B (g1624), .S0 (n_5799), .Y (n_5939));
MX2X1 g62300(.A (g1657), .B (n_5936), .S0 (n_5799), .Y (n_5937));
MX2X1 g62301(.A (g1677), .B (n_2469), .S0 (n_5799), .Y (n_5935));
MX2X1 g62304(.A (n_5932), .B (g2028), .S0 (n_5949), .Y (n_5934));
MX2X1 g62305(.A (g2060), .B (n_5932), .S0 (n_5949), .Y (n_5933));
MX2X1 g62306(.A (g2079), .B (n_2472), .S0 (n_5949), .Y (n_5931));
MX2X1 g62307(.A (n_5928), .B (g2587), .S0 (n_5944), .Y (n_5930));
MX2X1 g62308(.A (g2619), .B (n_5928), .S0 (n_5944), .Y (n_5929));
MX2X1 g62309(.A (g2638), .B (n_2466), .S0 (n_5944), .Y (n_5927));
MX2X1 g62311(.A (g1926), .B (n_5925), .S0 (n_5784), .Y (n_5926));
MX2X1 g62312(.A (g1945), .B (n_2738), .S0 (n_5784), .Y (n_5924));
MX2X1 g62314(.A (g2485), .B (n_5921), .S0 (n_5782), .Y (n_5922));
MX2X1 g62315(.A (g2504), .B (n_2969), .S0 (n_5782), .Y (n_5920));
MX2X1 g62320(.A (g2351), .B (n_5917), .S0 (n_5786), .Y (n_5918));
MX2X1 g62321(.A (g2370), .B (n_2967), .S0 (n_5786), .Y (n_5916));
NAND2X1 g61632(.A (n_5769), .B (n_5819), .Y (n_5914));
NOR2X1 g61633(.A (n_6153), .B (n_10261), .Y (n_5913));
NAND2X1 g62592(.A (n_5788), .B (n_1667), .Y (n_5992));
INVX1 g62596(.A (n_5909), .Y (n_5910));
INVX1 g62619(.A (n_5907), .Y (n_5908));
INVX1 g62626(.A (n_5905), .Y (n_5906));
NAND3X1 g62647(.A (n_10614), .B (g1691), .C (n_9894), .Y (n_5904));
NAND3X1 g62653(.A (n_5854), .B (g2093), .C (n_9894), .Y (n_5901));
NAND3X1 g62655(.A (n_5852), .B (g2250), .C (n_9139), .Y (n_5899));
NAND3X1 g62661(.A (n_10787), .B (g2652), .C (n_9811), .Y (n_5896));
DFFSRX1 g341_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5774), .Q (g_6192), .QN ());
NOR3X1 g62032(.A (n_9461), .B (g_13871), .C (n_6524), .Y (n_5891));
NAND3X1 g62056(.A (n_7395), .B (n_6523), .C (n_8793), .Y (n_5889));
NOR2X1 g62208(.A (n_884), .B (n_5977), .Y (n_5888));
NOR2X1 g62210(.A (n_886), .B (n_5974), .Y (n_5887));
NOR2X1 g62212(.A (n_867), .B (n_5971), .Y (n_5886));
NOR2X1 g62216(.A (n_859), .B (n_5968), .Y (n_5885));
DFFSRX1 g4575_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10388), .Q (g4575), .QN ());
DFFSRX1 g4578_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5772), .Q (g4578), .QN ());
DFFSRX1 g4388_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5777), .Q (g4388), .QN ());
DFFSRX1 g4401_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5776), .Q (g4401), .QN ());
DFFSRX1 g164_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5790), .Q (g_11293), .QN ());
DFFSRX1 g446_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5780), .Q (g_21576), .QN ());
DFFSRX1 g336_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5768), .Q (g_19304), .QN ());
NOR2X1 g62593(.A (n_5849), .B (n_1236), .Y (n_5884));
NOR2X1 g62597(.A (n_5839), .B (n_1063), .Y (n_5909));
NOR2X1 g62602(.A (n_5839), .B (n_1230), .Y (n_5883));
INVX1 g62607(.A (n_5881), .Y (n_5882));
NOR2X1 g62620(.A (n_5844), .B (n_1060), .Y (n_5907));
NOR2X1 g62623(.A (n_5844), .B (n_1160), .Y (n_5880));
NOR2X1 g62627(.A (n_5833), .B (n_1065), .Y (n_5905));
MX2X1 g61746(.A (g20901), .B (g_20208), .S0 (n_9359), .Y (n_5879));
NOR2X1 g62629(.A (n_5833), .B (n_1138), .Y (n_5878));
INVX1 g62634(.A (n_5876), .Y (n_5877));
NAND3X1 g62637(.A (n_5799), .B (n_2099), .C (n_9698), .Y (n_5875));
MX2X1 g61748(.A (g20901), .B (n_8799), .S0 (n_9019), .Y (n_5874));
INVX1 g62639(.A (n_5872), .Y (n_5873));
INVX1 g62642(.A (n_5870), .Y (n_5871));
AOI21X1 g60906(.A0 (n_3493), .A1 (g4521), .B0 (n_5767), .Y (n_5869));
MX2X1 g62694(.A (g2775), .B (n_5737), .S0 (n_9091), .Y (n_5868));
MX2X1 g62695(.A (g2783), .B (n_5736), .S0 (n_9797), .Y (n_5866));
MX2X1 g62696(.A (g2787), .B (n_5735), .S0 (n_9797), .Y (n_5865));
MX2X1 g62697(.A (g2795), .B (n_5734), .S0 (n_9834), .Y (n_5863));
MX2X1 g62699(.A (g2807), .B (n_5733), .S0 (n_9448), .Y (n_5862));
MX2X1 g62700(.A (g2815), .B (n_5731), .S0 (n_9797), .Y (n_5860));
MX2X1 g62701(.A (g2819), .B (n_5729), .S0 (n_9750), .Y (n_5859));
MX2X1 g62702(.A (g2827), .B (n_5727), .S0 (n_9000), .Y (n_5857));
INVX1 g62811(.A (n_5949), .Y (n_5854));
INVX1 g62841(.A (n_5947), .Y (n_5852));
INVX4 g62874(.A (n_5786), .Y (n_5844));
INVX2 g62883(.A (n_5784), .Y (n_5839));
OAI21X1 g60914(.A0 (g4512), .A1 (n_5711), .B0 (n_5756), .Y (n_5837));
INVX2 g62892(.A (n_5782), .Y (n_5833));
NOR2X1 g61937(.A (n_10416), .B (n_5506), .Y (n_5831));
AOI22X1 g62086(.A0 (n_2246), .A1 (n_5709), .B0 (g_16296), .B1(n_9599), .Y (n_5830));
DFFSRX1 g4226_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8870), .Q (g8918), .QN ());
NAND3X1 g61534(.A (n_5724), .B (n_6928), .C (n_9630), .Y (n_5828));
NAND2X1 g62209(.A (n_5508), .B (n_7395), .Y (n_5825));
NAND3X1 g62257(.A (n_7402), .B (n_10861), .C (g_16296), .Y (n_5824));
MX2X1 g62292(.A (g_16983), .B (n_5707), .S0 (n_9871), .Y (n_5822));
AND2X1 g61631(.A (n_5821), .B (n_3900), .Y (n_6254));
AOI21X1 g61643(.A0 (n_5755), .A1 (n_9351), .B0 (n_6005), .Y (n_6299));
DFFSRX1 g4382_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5738), .Q (g4382), .QN ());
DFFSRX1 g4408_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5714), .Q (g7243), .QN ());
DFFSRX1 g4392_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5716), .Q (g4392), .QN ());
DFFSRX1 g1_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5718), .Q (g12832), .QN ());
DFFSRX1 g4414_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5720), .Q (g7257), .QN ());
DFFSRX1 g294_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5725), .Q (g_18308), .QN ());
DFFSRX1 g4961_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5719), .Q (g4961), .QN ());
OAI21X1 g64026(.A0 (g_19459), .A1 (n_11056), .B0 (n_7395), .Y(n_5820));
DFFSRX1 g146_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5740), .Q (g_15691), .QN ());
DFFSRX1 g2767_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5762), .Q (g2767), .QN ());
DFFSRX1 g2779_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5760), .Q (g2779), .QN ());
DFFSRX1 g2791_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5759), .Q (g2791), .QN ());
DFFSRX1 g2795_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5758), .Q (g2795), .QN ());
DFFSRX1 g2811_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5757), .Q (g2811), .QN ());
DFFSRX1 g2823_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5746), .Q (g2823), .QN ());
DFFSRX1 g2827_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5745), .Q (g2827), .QN ());
NAND3X1 g61724(.A (n_5765), .B (g_16311), .C (n_10385), .Y (n_5819));
NAND2X1 g62563(.A (n_5788), .B (g1792), .Y (n_5818));
NAND2X1 g62566(.A (n_5786), .B (g2351), .Y (n_5817));
NAND2X1 g62567(.A (n_5784), .B (g1926), .Y (n_5816));
NAND2X1 g62568(.A (n_5782), .B (g2485), .Y (n_5815));
NAND2X1 g62586(.A (n_5944), .B (n_1522), .Y (n_5814));
MX2X1 g60905(.A (g4515), .B (n_2101), .S0 (g4521), .Y (n_5813));
INVX1 g62594(.A (n_5977), .Y (n_5811));
INVX1 g62603(.A (n_5974), .Y (n_5810));
NAND2X1 g62606(.A (n_5808), .B (g2060), .Y (n_5809));
NAND2X1 g62608(.A (n_5808), .B (n_1515), .Y (n_5881));
NAND2X1 g62610(.A (n_5808), .B (n_1524), .Y (n_5807));
NAND2X1 g62611(.A (n_5798), .B (g2217), .Y (n_5806));
NAND2X1 g62612(.A (n_5798), .B (n_1517), .Y (n_6067));
INVX1 g62624(.A (n_5971), .Y (n_5805));
INVX1 g62630(.A (n_5968), .Y (n_5804));
NAND2X1 g62633(.A (n_5944), .B (g2619), .Y (n_5803));
NAND2X1 g62632(.A (n_5799), .B (g1657), .Y (n_5801));
NAND2X1 g62635(.A (n_5944), .B (n_1506), .Y (n_5876));
NAND2X1 g62638(.A (n_5799), .B (n_1531), .Y (n_5800));
AND2X1 g62640(.A (n_5798), .B (n_1520), .Y (n_5872));
NAND2X1 g62641(.A (n_5798), .B (n_1527), .Y (n_5797));
AND2X1 g62643(.A (n_5799), .B (g25167), .Y (n_5870));
OAI21X1 g62663(.A0 (n_326), .A1 (n_9333), .B0 (n_5795), .Y (n_5796));
OAI21X1 g62664(.A0 (n_317), .A1 (n_9797), .B0 (n_5792), .Y (n_5794));
NAND2X1 g61823(.A (n_5624), .B (n_5700), .Y (n_5790));
CLKBUFX1 g62812(.A (n_5808), .Y (n_5949));
CLKBUFX1 g62842(.A (n_5798), .Y (n_5947));
INVX2 g62867(.A (n_5788), .Y (n_5849));
NOR2X1 g62036(.A (n_5695), .B (n_5284), .Y (n_5781));
MX2X1 g62137(.A (n_5663), .B (n_5639), .S0 (n_9218), .Y (n_5780));
AOI22X1 g61548(.A0 (n_2271), .A1 (n_7146), .B0 (g_18308), .B1(n_9193), .Y (n_5779));
MX2X1 g61026(.A (g4401), .B (n_5645), .S0 (n_9311), .Y (n_5777));
MX2X1 g61027(.A (g4405), .B (n_5644), .S0 (n_8955), .Y (n_5776));
AOI21X1 g62294(.A0 (g_10556), .A1 (n_9141), .B0 (n_5688), .Y(n_5775));
MX2X1 g62323(.A (g_22328), .B (g21176), .S0 (n_9599), .Y (n_5774));
DFFSRX1 g4749_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5693), .Q (g4749), .QN ());
DFFSRX1 g4894_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5690), .Q (g4894), .QN ());
DFFSRX1 g4771_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5692), .Q (g4771), .QN ());
DFFSRX1 g4760_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5689), .Q (g4760), .QN ());
DFFSRX1 g246_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5694), .Q (g_21813), .QN ());
AOI21X1 g61939(.A0 (n_5654), .A1 (n_816), .B0 (n_364), .Y (g33894));
OAI21X1 g61708(.A0 (n_5681), .A1 (n_9422), .B0 (n_10601), .Y(n_5772));
OR2X1 g62595(.A (n_5744), .B (n_561), .Y (n_5977));
AOI22X1 g61740(.A0 (n_2249), .A1 (n_8583), .B0 (g_11293), .B1(n_9772), .Y (n_5769));
OR2X1 g62604(.A (n_5742), .B (n_647), .Y (n_5974));
OR2X1 g62625(.A (n_5743), .B (n_592), .Y (n_5971));
OR2X1 g62631(.A (n_5741), .B (n_487), .Y (n_5968));
OAI22X1 g62676(.A0 (n_5668), .A1 (n_10952), .B0 (g_16983), .B1(n_9830), .Y (n_5768));
NOR2X1 g60908(.A (n_2100), .B (g4521), .Y (n_5767));
NOR2X1 g61810(.A (n_6153), .B (n_8583), .Y (n_5765));
OAI21X1 g62793(.A0 (n_5614), .A1 (n_5761), .B0 (n_5676), .Y (n_5762));
OAI21X1 g62794(.A0 (n_5613), .A1 (n_5761), .B0 (n_5674), .Y (n_5760));
OAI21X1 g62795(.A0 (n_5612), .A1 (n_5761), .B0 (n_5672), .Y (n_5759));
OAI21X1 g62796(.A0 (n_5611), .A1 (n_5761), .B0 (n_5671), .Y (n_5758));
OAI21X1 g62797(.A0 (n_5609), .A1 (n_5761), .B0 (n_5669), .Y (n_5757));
NAND2X1 g62800(.A (n_5667), .B (n_9091), .Y (n_5795));
NAND2X1 g62801(.A (n_5666), .B (n_9091), .Y (n_5792));
INVX1 g61836(.A (n_5755), .Y (n_5756));
INVX1 g62813(.A (n_10994), .Y (n_5808));
INVX4 g62830(.A (n_10787), .Y (n_5944));
INVX2 g62843(.A (n_5749), .Y (n_5798));
INVX4 g62855(.A (n_10614), .Y (n_5799));
OAI21X1 g62859(.A0 (n_5608), .A1 (n_5761), .B0 (n_5564), .Y (n_5746));
OAI21X1 g62860(.A0 (n_5607), .A1 (n_5761), .B0 (n_5563), .Y (n_5745));
INVX2 g62868(.A (n_5744), .Y (n_5788));
INVX2 g62877(.A (n_5743), .Y (n_5786));
INVX2 g62886(.A (n_5742), .Y (n_5784));
INVX2 g62895(.A (n_5741), .Y (n_5782));
DFFSRX1 g225_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5642), .Q (g_19515), .QN ());
DFFSRX1 g102_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5664), .Q (g20901), .QN ());
OAI21X1 g61945(.A0 (g_22605), .A1 (n_10013), .B0 (n_5678), .Y(n_5740));
NAND3X1 g61008(.A (n_5631), .B (n_2269), .C (n_5592), .Y (n_5738));
OAI21X1 g63287(.A0 (g2767), .A1 (n_5732), .B0 (n_5662), .Y (n_5737));
OAI21X1 g63288(.A0 (n_5730), .A1 (g2779), .B0 (n_5661), .Y (n_5736));
OAI21X1 g63289(.A0 (n_5728), .A1 (g2791), .B0 (n_5660), .Y (n_5735));
OAI21X1 g63290(.A0 (n_5726), .A1 (g2795), .B0 (n_5659), .Y (n_5734));
OAI21X1 g63291(.A0 (n_5732), .A1 (g2799), .B0 (n_5658), .Y (n_5733));
OAI21X1 g63292(.A0 (n_5730), .A1 (g2811), .B0 (n_5657), .Y (n_5731));
OAI21X1 g63293(.A0 (n_5728), .A1 (g2823), .B0 (n_5655), .Y (n_5729));
OAI21X1 g63294(.A0 (n_5726), .A1 (g2827), .B0 (n_5656), .Y (n_5727));
NAND2X1 g61571(.A (n_5602), .B (n_5652), .Y (n_5725));
NOR2X1 g61572(.A (n_5723), .B (n_7146), .Y (n_5724));
NAND3X1 g61030(.A (n_5641), .B (n_5273), .C (n_5578), .Y (n_5720));
NAND2X1 g61583(.A (n_3752), .B (n_5650), .Y (n_5719));
OAI21X1 g61031(.A0 (g4455), .A1 (n_9627), .B0 (n_5715), .Y (n_5718));
OAI21X1 g61050(.A0 (n_74), .A1 (n_9681), .B0 (n_5715), .Y (n_5716));
DFFSRX1 g1682_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6858), .Q (), .QN (g1682));
DFFSRX1 g4430_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5677), .Q (g4430), .QN ());
DFFSRX1 g5115_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_8706), .Q (n_3618), .QN ());
DFFSRX1 g6154_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5646), .Q (n_3589), .QN ());
DFFSRX1 g5808_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5686), .Q (n_3611), .QN ());
DFFSRX1 g4434_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5683), .Q (), .QN (g4434));
DFFSRX1 g5084_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5680), .Q (g5084), .QN ());
NAND2X1 g61051(.A (n_5643), .B (n_5637), .Y (n_5714));
AND2X1 g64156(.A (n_10310), .B (n_9874), .Y (n_7402));
DFFSRX1 g4222_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8917), .Q (g8870), .QN ());
OR2X1 g64274(.A (n_172), .B (n_10311), .Y (n_5712));
NAND3X1 g61733(.A (n_5711), .B (g4572), .C (n_10687), .Y (n_5821));
DFFSRX1 g4521_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5629), .Q (), .QN (g4521));
INVX1 g62761(.A (g_22328), .Y (n_5707));
AND2X1 g61837(.A (n_5711), .B (g20049), .Y (n_5755));
NAND2X1 g62845(.A (n_5622), .B (n_5705), .Y (n_5749));
AOI21X1 g62869(.A0 (n_5569), .A1 (n_5704), .B0 (n_5703), .Y (n_5744));
AOI21X1 g62878(.A0 (n_5567), .A1 (n_5704), .B0 (n_5703), .Y (n_5743));
AOI21X1 g62887(.A0 (n_5568), .A1 (n_5702), .B0 (n_5701), .Y (n_5742));
AOI21X1 g62896(.A0 (n_5566), .A1 (n_5702), .B0 (n_5701), .Y (n_5741));
NAND3X1 g61935(.A (n_5619), .B (g_11293), .C (n_9797), .Y (n_5700));
DFFSRX1 g128_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10690), .Q (g21245), .QN ());
NAND4X1 g62286(.A (n_2448), .B (n_2137), .C (n_5543), .D (n_1686), .Y(n_5695));
MX2X1 g62325(.A (g_20208), .B (n_5583), .S0 (n_9359), .Y (n_5694));
NAND2X1 g61634(.A (n_3582), .B (n_5599), .Y (n_5693));
NAND2X1 g61635(.A (n_3580), .B (n_5596), .Y (n_5692));
DFFSRX1 g5462_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10955), .Q (n_3616), .QN ());
DFFSRX1 g6500_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5600), .Q (n_3604), .QN ());
DFFSRX1 g4826_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5593), .Q (), .QN (g4826));
DFFSRX1 g4831_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5627), .Q (), .QN (g4831));
DFFSRX1 g4446_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5625), .Q (g7245), .QN ());
DFFSRX1 g4449_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5626), .Q (g7260), .QN ());
DFFSRX1 g5080_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5615), .Q (g5080), .QN ());
DFFSRX1 g269_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5590), .Q (g_20208), .QN ());
INVX1 g62589(.A (n_6523), .Y (n_5709));
NAND2X1 g61735(.A (n_5633), .B (n_3578), .Y (n_5690));
NAND2X1 g61734(.A (n_5634), .B (n_3581), .Y (n_5689));
NOR3X1 g62613(.A (n_10861), .B (g_16296), .C (n_9353), .Y (n_5688));
NAND3X1 g61801(.A (n_5576), .B (n_2560), .C (n_3613), .Y (n_5686));
DFFSRX1 g316_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5570), .Q (g_22328), .QN ());
DFFSRX1 g4219_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8916), .Q (g8917), .QN ());
MX2X1 g61842(.A (g4452), .B (n_5532), .S0 (n_8955), .Y (n_5683));
INVX1 g61885(.A (g4572), .Y (n_5681));
OAI21X1 g61915(.A0 (n_5515), .A1 (g5080), .B0 (n_5571), .Y (n_5680));
DFFSRX1 g291_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5557), .Q (g_12922), .QN ());
NAND4X1 g62061(.A (n_5547), .B (n_9834), .C (n_4126), .D (n_10264),.Y (n_5678));
OAI22X1 g61482(.A0 (n_5521), .A1 (n_9976), .B0 (g4434), .B1 (n_9627),.Y (n_5677));
AOI22X1 g63305(.A0 (g2763), .A1 (n_10078), .B0 (g2767), .B1 (n_5675),.Y (n_5676));
AOI22X1 g63306(.A0 (g2767), .A1 (n_9871), .B0 (g2779), .B1 (n_5675),.Y (n_5674));
AOI22X1 g63307(.A0 (g2779), .A1 (n_10078), .B0 (g2791), .B1 (n_5675),.Y (n_5672));
AOI22X1 g63308(.A0 (g2795), .A1 (n_5675), .B0 (g2791), .B1 (n_10376),.Y (n_5671));
AOI22X1 g63309(.A0 (g2799), .A1 (n_10078), .B0 (g2811), .B1 (n_5675),.Y (n_5669));
AOI21X1 g63330(.A0 (n_5440), .A1 (g_19304), .B0 (n_5565), .Y(n_5668));
AOI22X1 g63336(.A0 (n_5226), .A1 (n_5513), .B0 (n_5224), .B1(n_5665), .Y (n_5667));
AOI22X1 g63343(.A0 (n_5346), .A1 (n_5665), .B0 (n_5225), .B1(n_5513), .Y (n_5666));
MX2X1 g62108(.A (g_19136), .B (n_5663), .S0 (n_10005), .Y (n_5664));
NAND2X1 g63432(.A (n_5732), .B (g2771), .Y (n_5662));
NAND2X1 g63433(.A (n_5730), .B (g2775), .Y (n_5661));
NAND2X1 g63434(.A (n_5728), .B (g2783), .Y (n_5660));
NAND2X1 g63435(.A (n_5726), .B (g2787), .Y (n_5659));
NAND2X1 g63436(.A (n_5732), .B (g2803), .Y (n_5658));
NAND2X1 g63437(.A (n_5730), .B (g2807), .Y (n_5657));
NAND2X1 g63438(.A (n_5726), .B (g2819), .Y (n_5656));
NAND2X1 g63439(.A (n_5728), .B (g2815), .Y (n_5655));
NOR2X1 g62228(.A (g_8896), .B (n_5560), .Y (n_5654));
NAND3X1 g61626(.A (n_5556), .B (g_18308), .C (n_10063), .Y (n_5652));
NAND4X1 g61640(.A (n_5553), .B (n_2064), .C (n_9279), .D (n_10296),.Y (n_5650));
DFFSRX1 g1950_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5575), .Q (g1950), .QN ());
DFFSRX1 g4821_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10363), .Q (), .QN (g4821));
DFFSRX1 g5011_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5549), .Q (), .QN (g5011));
DFFSRX1 g4704_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5587), .Q (g4704), .QN ());
DFFSRX1 g324_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5574), .Q (g_13255), .QN ());
NAND3X1 g61717(.A (n_5584), .B (n_2540), .C (n_3590), .Y (n_5646));
OR2X1 g61065(.A (n_5581), .B (g4411), .Y (n_5645));
OR2X1 g61066(.A (n_5580), .B (g4405), .Y (n_5644));
AOI21X1 g61073(.A0 (n_5591), .A1 (n_5453), .B0 (n_5630), .Y (n_5715));
NAND3X1 g61075(.A (n_5640), .B (n_5363), .C (n_10005), .Y (n_5643));
MX2X1 g62678(.A (g_9584), .B (n_3559), .S0 (n_9256), .Y (n_5642));
NAND3X1 g61076(.A (n_5640), .B (g4382), .C (n_9359), .Y (n_5641));
MX2X1 g62681(.A (g_21576), .B (g_9584), .S0 (n_5582), .Y (n_5639));
AOI21X1 g61079(.A0 (g4411), .A1 (n_9856), .B0 (n_5579), .Y (n_5637));
NAND3X1 g61817(.A (n_5540), .B (n_2581), .C (n_2067), .Y (n_5634));
NAND3X1 g61819(.A (n_5539), .B (n_4091), .C (n_1626), .Y (n_5633));
INVX1 g61114(.A (n_5630), .Y (n_5631));
OAI21X1 g60915(.A0 (g4512), .A1 (n_9422), .B0 (n_5530), .Y (n_5629));
MX2X1 g61876(.A (g5965), .B (n_5460), .S0 (n_9218), .Y (n_5627));
DFFSRX1 g4572_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5536), .Q (g4572), .QN ());
DFFSRX1 g59_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5534), .Q (g20049), .QN ());
NAND3X1 g61914(.A (n_5517), .B (n_5221), .C (n_5455), .Y (n_5626));
OAI21X1 g61947(.A0 (n_5365), .A1 (n_5454), .B0 (n_5522), .Y (n_5625));
AOI22X1 g61956(.A0 (n_2260), .A1 (n_6655), .B0 (g_15691), .B1(n_9129), .Y (n_5624));
OAI21X1 g63221(.A0 (n_6892), .A1 (g2803), .B0 (n_8557), .Y (n_5622));
NOR2X1 g62047(.A (n_6153), .B (n_6655), .Y (n_5619));
OAI21X1 g63239(.A0 (n_6893), .A1 (g2771), .B0 (n_8557), .Y (n_5617));
OAI21X1 g62105(.A0 (g5077), .A1 (n_9422), .B0 (n_5519), .Y (n_5615));
NAND2X1 g63462(.A (g1632), .B (n_5675), .Y (n_5614));
NAND2X1 g63464(.A (g1768), .B (n_5675), .Y (n_5613));
NAND2X1 g63466(.A (g1902), .B (n_5675), .Y (n_5612));
NAND2X1 g63467(.A (g2036), .B (n_5675), .Y (n_5611));
NAND2X1 g63468(.A (g2193), .B (n_5675), .Y (n_5610));
NAND2X1 g63469(.A (g2327), .B (n_5675), .Y (n_5609));
NAND2X1 g63471(.A (g2461), .B (n_5675), .Y (n_5608));
NAND2X1 g63472(.A (n_5675), .B (g2595), .Y (n_5607));
AOI22X1 g61646(.A0 (n_2296), .A1 (n_11104), .B0 (g_12922), .B1(n_9903), .Y (n_5602));
DFFSRX1 g1816_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5538), .Q (g1816), .QN ());
DFFSRX1 g2161_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5529), .Q (), .QN (g2161));
DFFSRX1 g2169_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5527), .Q (), .QN (g2169));
DFFSRX1 g2173_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5526), .Q (), .QN (g2173));
DFFSRX1 g2181_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5524), .Q (), .QN (g2181));
DFFSRX1 g2084_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5531), .Q (g2084), .QN ());
DFFSRX1 g2555_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6664), .Q (g2555), .QN ());
DFFSRX1 g2153_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10377), .Q (g2153), .QN ());
DFFSRX1 g239_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5537), .Q (g_22371), .QN ());
NAND3X1 g61718(.A (n_5544), .B (n_2298), .C (n_3606), .Y (n_5600));
NAND4X1 g61741(.A (n_5542), .B (n_8906), .C (n_9279), .D (n_2067), .Y(n_5599));
NAND4X1 g61742(.A (n_5541), .B (n_2067), .C (n_9139), .D (n_8694), .Y(n_5596));
MX2X1 g61752(.A (g6311), .B (n_5481), .S0 (n_8955), .Y (n_5593));
NAND3X1 g61074(.A (n_5409), .B (n_5591), .C (n_9453), .Y (n_5592));
MX2X1 g62691(.A (g_22371), .B (n_5465), .S0 (n_9558), .Y (n_5590));
NAND2X1 g61816(.A (n_3588), .B (n_5483), .Y (n_5587));
NAND3X1 g61830(.A (n_7093), .B (n_3394), .C (n_9425), .Y (n_5584));
DFFSRX1 g1612_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5489), .Q (), .QN (g1612));
NOR2X1 g61115(.A (n_1657), .B (n_5591), .Y (n_5630));
MX2X1 g62937(.A (n_5663), .B (g14167), .S0 (n_5582), .Y (n_5583));
NOR2X1 g61124(.A (n_784), .B (n_5591), .Y (n_5581));
NOR2X1 g61125(.A (n_597), .B (n_5591), .Y (n_5580));
AND2X1 g61126(.A (n_5591), .B (g4375), .Y (n_5640));
NOR2X1 g61127(.A (n_5591), .B (n_5378), .Y (n_5579));
OR2X1 g61128(.A (n_5591), .B (n_1980), .Y (n_5578));
NAND3X1 g61940(.A (n_5458), .B (n_5459), .C (n_10385), .Y (n_5576));
NAND3X1 g61152(.A (n_5450), .B (n_2266), .C (n_4131), .Y (n_5575));
DFFSRX1 g4216_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8915), .Q (g8916), .QN ());
NAND3X1 g63208(.A (n_5573), .B (n_2531), .C (n_5370), .Y (n_5574));
AOI22X1 g62080(.A0 (n_5518), .A1 (g5073), .B0 (n_5514), .B1 (g5080),.Y (n_5571));
MX2X1 g63368(.A (g_13255), .B (n_6280), .S0 (n_9681), .Y (n_5570));
NOR2X1 g63476(.A (n_6895), .B (g2775), .Y (n_5569));
NOR2X1 g63486(.A (n_6895), .B (g2783), .Y (n_5568));
NOR2X1 g63504(.A (n_6892), .B (g2807), .Y (n_5567));
NOR2X1 g63508(.A (n_6895), .B (g2815), .Y (n_5566));
NOR2X1 g63518(.A (n_5440), .B (n_3519), .Y (n_5565));
AOI22X1 g63543(.A0 (n_2231), .A1 (n_5562), .B0 (g2811), .B1(n_10376), .Y (n_5564));
AOI22X1 g63544(.A0 (n_1968), .A1 (n_5562), .B0 (g2823), .B1 (n_9129),.Y (n_5563));
INVX1 g62335(.A (g_19136), .Y (n_5560));
NAND2X1 g63878(.A (n_5559), .B (n_8557), .Y (n_5732));
NAND2X1 g63879(.A (n_3866), .B (n_5559), .Y (n_5730));
NAND3X1 g63910(.A (n_5559), .B (n_10650), .C (n_3868), .Y (n_5728));
NAND3X1 g63911(.A (n_5559), .B (n_10650), .C (g2724), .Y (n_5726));
DFFSRX1 g1526_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5485), .Q (g1526), .QN ());
DFFSRX1 g1454_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5449), .Q (), .QN (g1454));
DFFSRX1 g1467_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5448), .Q (), .QN (g1467));
DFFSRX1 g1484_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5447), .Q (), .QN (g1484));
DFFSRX1 g1437_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5451), .Q (), .QN (g1437));
DFFSRX1 g1124_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5462), .Q (), .QN (g_20839));
DFFSRX1 g1141_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5461), .Q (), .QN (g_18200));
DFFSRX1 g1111_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5464), .Q (), .QN (g_18220));
DFFSRX1 g1094_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5466), .Q (), .QN (g_22236));
DFFSRX1 g2241_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5445), .Q (), .QN (g2241));
DFFSRX1 g2375_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5444), .Q (), .QN (g2375));
DFFSRX1 g2643_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5442), .Q (), .QN (g2643));
DFFSRX1 g2177_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5467), .Q (), .QN (g2177));
DFFSRX1 g2004_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5502), .Q (), .QN (g2004));
DFFSRX1 g2020_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5499), .Q (), .QN (g2020));
DFFSRX1 g2024_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5495), .Q (), .QN (g2024));
DFFSRX1 g1600_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5492), .Q (), .QN (g1600));
DFFSRX1 g1608_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5490), .Q (), .QN (g1608));
DFFSRX1 g1620_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5487), .Q (), .QN (g1620));
DFFSRX1 g2016_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5497), .Q (), .QN (g2016));
DFFSRX1 g4616_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5468), .Q (g4616), .QN ());
DFFSRX1 g4608_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5456), .Q (g4608), .QN ());
DFFSRX1 g714_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5437), .Q (), .QN (g_4449));
DFFSRX1 g890_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5504), .Q (g_16571), .QN ());
DFFSRX1 g691_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_10590), .Q (n_11065), .QN ());
DFFSRX1 g1996_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6757), .Q (g1996), .QN ());
DFFSRX1 g4040_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5486), .Q (g4040), .QN ());
DFFSRX1 g3831_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5476), .Q (g3831), .QN ());
DFFSRX1 g3835_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5474), .Q (), .QN (g3835));
NAND2X1 g61714(.A (n_5431), .B (n_5505), .Y (n_5557));
NOR2X1 g61715(.A (n_5723), .B (n_11104), .Y (n_5556));
AOI21X1 g61736(.A0 (n_5422), .A1 (n_2024), .B0 (n_6243), .Y (n_5553));
MX2X1 g61753(.A (g6657), .B (n_5420), .S0 (n_9234), .Y (n_5549));
INVX1 g62682(.A (n_6153), .Y (n_5547));
NAND3X1 g61831(.A (n_7333), .B (n_3547), .C (n_9558), .Y (n_5544));
DFFSRX1 g2421_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6631), .Q (g2421), .QN ());
NAND4X1 g62915(.A (g3897), .B (n_4988), .C (n_5402), .D (g4031), .Y(n_5543));
NOR2X1 g61928(.A (n_5408), .B (n_10947), .Y (n_5542));
NOR2X1 g61931(.A (n_5406), .B (n_3784), .Y (n_5541));
NOR2X1 g61930(.A (n_5407), .B (n_3612), .Y (n_5540));
NOR2X1 g61933(.A (n_5405), .B (n_3605), .Y (n_5539));
NAND3X1 g61151(.A (n_5377), .B (n_2242), .C (n_4133), .Y (n_5538));
MX2X1 g63138(.A (g_22600), .B (n_5271), .S0 (n_9091), .Y (n_5537));
INVX1 g62015(.A (n_10601), .Y (n_5536));
INVX1 g62017(.A (n_10386), .Y (n_5534));
OR2X1 g62020(.A (n_5375), .B (g4452), .Y (n_5532));
DFFSRX1 g872_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14167), .Q (g_9584), .QN ());
NAND3X1 g61161(.A (n_5373), .B (n_2272), .C (n_4614), .Y (n_5531));
DFFSRX1 g2509_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5369), .Q (), .QN (g2509));
OAI21X1 g62066(.A0 (g4531), .A1 (g4581), .B0 (n_10005), .Y (n_5530));
OAI22X1 g61170(.A0 (n_5268), .A1 (n_9884), .B0 (g2165), .B1 (n_9992),.Y (n_5529));
OAI22X1 g61172(.A0 (n_5267), .A1 (n_10952), .B0 (g2161), .B1(n_9627), .Y (n_5527));
OAI22X1 g61173(.A0 (n_5266), .A1 (n_9772), .B0 (g2177), .B1 (n_9651),.Y (n_5526));
OAI22X1 g61175(.A0 (n_5265), .A1 (n_9928), .B0 (g2169), .B1(n_10063), .Y (n_5524));
AOI21X1 g62111(.A0 (g4443), .A1 (n_9772), .B0 (n_5379), .Y (n_5522));
AOI21X1 g61529(.A0 (n_1015), .A1 (n_5454), .B0 (g4443), .Y (n_5521));
NAND3X1 g63532(.A (n_6280), .B (g_19304), .C (g_13901), .Y (n_5520));
NAND2X1 g62222(.A (n_5518), .B (n_5215), .Y (n_5519));
NAND3X1 g62242(.A (n_5374), .B (n_5364), .C (g4382), .Y (n_5517));
OR2X1 g62269(.A (n_5361), .B (n_5514), .Y (n_5515));
DFFSRX1 g479_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5430), .Q (g_19136), .QN ());
AND2X1 g63877(.A (n_5562), .B (n_9358), .Y (n_5675));
OAI21X1 g63884(.A0 (n_10841), .A1 (n_5362), .B0 (n_5436), .Y(n_5761));
INVX1 g63959(.A (n_5665), .Y (n_5513));
DFFSRX1 g1379_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5424), .Q (g1379), .QN ());
DFFSRX1 g2165_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5404), .Q (), .QN (g2165));
DFFSRX1 g2295_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5400), .Q (), .QN (g2295));
DFFSRX1 g2303_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5398), .Q (), .QN (g2303));
DFFSRX1 g2307_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5396), .Q (), .QN (g2307));
DFFSRX1 g2311_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5395), .Q (), .QN (g2311));
DFFSRX1 g2315_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5394), .Q (), .QN (g2315));
DFFSRX1 g2429_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5392), .Q (), .QN (g2429));
DFFSRX1 g2441_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5388), .Q (), .QN (g2441));
DFFSRX1 g2445_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5387), .Q (), .QN (g2445));
DFFSRX1 g2449_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5386), .Q (), .QN (g2449));
DFFSRX1 g2563_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5385), .Q (), .QN (g2563));
DFFSRX1 g2571_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5384), .Q (), .QN (g2571));
DFFSRX1 g2579_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5382), .Q (), .QN (g2579));
DFFSRX1 g2583_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5380), .Q (), .QN (g2583));
DFFSRX1 g2437_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5391), .Q (), .QN (g2437));
DFFSRX1 g2575_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5383), .Q (), .QN (g2575));
DFFSRX1 g1616_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5428), .Q (), .QN (g1616));
DFFSRX1 g723_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5393), .Q (g_15380), .QN ());
DFFSRX1 g287_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5423), .Q (g_19659), .QN ());
DFFSRX1 g1036_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5411), .Q (g_12465), .QN ());
DFFSRX1 g671_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5372), .Q (g_21447), .QN ());
DFFSRX1 g2287_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6639), .Q (g2287), .QN ());
DFFSRX1 g2089_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5359), .Q (), .QN (g2089));
DFFSRX1 g2246_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5358), .Q (), .QN (g2246));
DFFSRX1 g2269_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5357), .Q (g2269), .QN ());
DFFSRX1 g2273_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5356), .Q (), .QN (g2273));
DFFSRX1 g5156_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5432), .Q (g5156), .QN ());
DFFSRX1 g3827_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5415), .Q (), .QN (g3827));
DFFSRX1 g2197_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5414), .Q (g2197), .QN ());
DFFSRX1 g2227_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5412), .Q (g2227), .QN ());
DFFSRX1 g3817_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5410), .Q (g3817), .QN ());
DFFSRX1 g262_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5397), .Q (g_22600), .QN ());
XOR2X1 g62665(.A (g_10556), .B (n_5287), .Y (n_5508));
NAND4X1 g62671(.A (n_5403), .B (n_4607), .C (n_4088), .D (n_4984), .Y(n_5506));
CLKBUFX2 g62683(.A (n_6801), .Y (n_6153));
NAND3X1 g61800(.A (n_5323), .B (g_12922), .C (n_9797), .Y (n_5505));
NAND3X1 g61804(.A (n_5311), .B (n_2255), .C (n_2852), .Y (n_5504));
OAI22X1 g61343(.A0 (n_5068), .A1 (n_9371), .B0 (g2008), .B1 (n_9862),.Y (n_5502));
NAND3X1 g62806(.A (n_5290), .B (g3211), .C (n_8586), .Y (n_5501));
NAND3X1 g62809(.A (n_5289), .B (g3562), .C (n_4682), .Y (n_5500));
OAI22X1 g61347(.A0 (n_5045), .A1 (n_9903), .B0 (g2024), .B1 (n_9811),.Y (n_5499));
OAI22X1 g61346(.A0 (n_5058), .A1 (n_9976), .B0 (g2020), .B1 (n_9664),.Y (n_5497));
OAI22X1 g61348(.A0 (n_5044), .A1 (n_10952), .B0 (g2012), .B1(n_9627), .Y (n_5495));
OAI22X1 g61349(.A0 (n_5039), .A1 (n_9431), .B0 (g1604), .B1 (n_9627),.Y (n_5492));
DFFSRX1 g2008_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5337), .Q (), .QN (g2008));
OAI22X1 g61351(.A0 (n_5030), .A1 (n_9772), .B0 (g1600), .B1 (n_9992),.Y (n_5490));
OAI22X1 g61352(.A0 (n_5022), .A1 (n_9836), .B0 (g1616), .B1 (n_9830),.Y (n_5489));
DFFSRX1 g2116_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5238), .Q (), .QN (g2116));
OAI22X1 g61354(.A0 (n_5019), .A1 (n_9976), .B0 (g1608), .B1(n_10063), .Y (n_5487));
DFFSRX1 g1821_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5246), .Q (), .QN (g1821));
MX2X1 g62925(.A (g4031), .B (n_3430), .S0 (n_9218), .Y (n_5486));
DFFSRX1 g1886_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5340), .Q (), .QN (g1886));
DFFSRX1 g1870_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5345), .Q (), .QN (g1870));
OAI21X1 g60919(.A0 (n_4285), .A1 (n_9693), .B0 (n_5283), .Y (n_5485));
NAND4X1 g61938(.A (n_5288), .B (n_2067), .C (n_9940), .D (n_8777), .Y(n_5483));
NAND3X1 g61948(.A (g4372), .B (g4581), .C (n_9466), .Y (n_6011));
MX2X1 g61966(.A (n_19), .B (n_11196), .S0 (n_3626), .Y (n_5481));
DFFSRX1 g2567_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5278), .Q (), .QN (g2567));
OAI22X1 g63110(.A0 (n_4985), .A1 (n_9269), .B0 (g3827), .B1 (n_9651),.Y (n_5476));
MX2X1 g63111(.A (g3831), .B (n_4971), .S0 (n_9894), .Y (n_5474));
OR4X1 g61153(.A (g4411), .B (g4405), .C (g4375), .D (n_316), .Y(n_5591));
DFFSRX1 g2299_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5282), .Q (), .QN (g2299));
NAND3X1 g61484(.A (n_2564), .B (n_4976), .C (n_4844), .Y (n_5468));
OAI22X1 g61174(.A0 (n_4967), .A1 (n_9903), .B0 (g2181), .B1 (n_9992),.Y (n_5467));
OAI21X1 g61013(.A0 (n_4966), .A1 (n_10952), .B0 (n_3164), .Y(n_5466));
MX2X1 g63335(.A (g_20208), .B (g14147), .S0 (n_5582), .Y (n_5465));
OAI21X1 g61014(.A0 (n_4960), .A1 (n_9693), .B0 (n_3162), .Y (n_5464));
OAI21X1 g61015(.A0 (n_4959), .A1 (n_10078), .B0 (n_3161), .Y(n_5462));
OAI21X1 g61016(.A0 (n_4954), .A1 (n_9672), .B0 (n_3363), .Y (n_5461));
MX2X1 g62127(.A (n_1299), .B (n_5457), .S0 (n_5459), .Y (n_5460));
XOR2X1 g62132(.A (n_2072), .B (n_5457), .Y (n_5458));
DFFSRX1 g4213_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g11770), .Q (g8915), .QN ());
OAI22X1 g61554(.A0 (n_4955), .A1 (n_4956), .B0 (n_262), .B1 (n_9627),.Y (n_5456));
NAND2X1 g62243(.A (n_5454), .B (n_5453), .Y (n_5455));
OAI21X1 g60940(.A0 (n_5223), .A1 (n_9628), .B0 (n_3197), .Y (n_5451));
NAND3X1 g61203(.A (n_5258), .B (n_6677), .C (n_9834), .Y (n_5450));
OAI21X1 g60941(.A0 (n_5222), .A1 (n_9371), .B0 (n_3196), .Y (n_5449));
OAI21X1 g60942(.A0 (n_5219), .A1 (n_9903), .B0 (n_3191), .Y (n_5448));
OAI21X1 g60943(.A0 (n_5218), .A1 (n_9775), .B0 (n_3384), .Y (n_5447));
NAND3X1 g61042(.A (n_5259), .B (n_2558), .C (n_4864), .Y (n_5445));
NAND3X1 g61044(.A (n_10548), .B (n_2247), .C (n_10549), .Y (n_5444));
NAND3X1 g63961(.A (n_6897), .B (n_8557), .C (n_11), .Y (n_5665));
NAND3X1 g61046(.A (n_5253), .B (n_2284), .C (n_4611), .Y (n_5442));
DFFSRX1 g1373_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5291), .Q (g1373), .QN ());
DFFSRX1 g2433_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5279), .Q (), .QN (g2433));
DFFSRX1 g1744_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5349), .Q (), .QN (g1744));
DFFSRX1 g1748_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5354), .Q (), .QN (g1748));
DFFSRX1 g1752_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5348), .Q (), .QN (g1752));
DFFSRX1 g1756_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5347), .Q (), .QN (g1756));
DFFSRX1 g1736_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5235), .Q (), .QN (g1736));
DFFSRX1 g1878_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5342), .Q (), .QN (g1878));
DFFSRX1 g1882_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5341), .Q (), .QN (g1882));
DFFSRX1 g1740_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5233), .Q (), .QN (g1740));
DFFSRX1 g1890_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5338), .Q (), .QN (g1890));
DFFSRX1 g1874_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5344), .Q (), .QN (g1874));
DFFSRX1 g2012_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5336), .Q (), .QN (g2012));
DFFSRX1 g1604_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5335), .Q (), .QN (g1604));
DFFSRX1 g676_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5310), .Q (), .QN (g_16063));
DFFSRX1 g1183_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_8620), .Q (g1183), .QN ());
DFFSRX1 g686_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5270), .Q (g_17426), .QN ());
DFFSRX1 g1030_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5276), .Q (g_20159), .QN ());
DFFSRX1 g5052_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5272), .Q (g5052), .QN ());
DFFSRX1 g1862_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6684), .Q (g1862), .QN ());
DFFSRX1 g1728_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_6866), .Q (g1728), .QN ());
DFFSRX1 g2675_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5251), .Q (), .QN (g2675));
DFFSRX1 g2671_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5252), .Q (g2671), .QN ());
DFFSRX1 g1710_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5249), .Q (g1710), .QN ());
DFFSRX1 g1714_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5248), .Q (), .QN (g1714));
DFFSRX1 g1844_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5245), .Q (g1844), .QN ());
DFFSRX1 g1848_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5244), .Q (), .QN (g1848));
DFFSRX1 g1955_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5242), .Q (), .QN (g1955));
DFFSRX1 g1978_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5241), .Q (g1978), .QN ());
DFFSRX1 g1982_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5240), .Q (), .QN (g1982));
DFFSRX1 g2112_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5239), .Q (g2112), .QN ());
DFFSRX1 g2265_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5236), .Q (), .QN (g2265));
DFFSRX1 g2407_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5355), .Q (), .QN (g2407));
DFFSRX1 g2537_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5353), .Q (g2537), .QN ());
DFFSRX1 g2541_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5352), .Q (), .QN (g2541));
DFFSRX1 g2648_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5350), .Q (), .QN (g2648));
DFFSRX1 g5057_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5254), .Q (g5057), .QN ());
DFFSRX1 g2403_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5232), .Q (g2403), .QN ());
DFFSRX1 g3689_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5331), .Q (g3689), .QN ());
DFFSRX1 g3338_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5333), .Q (g3338), .QN ());
DFFSRX1 g5252_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5329), .Q (g5252), .QN ());
DFFSRX1 g5260_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5328), .Q (g5260), .QN ());
DFFSRX1 g5236_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5330), .Q (g5236), .QN ());
DFFSRX1 g5264_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5327), .Q (g5264), .QN ());
DFFSRX1 g5583_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5326), .Q (g5583), .QN ());
DFFSRX1 g5599_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5325), .Q (g5599), .QN ());
DFFSRX1 g5929_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5324), .Q (g5929), .QN ());
DFFSRX1 g5957_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5321), .Q (g5957), .QN ());
DFFSRX1 g3129_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5319), .Q (g3129), .QN ());
DFFSRX1 g3133_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5318), .Q (), .QN (g3133));
DFFSRX1 g6275_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5317), .Q (g6275), .QN ());
DFFSRX1 g6299_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5315), .Q (g6299), .QN ());
DFFSRX1 g6303_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5313), .Q (g6303), .QN ());
DFFSRX1 g6307_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5312), .Q (g6307), .QN ());
DFFSRX1 g6637_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5309), .Q (g6637), .QN ());
DFFSRX1 g6645_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5308), .Q (g6645), .QN ());
DFFSRX1 g3480_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5307), .Q (g3480), .QN ());
DFFSRX1 g3484_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5306), .Q (), .QN (g3484));
DFFSRX1 g2040_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5304), .Q (g2040), .QN ());
DFFSRX1 g2070_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5302), .Q (g2070), .QN ());
DFFSRX1 g3945_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5300), .Q (g3945), .QN ());
DFFSRX1 g3953_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5299), .Q (g3953), .QN ());
DFFSRX1 g1592_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5339), .Q (g1592), .QN ());
DFFSRX1 g1636_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5297), .Q (g1636), .QN ());
DFFSRX1 g2599_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5296), .Q (g2599), .QN ());
DFFSRX1 g1668_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5294), .Q (n_4120), .QN ());
DFFSRX1 g2629_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5293), .Q (g2629), .QN ());
DFFSRX1 g4473_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5275), .Q (g4473), .QN ());
INVX1 g64074(.A (n_6280), .Y (n_5440));
DFFSRX1 g2756_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5247), .Q (g2756), .QN ());
NAND3X1 g61739(.A (n_2797), .B (n_4921), .C (n_4961), .Y (n_5437));
INVX1 g64379(.A (n_5436), .Y (n_5559));
DFFSRX1 g6287_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5127), .Q (g6287), .QN ());
OAI21X1 g62792(.A0 (n_4896), .A1 (n_5007), .B0 (n_4990), .Y (n_5432));
AOI22X1 g61839(.A0 (n_2265), .A1 (n_6549), .B0 (g_19659), .B1(n_10376), .Y (n_5431));
NAND2X1 g62824(.A (n_4889), .B (n_4991), .Y (n_5430));
DFFSRX1 g2399_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4943), .Q (), .QN (g2399));
DFFSRX1 g6255_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5135), .Q (g6255), .QN ());
OAI22X1 g61353(.A0 (n_4913), .A1 (n_9903), .B0 (g1620), .B1 (n_9862),.Y (n_5428));
NAND4X1 g62914(.A (g3546), .B (n_10576), .C (n_10897), .D (g3680), .Y(n_5425));
DFFSRX1 g6239_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5141), .Q (g6239), .QN ());
DFFSRX1 g3602_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5050), .Q (g3602), .QN ());
DFFSRX1 g3594_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5052), .Q (g3594), .QN ());
DFFSRX1 g5949_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5150), .Q (g5949), .QN ());
DFFSRX1 g5933_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5155), .Q (g5933), .QN ());
DFFSRX1 g5917_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5159), .Q (g5917), .QN ());
NAND3X1 g60918(.A (n_5000), .B (n_2288), .C (n_4888), .Y (n_5424));
DFFSRX1 g3578_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5059), .Q (g3578), .QN ());
NAND2X1 g61918(.A (n_4999), .B (n_4911), .Y (n_5423));
AOI21X1 g61934(.A0 (n_4874), .A1 (n_3769), .B0 (g4961), .Y (n_5422));
MX2X1 g61967(.A (n_843), .B (n_7329), .S0 (n_3547), .Y (n_5420));
DFFSRX1 g5607_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5173), .Q (g5607), .QN ());
MX2X1 g63109(.A (g3821), .B (n_4886), .S0 (n_9091), .Y (n_5415));
MX2X1 g63132(.A (g2204), .B (n_4884), .S0 (n_10005), .Y (n_5414));
MX2X1 g63133(.A (g2197), .B (n_4881), .S0 (n_9000), .Y (n_5412));
NAND3X1 g62031(.A (n_4974), .B (n_2526), .C (n_4842), .Y (n_5411));
NAND2X1 g63219(.A (n_4879), .B (n_4987), .Y (n_5410));
XOR2X1 g61167(.A (g4382), .B (g4375), .Y (n_5409));
AOI21X1 g62074(.A0 (n_4021), .A1 (n_4982), .B0 (n_4983), .Y (n_5408));
AOI21X1 g62075(.A0 (n_4020), .A1 (n_4980), .B0 (n_4981), .Y (n_5407));
AOI21X1 g62076(.A0 (n_4019), .A1 (n_4978), .B0 (n_4979), .Y (n_5406));
AOI21X1 g62077(.A0 (n_4018), .A1 (n_11070), .B0 (n_4977), .Y(n_5405));
MX2X1 g61171(.A (n_4906), .B (n_4865), .S0 (n_9358), .Y (n_5404));
NAND4X1 g63298(.A (g3949), .B (n_5402), .C (g16748), .D (n_8917), .Y(n_5403));
OAI22X1 g61176(.A0 (n_4861), .A1 (n_9505), .B0 (g2299), .B1 (n_9651),.Y (n_5400));
OAI22X1 g61178(.A0 (n_4860), .A1 (n_9599), .B0 (g2295), .B1 (n_9992),.Y (n_5398));
MX2X1 g63370(.A (n_11106), .B (n_4857), .S0 (n_8955), .Y (n_5397));
OAI22X1 g61179(.A0 (n_4859), .A1 (n_10952), .B0 (g2311), .B1(n_9992), .Y (n_5396));
DFFSRX1 g3562_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5064), .Q (g3562), .QN ());
DFFSRX1 g887_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14147), .Q (g14167), .QN ());
OAI22X1 g61180(.A0 (n_4858), .A1 (n_10078), .B0 (g2315), .B1(n_9830), .Y (n_5395));
OAI22X1 g61181(.A0 (n_4856), .A1 (n_9903), .B0 (g2303), .B1 (n_9992),.Y (n_5394));
NAND3X1 g61517(.A (n_2543), .B (n_4820), .C (n_4875), .Y (n_5393));
OAI22X1 g61183(.A0 (n_4930), .A1 (n_9505), .B0 (g2433), .B1 (n_9811),.Y (n_5392));
OAI22X1 g61185(.A0 (n_4854), .A1 (n_9928), .B0 (g2429), .B1 (n_9992),.Y (n_5391));
OAI22X1 g61186(.A0 (n_4853), .A1 (n_9884), .B0 (g2445), .B1 (n_9862),.Y (n_5388));
OAI22X1 g61187(.A0 (n_4852), .A1 (n_9599), .B0 (g2449), .B1 (n_9811),.Y (n_5387));
OAI22X1 g61188(.A0 (n_4851), .A1 (n_9461), .B0 (g2437), .B1 (n_9651),.Y (n_5386));
OAI22X1 g61189(.A0 (n_4850), .A1 (n_9461), .B0 (g2567), .B1 (n_9992),.Y (n_5385));
DFFSRX1 g5567_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5184), .Q (g5567), .QN ());
OAI22X1 g61191(.A0 (n_4849), .A1 (n_9431), .B0 (g2563), .B1 (n_9862),.Y (n_5384));
OAI22X1 g61192(.A0 (n_4847), .A1 (n_10952), .B0 (g2579), .B1(n_9992), .Y (n_5383));
OAI22X1 g61193(.A0 (n_4846), .A1 (n_9193), .B0 (g2583), .B1 (n_9862),.Y (n_5382));
OAI22X1 g61194(.A0 (n_4845), .A1 (n_9269), .B0 (g2571), .B1 (n_9992),.Y (n_5380));
NOR2X1 g62241(.A (n_5374), .B (n_5378), .Y (n_5379));
NAND3X1 g61200(.A (n_4965), .B (n_10911), .C (n_9558), .Y (n_5377));
NOR2X1 g62263(.A (n_595), .B (n_5374), .Y (n_5375));
NAND3X1 g61210(.A (n_4962), .B (n_4296), .C (n_9209), .Y (n_5373));
DFFSRX1 g2465_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5015), .Q (g2465), .QN ());
OAI21X1 g62284(.A0 (n_95), .A1 (n_9333), .B0 (n_4964), .Y (n_5372));
DFFSRX1 g3961_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5021), .Q (g3961), .QN ());
NAND3X1 g63924(.A (g_13255), .B (g_16983), .C (n_9811), .Y (n_5370));
NAND3X1 g61045(.A (n_4953), .B (n_2533), .C (n_4308), .Y (n_5369));
DFFSRX1 g6653_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5076), .Q (g6653), .QN ());
DFFSRX1 g1514_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4986), .Q (n_10197), .QN ());
DFFSRX1 g1413_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4975), .Q (), .QN (g1413));
DFFSRX1 g827_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4972), .Q (g_14342), .QN ());
DFFSRX1 g4601_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4957), .Q (g4601), .QN ());
DFFSRX1 g3909_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5037), .Q (g3909), .QN ());
DFFSRX1 g3259_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5085), .Q (g3259), .QN ());
DFFSRX1 g3941_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5025), .Q (g3941), .QN ());
DFFSRX1 g6617_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5088), .Q (g6617), .QN ());
DFFSRX1 g3957_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5023), .Q (g3957), .QN ());
DFFSRX1 g6605_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5093), .Q (g6605), .QN ());
DFFSRX1 g5268_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5195), .Q (g5268), .QN ());
DFFSRX1 g3191_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5122), .Q (g3191), .QN ());
DFFSRX1 g6581_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5106), .Q (g6581), .QN ());
DFFSRX1 g5256_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5197), .Q (g5256), .QN ());
DFFSRX1 g5228_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5204), .Q (g5228), .QN ());
DFFSRX1 g490_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5009), .Q (g_15016), .QN ());
DFFSRX1 g5216_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5207), .Q (g5216), .QN ());
DFFSRX1 g1687_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4952), .Q (), .QN (g1687));
DFFSRX1 g2667_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4951), .Q (), .QN (g2667));
DFFSRX1 g1706_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4950), .Q (), .QN (g1706));
DFFSRX1 g1840_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4949), .Q (), .QN (g1840));
DFFSRX1 g1974_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4947), .Q (), .QN (g1974));
DFFSRX1 g2108_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4945), .Q (), .QN (g2108));
DFFSRX1 g2380_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4944), .Q (), .QN (g2380));
DFFSRX1 g2514_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5231), .Q (), .QN (g2514));
DFFSRX1 g2533_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5230), .Q (), .QN (g2533));
DFFSRX1 g5196_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5214), .Q (g5196), .QN ());
DFFSRX1 g5200_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5213), .Q (g5200), .QN ());
DFFSRX1 g5208_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5210), .Q (g5208), .QN ());
DFFSRX1 g5212_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5209), .Q (g5212), .QN ());
DFFSRX1 g5204_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5212), .Q (g5204), .QN ());
DFFSRX1 g5224_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5205), .Q (g5224), .QN ());
DFFSRX1 g5220_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5206), .Q (g5220), .QN ());
DFFSRX1 g5240_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5201), .Q (g5240), .QN ());
DFFSRX1 g5244_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5200), .Q (g5244), .QN ());
DFFSRX1 g5248_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5199), .Q (g5248), .QN ());
DFFSRX1 g5232_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5202), .Q (g5232), .QN ());
DFFSRX1 g5272_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5193), .Q (g5272), .QN ());
DFFSRX1 g5547_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5190), .Q (g5547), .QN ());
DFFSRX1 g5551_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5189), .Q (g5551), .QN ());
DFFSRX1 g5555_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5187), .Q (g5555), .QN ());
DFFSRX1 g5559_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5186), .Q (g5559), .QN ());
DFFSRX1 g5563_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5185), .Q (g5563), .QN ());
DFFSRX1 g5571_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5183), .Q (g5571), .QN ());
DFFSRX1 g5575_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5182), .Q (g5575), .QN ());
DFFSRX1 g5579_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5181), .Q (g5579), .QN ());
DFFSRX1 g5543_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5192), .Q (g5543), .QN ());
DFFSRX1 g5591_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5177), .Q (g5591), .QN ());
DFFSRX1 g5595_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5175), .Q (g5595), .QN ());
DFFSRX1 g5587_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5179), .Q (g5587), .QN ());
DFFSRX1 g5603_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5174), .Q (g5603), .QN ());
DFFSRX1 g5611_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5172), .Q (g5611), .QN ());
DFFSRX1 g5615_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5171), .Q (g5615), .QN ());
DFFSRX1 g5619_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5170), .Q (g5619), .QN ());
DFFSRX1 g5889_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5168), .Q (g5889), .QN ());
DFFSRX1 g5897_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5165), .Q (g5897), .QN ());
DFFSRX1 g5901_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5164), .Q (g5901), .QN ());
DFFSRX1 g5905_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5163), .Q (g5905), .QN ());
DFFSRX1 g5909_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5161), .Q (g5909), .QN ());
DFFSRX1 g5913_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5160), .Q (g5913), .QN ());
DFFSRX1 g5893_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5167), .Q (g5893), .QN ());
DFFSRX1 g5921_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5158), .Q (g5921), .QN ());
DFFSRX1 g5925_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5156), .Q (g5925), .QN ());
DFFSRX1 g5937_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5154), .Q (g5937), .QN ());
DFFSRX1 g5941_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5152), .Q (g5941), .QN ());
DFFSRX1 g5945_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5151), .Q (g5945), .QN ());
DFFSRX1 g5953_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5149), .Q (g5953), .QN ());
DFFSRX1 g5961_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5148), .Q (g5961), .QN ());
DFFSRX1 g5965_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5146), .Q (g5965), .QN ());
DFFSRX1 g3125_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5144), .Q (), .QN (g3125));
DFFSRX1 g6235_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5143), .Q (g6235), .QN ());
DFFSRX1 g6243_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5139), .Q (g6243), .QN ());
DFFSRX1 g6247_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5137), .Q (g6247), .QN ());
DFFSRX1 g6251_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5136), .Q (g6251), .QN ());
DFFSRX1 g6259_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5134), .Q (g6259), .QN ());
DFFSRX1 g6267_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5131), .Q (g6267), .QN ());
DFFSRX1 g6271_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5130), .Q (g6271), .QN ());
DFFSRX1 g6263_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5133), .Q (g6263), .QN ());
DFFSRX1 g6279_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5129), .Q (g6279), .QN ());
DFFSRX1 g6283_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5128), .Q (g6283), .QN ());
DFFSRX1 g6291_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5126), .Q (g6291), .QN ());
DFFSRX1 g6295_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5125), .Q (g6295), .QN ());
DFFSRX1 g3187_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5123), .Q (g3187), .QN ());
DFFSRX1 g6311_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5124), .Q (g6311), .QN ());
DFFSRX1 g3195_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5121), .Q (g3195), .QN ());
DFFSRX1 g3199_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5119), .Q (g3199), .QN ());
DFFSRX1 g3203_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5118), .Q (g3203), .QN ());
DFFSRX1 g3207_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5116), .Q (g3207), .QN ());
DFFSRX1 g3211_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5115), .Q (g3211), .QN ());
DFFSRX1 g3215_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5113), .Q (g3215), .QN ());
DFFSRX1 g3219_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5112), .Q (g3219), .QN ());
DFFSRX1 g3223_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5111), .Q (g3223), .QN ());
DFFSRX1 g3227_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5110), .Q (g3227), .QN ());
DFFSRX1 g3231_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5109), .Q (g3231), .QN ());
DFFSRX1 g3235_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5107), .Q (g3235), .QN ());
DFFSRX1 g3239_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5104), .Q (g3239), .QN ());
DFFSRX1 g6585_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5103), .Q (g6585), .QN ());
DFFSRX1 g3243_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5101), .Q (g3243), .QN ());
DFFSRX1 g6589_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5100), .Q (g6589), .QN ());
DFFSRX1 g6593_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5098), .Q (g6593), .QN ());
DFFSRX1 g3247_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5097), .Q (g3247), .QN ());
DFFSRX1 g6597_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5095), .Q (g6597), .QN ());
DFFSRX1 g6601_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5094), .Q (g6601), .QN ());
DFFSRX1 g6609_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5092), .Q (g6609), .QN ());
DFFSRX1 g3251_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5091), .Q (g3251), .QN ());
DFFSRX1 g6613_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5090), .Q (g6613), .QN ());
DFFSRX1 g3255_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5087), .Q (g3255), .QN ());
DFFSRX1 g6621_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5086), .Q (g6621), .QN ());
DFFSRX1 g6625_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5084), .Q (g6625), .QN ());
DFFSRX1 g3263_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5082), .Q (g3263), .QN ());
DFFSRX1 g6633_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5081), .Q (g6633), .QN ());
DFFSRX1 g6629_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5083), .Q (g6629), .QN ());
DFFSRX1 g6641_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5079), .Q (g6641), .QN ());
DFFSRX1 g6649_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5077), .Q (g6649), .QN ());
DFFSRX1 g6657_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5075), .Q (g6657), .QN ());
DFFSRX1 g3476_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5016), .Q (), .QN (g3476));
DFFSRX1 g3538_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5073), .Q (g3538), .QN ());
DFFSRX1 g3542_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5072), .Q (g3542), .QN ());
DFFSRX1 g3546_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5071), .Q (g3546), .QN ());
DFFSRX1 g3550_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5069), .Q (g3550), .QN ());
DFFSRX1 g3554_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5067), .Q (g3554), .QN ());
DFFSRX1 g3558_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5065), .Q (g3558), .QN ());
DFFSRX1 g3566_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5063), .Q (g3566), .QN ());
DFFSRX1 g3570_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5062), .Q (g3570), .QN ());
DFFSRX1 g3574_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5060), .Q (g3574), .QN ());
DFFSRX1 g3582_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5056), .Q (g3582), .QN ());
DFFSRX1 g3586_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5055), .Q (g3586), .QN ());
DFFSRX1 g3590_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5053), .Q (g3590), .QN ());
DFFSRX1 g3606_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5048), .Q (g3606), .QN ());
DFFSRX1 g3610_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5047), .Q (g3610), .QN ());
DFFSRX1 g3614_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5046), .Q (g3614), .QN ());
DFFSRX1 g3598_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5051), .Q (g3598), .QN ());
DFFSRX1 g3889_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5043), .Q (g3889), .QN ());
DFFSRX1 g3893_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5042), .Q (g3893), .QN ());
DFFSRX1 g3897_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5041), .Q (g3897), .QN ());
DFFSRX1 g3901_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5040), .Q (g3901), .QN ());
DFFSRX1 g3905_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5038), .Q (g3905), .QN ());
DFFSRX1 g3925_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5032), .Q (g3925), .QN ());
DFFSRX1 g3929_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5029), .Q (g3929), .QN ());
DFFSRX1 g3933_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5028), .Q (g3933), .QN ());
DFFSRX1 g3937_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5026), .Q (g3937), .QN ());
DFFSRX1 g3921_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5033), .Q (g3921), .QN ());
DFFSRX1 g3949_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5024), .Q (g3949), .QN ());
DFFSRX1 g3913_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5035), .Q (g3913), .QN ());
DFFSRX1 g3965_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5020), .Q (g3965), .QN ());
DFFSRX1 g3917_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5034), .Q (g3917), .QN ());
DFFSRX1 g2331_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5018), .Q (g2331), .QN ());
DFFSRX1 g2361_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5017), .Q (g2361), .QN ());
DFFSRX1 g2495_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5014), .Q (n_4339), .QN ());
DFFSRX1 g5503_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5008), .Q (), .QN (g5503));
DFFSRX1 g5849_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5006), .Q (), .QN (g5849));
DFFSRX1 g3115_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5013), .Q (g3115), .QN ());
DFFSRX1 g6195_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5005), .Q (), .QN (g6195));
DFFSRX1 g3147_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5004), .Q (), .QN (g3147));
DFFSRX1 g3498_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5002), .Q (), .QN (g3498));
DFFSRX1 g3849_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5001), .Q (), .QN (g3849));
DFFSRX1 g3466_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5012), .Q (g3466), .QN ());
DFFSRX1 g6541_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_5003), .Q (), .QN (g6541));
DFFSRX1 g232_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4970), .Q (g_20244), .QN ());
OAI21X1 g64075(.A0 (g_13255), .A1 (g_16983), .B0 (n_3522), .Y(n_6280));
OR2X1 g64154(.A (n_5227), .B (n_10841), .Y (n_5562));
NOR2X1 g62585(.A (g5077), .B (n_9856), .Y (n_5518));
NAND2X1 g62618(.A (n_5364), .B (n_5363), .Y (n_5365));
NAND4X1 g64380(.A (n_10841), .B (n_5362), .C (g2735), .D (n_11012),.Y (n_5436));
NOR2X1 g62645(.A (g5069), .B (g5077), .Y (n_5361));
MX2X1 g62711(.A (g2084), .B (n_4905), .S0 (n_9000), .Y (n_5359));
OAI22X1 g62715(.A0 (n_4907), .A1 (n_9371), .B0 (g2241), .B1 (n_9992),.Y (n_5358));
OAI22X1 g62717(.A0 (n_4904), .A1 (n_9903), .B0 (g2265), .B1(n_10063), .Y (n_5357));
MX2X1 g62718(.A (g2269), .B (n_4899), .S0 (n_9279), .Y (n_5356));
MX2X1 g62722(.A (g2403), .B (n_4708), .S0 (n_9167), .Y (n_5355));
OAI22X1 g61333(.A0 (n_4780), .A1 (n_9976), .B0 (g1752), .B1 (n_9664),.Y (n_5354));
OAI22X1 g62725(.A0 (n_4716), .A1 (n_9431), .B0 (g2533), .B1 (n_9698),.Y (n_5353));
MX2X1 g62726(.A (g2537), .B (n_4707), .S0 (n_9218), .Y (n_5352));
OAI22X1 g62728(.A0 (n_4727), .A1 (n_9772), .B0 (g2643), .B1 (n_9651),.Y (n_5350));
OAI22X1 g61334(.A0 (n_4781), .A1 (n_10952), .B0 (g1736), .B1(n_9664), .Y (n_5349));
OAI22X1 g61335(.A0 (n_4779), .A1 (n_9461), .B0 (g1756), .B1 (n_9209),.Y (n_5348));
OAI22X1 g61336(.A0 (n_4777), .A1 (n_10952), .B0 (g1744), .B1(n_9992), .Y (n_5347));
AOI21X1 g64708(.A0 (n_4224), .A1 (n_8895), .B0 (n_4935), .Y (n_5346));
OAI22X1 g61337(.A0 (n_4776), .A1 (n_9129), .B0 (g1874), .B1(n_10005), .Y (n_5345));
MX2X1 g61338(.A (n_4187), .B (n_4775), .S0 (n_8955), .Y (n_5344));
OAI22X1 g61339(.A0 (n_4774), .A1 (n_9431), .B0 (g1870), .B1 (n_9521),.Y (n_5342));
OAI22X1 g61340(.A0 (n_4773), .A1 (n_9976), .B0 (g1886), .B1 (n_9651),.Y (n_5341));
OAI22X1 g61341(.A0 (n_4772), .A1 (n_9431), .B0 (g1890), .B1 (n_9811),.Y (n_5340));
NOR2X1 g62790(.A (n_4900), .B (n_9019), .Y (n_5339));
OAI22X1 g61342(.A0 (n_4770), .A1 (n_9772), .B0 (g1878), .B1 (n_9651),.Y (n_5338));
MX2X1 g61344(.A (n_4183), .B (n_4769), .S0 (n_9156), .Y (n_5337));
OAI22X1 g61345(.A0 (n_4768), .A1 (n_9976), .B0 (g2004), .B1 (n_9627),.Y (n_5336));
MX2X1 g61350(.A (n_4527), .B (n_4767), .S0 (n_9279), .Y (n_5335));
MX2X1 g62922(.A (g3329), .B (n_3020), .S0 (n_9553), .Y (n_5333));
MX2X1 g62924(.A (g3680), .B (n_3019), .S0 (n_8955), .Y (n_5331));
MX2X1 g62954(.A (g5216), .B (n_4670), .S0 (n_9750), .Y (n_5330));
MX2X1 g62958(.A (g5236), .B (n_4669), .S0 (n_9333), .Y (n_5329));
MX2X1 g62960(.A (g5244), .B (n_4656), .S0 (n_9000), .Y (n_5328));
MX2X1 g62961(.A (g5248), .B (n_4667), .S0 (n_8955), .Y (n_5327));
MX2X1 g62977(.A (g5563), .B (n_4666), .S0 (n_9256), .Y (n_5326));
MX2X1 g62981(.A (g5583), .B (n_4665), .S0 (n_9240), .Y (n_5325));
MX2X1 g63002(.A (g5909), .B (n_4662), .S0 (n_9834), .Y (n_5324));
NOR2X1 g61921(.A (n_5723), .B (n_6549), .Y (n_5323));
MX2X1 g63009(.A (g5941), .B (n_4661), .S0 (n_9797), .Y (n_5321));
OAI22X1 g63016(.A0 (n_4689), .A1 (n_10952), .B0 (g3125), .B1(n_9651), .Y (n_5319));
MX2X1 g63019(.A (g3129), .B (n_4651), .S0 (n_9358), .Y (n_5318));
MX2X1 g63028(.A (g6255), .B (n_4660), .S0 (n_8955), .Y (n_5317));
MX2X1 g63034(.A (g6283), .B (n_4659), .S0 (n_9894), .Y (n_5315));
MX2X1 g63035(.A (g6287), .B (n_4658), .S0 (n_10005), .Y (n_5313));
MX2X1 g63036(.A (g6291), .B (n_4657), .S0 (n_8955), .Y (n_5312));
NAND3X1 g61958(.A (n_4912), .B (g_22552), .C (n_10385), .Y (n_5311));
OAI22X1 g61960(.A0 (n_4963), .A1 (n_3916), .B0 (n_3310), .B1(n_9651), .Y (n_5310));
MX2X1 g63075(.A (g6621), .B (n_4653), .S0 (n_9797), .Y (n_5309));
MX2X1 g63077(.A (g6629), .B (n_4652), .S0 (n_9218), .Y (n_5308));
OAI22X1 g63085(.A0 (n_4688), .A1 (n_9976), .B0 (g3476), .B1 (n_9627),.Y (n_5307));
DFFSRX1 g1772_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4927), .Q (g1772), .QN ());
MX2X1 g63086(.A (g3480), .B (n_4650), .S0 (n_9218), .Y (n_5306));
MX2X1 g63107(.A (g2047), .B (n_4649), .S0 (n_9834), .Y (n_5304));
MX2X1 g63108(.A (g2040), .B (n_4647), .S0 (n_8955), .Y (n_5302));
DFFSRX1 g822_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4940), .Q (g_15381), .QN ());
DFFSRX1 g283_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4876), .Q (g_5450), .QN ());
MX2X1 g63126(.A (g3929), .B (n_4655), .S0 (n_9256), .Y (n_5300));
MX2X1 g63128(.A (g3937), .B (n_4654), .S0 (n_9750), .Y (n_5299));
DFFSRX1 g4372_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4887), .Q (g4372), .QN ());
MX2X1 g63143(.A (g1644), .B (n_4676), .S0 (n_9234), .Y (n_5297));
MX2X1 g63144(.A (g2606), .B (n_4645), .S0 (n_9167), .Y (n_5296));
MX2X1 g63145(.A (g1636), .B (n_4673), .S0 (n_10005), .Y (n_5294));
MX2X1 g63146(.A (g2599), .B (n_4640), .S0 (n_10005), .Y (n_5293));
NAND3X1 g60928(.A (n_4867), .B (n_2794), .C (n_4598), .Y (n_5291));
NOR2X1 g63203(.A (n_4898), .B (n_8588), .Y (n_5290));
NOR2X1 g63211(.A (n_4897), .B (n_10895), .Y (n_5289));
AOI21X1 g62050(.A0 (n_4590), .A1 (n_4251), .B0 (n_8707), .Y (n_5288));
INVX1 g63249(.A (n_6570), .Y (n_5287));
NAND4X1 g63316(.A (n_3219), .B (n_4605), .C (n_4098), .D (n_3895), .Y(n_5284));
AOI22X1 g60931(.A0 (n_4600), .A1 (n_9521), .B0 (n_10196), .B1(n_10952), .Y (n_5283));
MX2X1 g61177(.A (n_4529), .B (n_4603), .S0 (n_9894), .Y (n_5282));
MX2X1 g61184(.A (n_4531), .B (n_4597), .S0 (n_9234), .Y (n_5279));
MX2X1 g61190(.A (n_4726), .B (n_4594), .S0 (n_9172), .Y (n_5278));
NAND3X1 g62240(.A (n_4833), .B (n_2783), .C (n_4809), .Y (n_5276));
OAI22X1 g63645(.A0 (n_4049), .A1 (n_9193), .B0 (g4369), .B1 (n_9992),.Y (n_5275));
NAND2X1 g61212(.A (g4375), .B (n_9019), .Y (n_5273));
MX2X1 g62303(.A (g5046), .B (n_4813), .S0 (n_10063), .Y (n_5272));
MX2X1 g63757(.A (g_22371), .B (g14125), .S0 (n_5582), .Y (n_5271));
MX2X1 g62322(.A (n_11055), .B (n_4806), .S0 (n_9167), .Y (n_5270));
DFFSRX1 g4185_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4824), .Q (g11770), .QN ());
AOI21X1 g61262(.A0 (n_4836), .A1 (n_1528), .B0 (n_4838), .Y (n_5268));
AOI21X1 g61264(.A0 (n_4834), .A1 (n_1529), .B0 (n_4835), .Y (n_5267));
AOI21X1 g61265(.A0 (n_4829), .A1 (n_2258), .B0 (n_4830), .Y (n_5266));
DFFSRX1 g411_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4915), .Q (g_19113), .QN ());
AOI21X1 g61267(.A0 (n_4827), .A1 (n_1519), .B0 (n_4828), .Y (n_5265));
DFFSRX1 g5481_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4929), .Q (), .QN (g5481));
DFFSRX1 g5485_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4928), .Q (g5485), .QN ());
DFFSRX1 g5827_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4926), .Q (), .QN (g5827));
DFFSRX1 g5831_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4925), .Q (g5831), .QN ());
DFFSRX1 g1802_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4924), .Q (n_4139), .QN ());
DFFSRX1 g6177_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4922), .Q (g6177), .QN ());
DFFSRX1 g6173_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4923), .Q (), .QN (g6173));
DFFSRX1 g1906_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4918), .Q (g1906), .QN ());
DFFSRX1 g1936_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4917), .Q (g1936), .QN ());
DFFSRX1 g4112_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4877), .Q (), .QN (g4112));
DFFSRX1 g4116_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4870), .Q (), .QN (g4116));
DFFSRX1 g4119_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4869), .Q (), .QN (g4119));
DFFSRX1 g4122_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4868), .Q (), .QN (g4122));
DFFSRX1 g4005_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4891), .Q (g_3974), .QN ());
DFFSRX1 g5062_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4841), .Q (n_1356), .QN ());
OAI21X1 g64370(.A0 (n_4803), .A1 (n_10650), .B0 (n_4822), .Y(g33079));
OAI21X1 g64371(.A0 (n_4804), .A1 (n_10650), .B0 (n_4823), .Y(g33435));
DFFSRX1 g4531_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4934), .Q (), .QN (g4531));
NAND3X1 g61064(.A (n_4787), .B (n_10372), .C (n_10949), .Y (n_5259));
XOR2X1 g61289(.A (n_1261), .B (n_4798), .Y (n_5258));
NAND3X1 g61069(.A (n_4920), .B (n_10669), .C (n_9894), .Y (n_10548));
INVX1 g62616(.A (n_5374), .Y (n_5454));
NAND2X1 g62636(.A (n_4931), .B (n_4572), .Y (n_5254));
NAND3X1 g61072(.A (n_4919), .B (n_10978), .C (n_9209), .Y (n_5253));
OAI22X1 g62689(.A0 (n_4725), .A1 (n_9371), .B0 (g2667), .B1 (n_9992),.Y (n_5252));
MX2X1 g62690(.A (g2671), .B (n_4712), .S0 (n_8955), .Y (n_5251));
OAI22X1 g62693(.A0 (n_4730), .A1 (n_10952), .B0 (g1706), .B1(n_9992), .Y (n_5249));
MX2X1 g62698(.A (g1710), .B (n_4715), .S0 (n_9279), .Y (n_5248));
OR2X1 g64528(.A (n_5362), .B (n_9398), .Y (n_5247));
MX2X1 g62703(.A (g1816), .B (n_10467), .S0 (n_9172), .Y (n_5246));
OAI22X1 g62705(.A0 (n_4723), .A1 (n_9976), .B0 (g1840), .B1 (n_9992),.Y (n_5245));
MX2X1 g62706(.A (g1844), .B (n_4711), .S0 (n_9240), .Y (n_5244));
MX2X1 g62707(.A (g1950), .B (n_4731), .S0 (n_9172), .Y (n_5242));
OAI22X1 g62709(.A0 (n_4721), .A1 (n_9193), .B0 (g1974), .B1 (n_9992),.Y (n_5241));
MX2X1 g62710(.A (g1978), .B (n_4710), .S0 (n_8955), .Y (n_5240));
OAI22X1 g62713(.A0 (n_4719), .A1 (n_10952), .B0 (g2108), .B1(n_9830), .Y (n_5239));
MX2X1 g62714(.A (g2112), .B (n_4709), .S0 (n_9750), .Y (n_5238));
MX2X1 g62716(.A (n_5961), .B (n_4713), .S0 (n_9501), .Y (n_5236));
OAI22X1 g61331(.A0 (n_4783), .A1 (n_10952), .B0 (g1740), .B1(n_9651), .Y (n_5235));
MX2X1 g61332(.A (n_4190), .B (n_4782), .S0 (n_8955), .Y (n_5233));
OAI22X1 g62721(.A0 (n_4717), .A1 (n_9599), .B0 (g2399), .B1 (n_9992),.Y (n_5232));
OAI22X1 g62723(.A0 (n_4532), .A1 (n_9772), .B0 (g2509), .B1 (n_9558),.Y (n_5231));
MX2X1 g62724(.A (n_5229), .B (n_4520), .S0 (n_9311), .Y (n_5230));
NAND2X1 g64655(.A (n_4936), .B (n_11012), .Y (n_5227));
DFFSRX1 g1070_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4587), .Q (), .QN (g_6283));
MX2X1 g64698(.A (n_4556), .B (n_4232), .S0 (n_8895), .Y (n_5226));
DFFSRX1 g5077_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4746), .Q (), .QN (g5077));
MX2X1 g64705(.A (n_4555), .B (n_4230), .S0 (n_8895), .Y (n_5225));
AOI21X1 g64706(.A0 (n_4225), .A1 (n_8895), .B0 (n_4812), .Y (n_5224));
AND2X1 g60974(.A (n_4639), .B (n_4690), .Y (n_5223));
AND2X1 g60975(.A (n_4634), .B (n_4680), .Y (n_5222));
AND2X1 g62821(.A (g4438), .B (n_10687), .Y (n_5364));
NAND2X1 g62822(.A (g4438), .B (n_9107), .Y (n_5221));
AND2X1 g60976(.A (n_4630), .B (n_4678), .Y (n_5219));
AND2X1 g60977(.A (n_4619), .B (n_4677), .Y (n_5218));
AOI21X1 g62921(.A0 (g5069), .A1 (g5084), .B0 (n_4753), .Y (n_5215));
DFFSRX1 g1024_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4589), .Q (g_22306), .QN ());
DFFSRX1 g6181_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4789), .Q (), .QN (g6181));
MX2X1 g62944(.A (g5188), .B (n_4442), .S0 (n_9469), .Y (n_5214));
MX2X1 g62945(.A (g5204), .B (n_4441), .S0 (n_8955), .Y (n_5213));
MX2X1 g62946(.A (g5256), .B (n_4440), .S0 (n_9000), .Y (n_5212));
MX2X1 g62947(.A (g5212), .B (n_4439), .S0 (n_9256), .Y (n_5210));
MX2X1 g62948(.A (g5260), .B (n_4347), .S0 (n_9311), .Y (n_5209));
MX2X1 g62949(.A (g5220), .B (n_4493), .S0 (n_9172), .Y (n_5207));
MX2X1 g62950(.A (g5264), .B (n_4438), .S0 (n_9000), .Y (n_5206));
MX2X1 g62951(.A (g5196), .B (n_4437), .S0 (n_8955), .Y (n_5205));
MX2X1 g62952(.A (g5200), .B (n_4458), .S0 (n_9091), .Y (n_5204));
MX2X1 g62953(.A (g5208), .B (n_4459), .S0 (n_9240), .Y (n_5202));
MX2X1 g62955(.A (g5224), .B (n_4381), .S0 (n_9000), .Y (n_5201));
MX2X1 g62956(.A (g5228), .B (n_4507), .S0 (n_9156), .Y (n_5200));
MX2X1 g62957(.A (g5232), .B (n_4504), .S0 (n_9167), .Y (n_5199));
MX2X1 g62959(.A (g5240), .B (n_4503), .S0 (n_9256), .Y (n_5197));
MX2X1 g62962(.A (g5252), .B (n_4400), .S0 (n_8955), .Y (n_5195));
MX2X1 g62963(.A (g5268), .B (n_4434), .S0 (n_9256), .Y (n_5193));
MX2X1 g62967(.A (g5535), .B (n_4433), .S0 (n_9091), .Y (n_5192));
MX2X1 g62968(.A (g5551), .B (n_4432), .S0 (n_9797), .Y (n_5190));
MX2X1 g62969(.A (g5603), .B (n_4431), .S0 (n_9359), .Y (n_5189));
MX2X1 g62970(.A (g5559), .B (n_4345), .S0 (n_10687), .Y (n_5187));
MX2X1 g62971(.A (g5607), .B (n_4430), .S0 (n_9172), .Y (n_5186));
MX2X1 g62972(.A (g5567), .B (n_4502), .S0 (n_9240), .Y (n_5185));
MX2X1 g62973(.A (g5611), .B (n_4429), .S0 (n_10005), .Y (n_5184));
MX2X1 g62974(.A (g5543), .B (n_4428), .S0 (n_9834), .Y (n_5183));
MX2X1 g62975(.A (g5547), .B (n_4501), .S0 (n_9311), .Y (n_5182));
MX2X1 g62976(.A (g5555), .B (n_4500), .S0 (n_9000), .Y (n_5181));
MX2X1 g62978(.A (g5571), .B (n_4427), .S0 (n_9992), .Y (n_5179));
MX2X1 g62979(.A (g5575), .B (n_4498), .S0 (n_9797), .Y (n_5177));
MX2X1 g62980(.A (g5579), .B (n_4496), .S0 (n_8955), .Y (n_5175));
MX2X1 g62982(.A (g5587), .B (n_4495), .S0 (n_8955), .Y (n_5174));
MX2X1 g62983(.A (g5591), .B (n_4426), .S0 (n_8955), .Y (n_5173));
MX2X1 g62984(.A (g5595), .B (n_4425), .S0 (n_9000), .Y (n_5172));
MX2X1 g62985(.A (g5599), .B (n_4423), .S0 (n_9992), .Y (n_5171));
MX2X1 g62986(.A (g5615), .B (n_4421), .S0 (n_8955), .Y (n_5170));
MX2X1 g62992(.A (g5881), .B (n_4420), .S0 (n_9466), .Y (n_5168));
MX2X1 g62993(.A (g5897), .B (n_4419), .S0 (n_9834), .Y (n_5167));
MX2X1 g62994(.A (g5949), .B (n_4418), .S0 (n_9156), .Y (n_5165));
MX2X1 g62995(.A (g5905), .B (n_4417), .S0 (n_9167), .Y (n_5164));
MX2X1 g62996(.A (g5953), .B (n_4416), .S0 (n_9156), .Y (n_5163));
MX2X1 g62997(.A (g5913), .B (n_4492), .S0 (n_9000), .Y (n_5161));
MX2X1 g62998(.A (g5957), .B (n_4415), .S0 (n_9359), .Y (n_5160));
MX2X1 g62999(.A (g5889), .B (n_4414), .S0 (n_9000), .Y (n_5159));
MX2X1 g63000(.A (g5893), .B (n_4490), .S0 (n_9992), .Y (n_5158));
MX2X1 g63001(.A (g5901), .B (n_4489), .S0 (n_9156), .Y (n_5156));
MX2X1 g63003(.A (g5917), .B (n_4413), .S0 (n_9311), .Y (n_5155));
MX2X1 g63004(.A (g5921), .B (n_4488), .S0 (n_9218), .Y (n_5154));
MX2X1 g63005(.A (g5925), .B (n_4487), .S0 (n_8955), .Y (n_5152));
MX2X1 g63006(.A (g5929), .B (n_4411), .S0 (n_9000), .Y (n_5151));
MX2X1 g63007(.A (g5933), .B (n_4486), .S0 (n_9359), .Y (n_5150));
MX2X1 g63008(.A (g5937), .B (n_4403), .S0 (n_9172), .Y (n_5149));
MX2X1 g63010(.A (g5945), .B (n_4410), .S0 (n_9797), .Y (n_5148));
MX2X1 g63011(.A (g5961), .B (n_4409), .S0 (n_9992), .Y (n_5146));
MX2X1 g63015(.A (g3119), .B (n_4485), .S0 (n_9664), .Y (n_5144));
MX2X1 g63017(.A (g6227), .B (n_4436), .S0 (n_9172), .Y (n_5143));
MX2X1 g63018(.A (g6243), .B (n_4360), .S0 (n_9358), .Y (n_5141));
MX2X1 g63020(.A (g6295), .B (n_4408), .S0 (n_9091), .Y (n_5139));
MX2X1 g63021(.A (g6251), .B (n_4407), .S0 (n_8955), .Y (n_5137));
MX2X1 g63022(.A (g6299), .B (n_4406), .S0 (n_9333), .Y (n_5136));
MX2X1 g63023(.A (g6259), .B (n_4483), .S0 (n_9000), .Y (n_5135));
MX2X1 g63024(.A (g6303), .B (n_4405), .S0 (n_9234), .Y (n_5134));
MX2X1 g63025(.A (g6235), .B (n_4404), .S0 (n_9311), .Y (n_5133));
MX2X1 g63026(.A (g6239), .B (n_4481), .S0 (n_9681), .Y (n_5131));
MX2X1 g63027(.A (g6247), .B (n_4479), .S0 (n_9681), .Y (n_5130));
MX2X1 g63029(.A (g6263), .B (n_4402), .S0 (n_9333), .Y (n_5129));
MX2X1 g63030(.A (g6267), .B (n_4478), .S0 (n_9240), .Y (n_5128));
MX2X1 g63031(.A (g6271), .B (n_4477), .S0 (n_9894), .Y (n_5127));
MX2X1 g63032(.A (g6275), .B (n_4401), .S0 (n_9797), .Y (n_5126));
MX2X1 g63033(.A (g6279), .B (n_4450), .S0 (n_9797), .Y (n_5125));
MX2X1 g63037(.A (g6307), .B (n_4399), .S0 (n_9311), .Y (n_5124));
MX2X1 g63038(.A (g3179), .B (n_4398), .S0 (n_9256), .Y (n_5123));
MX2X1 g63039(.A (g3195), .B (n_4397), .S0 (n_9234), .Y (n_5122));
MX2X1 g63040(.A (g3247), .B (n_4396), .S0 (n_9234), .Y (n_5121));
MX2X1 g63041(.A (g3203), .B (n_4395), .S0 (n_9156), .Y (n_5119));
MX2X1 g63042(.A (g3251), .B (n_4393), .S0 (n_9000), .Y (n_5118));
MX2X1 g63043(.A (g3211), .B (n_4475), .S0 (n_9000), .Y (n_5116));
MX2X1 g63044(.A (g3255), .B (n_4394), .S0 (n_9172), .Y (n_5115));
MX2X1 g63045(.A (g3187), .B (n_4392), .S0 (n_9172), .Y (n_5113));
MX2X1 g63048(.A (g3191), .B (n_4474), .S0 (n_10687), .Y (n_5112));
DFFSRX1 g5835_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4796), .Q (), .QN (g5835));
MX2X1 g63050(.A (g3199), .B (n_4473), .S0 (n_9000), .Y (n_5111));
MX2X1 g63051(.A (g3207), .B (n_4391), .S0 (n_9000), .Y (n_5110));
MX2X1 g63052(.A (g3215), .B (n_4390), .S0 (n_9000), .Y (n_5109));
MX2X1 g63053(.A (g3219), .B (n_4472), .S0 (n_10005), .Y (n_5107));
MX2X1 g63054(.A (g6573), .B (n_4388), .S0 (n_9139), .Y (n_5106));
MX2X1 g63055(.A (g3223), .B (n_4471), .S0 (n_9311), .Y (n_5104));
MX2X1 g63056(.A (g6589), .B (n_4346), .S0 (n_9256), .Y (n_5103));
MX2X1 g63057(.A (g3227), .B (n_4387), .S0 (n_9091), .Y (n_5101));
MX2X1 g63058(.A (g6641), .B (n_4366), .S0 (n_9797), .Y (n_5100));
MX2X1 g63059(.A (g6597), .B (n_4389), .S0 (n_8955), .Y (n_5098));
MX2X1 g63060(.A (g3231), .B (n_4469), .S0 (n_9172), .Y (n_5097));
MX2X1 g63061(.A (g6645), .B (n_4363), .S0 (n_9359), .Y (n_5095));
MX2X1 g63062(.A (g6605), .B (n_4468), .S0 (n_9359), .Y (n_5094));
MX2X1 g63063(.A (g6649), .B (n_4349), .S0 (n_8955), .Y (n_5093));
MX2X1 g63064(.A (g6581), .B (n_4369), .S0 (n_8955), .Y (n_5092));
MX2X1 g63065(.A (g3235), .B (n_4380), .S0 (n_8955), .Y (n_5091));
MX2X1 g63066(.A (g6585), .B (n_4470), .S0 (n_8955), .Y (n_5090));
MX2X1 g63067(.A (g6593), .B (n_4446), .S0 (n_9172), .Y (n_5088));
MX2X1 g63068(.A (g3239), .B (n_4386), .S0 (n_9218), .Y (n_5087));
MX2X1 g63069(.A (g6601), .B (n_4412), .S0 (n_10005), .Y (n_5086));
MX2X1 g63070(.A (g3243), .B (n_4385), .S0 (n_9256), .Y (n_5085));
MX2X1 g63071(.A (g6609), .B (n_4344), .S0 (n_9000), .Y (n_5084));
MX2X1 g63072(.A (g6613), .B (n_4449), .S0 (n_9894), .Y (n_5083));
MX2X1 g63073(.A (g3259), .B (n_4348), .S0 (n_9234), .Y (n_5082));
MX2X1 g63074(.A (g6617), .B (n_4451), .S0 (n_9978), .Y (n_5081));
MX2X1 g63076(.A (g6625), .B (n_4467), .S0 (n_9218), .Y (n_5079));
MX2X1 g63078(.A (g6633), .B (n_4384), .S0 (n_8955), .Y (n_5077));
MX2X1 g63079(.A (g6637), .B (n_4383), .S0 (n_8955), .Y (n_5076));
MX2X1 g63080(.A (g6653), .B (n_4382), .S0 (n_9797), .Y (n_5075));
MX2X1 g63087(.A (g3530), .B (n_4379), .S0 (n_9466), .Y (n_5073));
MX2X1 g63088(.A (g3546), .B (n_4378), .S0 (n_8955), .Y (n_5072));
MX2X1 g63089(.A (g3598), .B (n_4377), .S0 (n_9311), .Y (n_5071));
MX2X1 g63090(.A (g3554), .B (n_4376), .S0 (n_9311), .Y (n_5069));
MX2X1 g61418(.A (g2004), .B (n_5057), .S0 (n_4306), .Y (n_5068));
MX2X1 g63091(.A (g3602), .B (n_4375), .S0 (n_9167), .Y (n_5067));
MX2X1 g63092(.A (g3562), .B (n_4466), .S0 (n_9750), .Y (n_5065));
MX2X1 g63093(.A (g3606), .B (n_4374), .S0 (n_9234), .Y (n_5064));
MX2X1 g63094(.A (g3538), .B (n_4373), .S0 (n_9750), .Y (n_5063));
MX2X1 g63095(.A (g3542), .B (n_4465), .S0 (n_9218), .Y (n_5062));
MX2X1 g63096(.A (g3550), .B (n_4464), .S0 (n_9359), .Y (n_5060));
MX2X1 g63097(.A (g3558), .B (n_4372), .S0 (n_9359), .Y (n_5059));
MX2X1 g61421(.A (g2016), .B (n_5057), .S0 (n_4305), .Y (n_5058));
MX2X1 g63098(.A (g3566), .B (n_4371), .S0 (n_8955), .Y (n_5056));
MX2X1 g63099(.A (g3570), .B (n_4462), .S0 (n_8955), .Y (n_5055));
MX2X1 g63100(.A (g3574), .B (n_4461), .S0 (n_9156), .Y (n_5053));
MX2X1 g63101(.A (g3578), .B (n_4370), .S0 (n_9156), .Y (n_5052));
MX2X1 g63102(.A (g3582), .B (n_4460), .S0 (n_9311), .Y (n_5051));
MX2X1 g63103(.A (g3586), .B (n_4368), .S0 (n_9172), .Y (n_5050));
MX2X1 g63104(.A (g3590), .B (n_4367), .S0 (n_9234), .Y (n_5048));
MX2X1 g63105(.A (g3594), .B (n_4365), .S0 (n_9311), .Y (n_5047));
MX2X1 g63106(.A (g3610), .B (n_4364), .S0 (n_9000), .Y (n_5046));
MX2X1 g61422(.A (g2020), .B (n_5057), .S0 (n_4319), .Y (n_5045));
MX2X1 g61423(.A (g2024), .B (n_5057), .S0 (n_4303), .Y (n_5044));
MX2X1 g63112(.A (g3881), .B (n_4362), .S0 (n_9553), .Y (n_5043));
MX2X1 g63113(.A (g3897), .B (n_4361), .S0 (n_9000), .Y (n_5042));
MX2X1 g63114(.A (g3949), .B (n_4359), .S0 (n_9750), .Y (n_5041));
MX2X1 g63115(.A (g3905), .B (n_4358), .S0 (n_9000), .Y (n_5040));
AOI21X1 g61424(.A0 (n_4742), .A1 (n_1532), .B0 (n_4744), .Y (n_5039));
MX2X1 g63116(.A (g3953), .B (n_4357), .S0 (n_9240), .Y (n_5038));
MX2X1 g63117(.A (g3913), .B (n_4457), .S0 (n_9553), .Y (n_5037));
MX2X1 g63118(.A (g3957), .B (n_4356), .S0 (n_10687), .Y (n_5035));
MX2X1 g63119(.A (g3889), .B (n_4355), .S0 (n_9311), .Y (n_5034));
MX2X1 g63120(.A (g3893), .B (n_4456), .S0 (n_9000), .Y (n_5033));
MX2X1 g63121(.A (g3901), .B (n_4455), .S0 (n_9000), .Y (n_5032));
AOI21X1 g61426(.A0 (n_4740), .A1 (n_1533), .B0 (n_4741), .Y (n_5030));
MX2X1 g63122(.A (g3909), .B (n_4354), .S0 (n_9000), .Y (n_5029));
MX2X1 g63123(.A (g3917), .B (n_4353), .S0 (n_9359), .Y (n_5028));
MX2X1 g63124(.A (g3921), .B (n_4454), .S0 (n_9000), .Y (n_5026));
MX2X1 g63125(.A (g3925), .B (n_4453), .S0 (n_9000), .Y (n_5025));
MX2X1 g63127(.A (g3933), .B (n_4452), .S0 (n_10005), .Y (n_5024));
MX2X1 g63129(.A (g3941), .B (n_4352), .S0 (n_9750), .Y (n_5023));
AOI21X1 g61428(.A0 (n_4738), .A1 (n_2521), .B0 (n_4739), .Y (n_5022));
MX2X1 g63130(.A (g3945), .B (n_4351), .S0 (n_9091), .Y (n_5021));
MX2X1 g63131(.A (g3961), .B (n_4350), .S0 (n_8955), .Y (n_5020));
AOI21X1 g61430(.A0 (n_4736), .A1 (n_1510), .B0 (n_4737), .Y (n_5019));
MX2X1 g63136(.A (g2338), .B (n_4336), .S0 (n_8955), .Y (n_5018));
MX2X1 g63137(.A (g2331), .B (n_4333), .S0 (n_9240), .Y (n_5017));
MX2X1 g63139(.A (g3470), .B (n_4448), .S0 (n_9091), .Y (n_5016));
MX2X1 g63140(.A (g2472), .B (n_4343), .S0 (n_9000), .Y (n_5015));
MX2X1 g63141(.A (g2465), .B (n_4340), .S0 (n_9000), .Y (n_5014));
NAND2X1 g63205(.A (n_4445), .B (n_4700), .Y (n_5013));
NAND2X1 g63215(.A (n_4444), .B (n_4695), .Y (n_5012));
NAND2X1 g62053(.A (n_3774), .B (n_4642), .Y (n_5009));
AOI22X1 g63248(.A0 (n_4330), .A1 (n_2943), .B0 (n_2944), .B1(n_5007), .Y (n_5008));
AOI22X1 g63252(.A0 (n_4328), .A1 (n_2940), .B0 (n_2941), .B1(n_5007), .Y (n_5006));
AOI22X1 g63254(.A0 (n_4325), .A1 (n_2936), .B0 (n_2937), .B1(n_5007), .Y (n_5005));
AOI22X1 g63256(.A0 (n_4317), .A1 (n_3253), .B0 (n_2933), .B1(n_5007), .Y (n_5004));
AOI22X1 g63258(.A0 (n_4323), .A1 (n_2930), .B0 (n_2931), .B1(n_5007), .Y (n_5003));
AOI22X1 g63263(.A0 (n_4321), .A1 (n_2928), .B0 (n_2929), .B1(n_5007), .Y (n_5002));
AOI22X1 g63264(.A0 (n_4315), .A1 (n_2923), .B0 (n_2924), .B1(n_5007), .Y (n_5001));
NAND4X1 g60930(.A (n_4593), .B (n_4866), .C (n_9750), .D (n_263), .Y(n_5000));
AOI21X1 g62082(.A0 (g_5450), .A1 (n_9856), .B0 (n_4672), .Y (n_4999));
NAND4X1 g63297(.A (n_6973), .B (n_10897), .C (g16722), .D (g3598), .Y(n_4996));
NAND3X1 g63325(.A (n_4693), .B (g_22379), .C (n_9351), .Y (n_4991));
DFFSRX1 g4031_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16748), .Q (g4031), .QN ());
NAND3X1 g63461(.A (n_4616), .B (n_2973), .C (g5156), .Y (n_4990));
NAND3X1 g63492(.A (n_868), .B (n_4293), .C (n_9874), .Y (n_4987));
AOI21X1 g60936(.A0 (n_4575), .A1 (n_2309), .B0 (n_9193), .Y (n_4986));
AOI22X1 g63553(.A0 (n_688), .A1 (n_4293), .B0 (n_4885), .B1 (g3831),.Y (n_4985));
NAND4X1 g63561(.A (n_6787), .B (g3933), .C (g13906), .D (n_5402), .Y(n_4984));
OAI21X1 g62213(.A0 (n_4567), .A1 (n_4982), .B0 (n_1283), .Y (n_4983));
OAI21X1 g62214(.A0 (n_4566), .A1 (n_4980), .B0 (n_1561), .Y (n_4981));
OAI21X1 g62215(.A0 (n_4565), .A1 (n_4978), .B0 (n_1282), .Y (n_4979));
OAI21X1 g62217(.A0 (n_4564), .A1 (n_11070), .B0 (n_1560), .Y(n_4977));
NAND4X1 g61553(.A (n_4581), .B (n_4843), .C (n_10013), .D (g4616), .Y(n_4976));
NAND2X1 g60939(.A (n_4586), .B (n_4243), .Y (n_4975));
NAND4X1 g62268(.A (n_4811), .B (n_4832), .C (n_9279), .D (n_287), .Y(n_4974));
OAI22X1 g61592(.A0 (n_4939), .A1 (n_4579), .B0 (n_79), .B1 (n_9862),.Y (n_4972));
XOR2X1 g63769(.A (n_2692), .B (n_4293), .Y (n_4971));
MX2X1 g63804(.A (g_21318), .B (n_4288), .S0 (n_9000), .Y (n_4970));
DFFSRX1 g884_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14125), .Q (g14147), .QN ());
OR2X1 g61258(.A (n_4968), .B (g1682), .Y (n_4969));
DFFSRX1 g1367_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4684), .Q (g1367), .QN ());
DFFSRX1 g1542_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4591), .Q (g1542), .QN ());
DFFSRX1 g1312_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4821), .Q (g1312), .QN ());
DFFSRX1 g1233_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4794), .Q (g10500), .QN ());
DFFSRX1 g4950_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4626), .Q (g4950), .QN ());
DFFSRX1 g4939_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4627), .Q (g4939), .QN ());
DFFSRX1 g6527_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4785), .Q (), .QN (g6527));
DFFSRX1 g4593_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4706), .Q (g4593), .QN ());
DFFSRX1 g4332_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4714), .Q (g4332), .QN ());
DFFSRX1 g812_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4663), .Q (g_10715), .QN ());
DFFSRX1 g4049_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4585), .Q (g4049), .QN ());
AOI21X1 g61266(.A0 (n_4583), .A1 (n_919), .B0 (n_4584), .Y (n_4967));
DFFSRX1 g5134_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4800), .Q (), .QN (g5134));
DFFSRX1 g5138_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4799), .Q (g5138), .QN ());
DFFSRX1 g5489_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4797), .Q (), .QN (g5489));
DFFSRX1 g6523_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4786), .Q (g6523), .QN ());
DFFSRX1 g3639_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4734), .Q (g3639), .QN ());
DFFSRX1 g3990_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4732), .Q (g3990), .QN ());
DFFSRX1 g5471_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4752), .Q (g5471), .QN ());
DFFSRX1 g5817_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4751), .Q (g5817), .QN ());
DFFSRX1 g6163_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4750), .Q (g6163), .QN ());
DFFSRX1 g3288_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4735), .Q (g3288), .QN ());
DFFSRX1 g3352_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4705), .Q (n_7004), .QN ());
DFFSRX1 g3703_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4704), .Q (n_6979), .QN ());
DFFSRX1 g5046_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4747), .Q (g5046), .QN ());
DFFSRX1 g255_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4636), .Q (g_21318), .QN ());
DFFSRX1 g3050_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4624), .Q (g3050), .QN ());
DFFSRX1 g6098_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4623), .Q (g6098), .QN ());
DFFSRX1 g6444_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4622), .Q (g6444), .QN ());
DFFSRX1 g3401_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4620), .Q (g3401), .QN ());
DFFSRX1 g3752_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4621), .Q (g3752), .QN ());
DFFSRX1 g5752_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4625), .Q (g5752), .QN ());
AOI21X1 g62254(.A0 (n_4262), .A1 (n_1972), .B0 (g4369), .Y (g34839));
AND2X1 g61063(.A (n_4766), .B (n_4795), .Y (n_4966));
XOR2X1 g61287(.A (n_1260), .B (n_4559), .Y (n_4965));
OR2X1 g62584(.A (n_4963), .B (n_3654), .Y (n_4964));
XOR2X1 g61290(.A (n_1257), .B (n_4562), .Y (n_4962));
NAND4X1 g62600(.A (n_4815), .B (g_4449), .C (n_10013), .D (n_3914),.Y (n_4961));
AND2X1 g61067(.A (n_4763), .B (n_4792), .Y (n_4960));
AND2X1 g61068(.A (n_4759), .B (n_4790), .Y (n_4959));
OR4X1 g62617(.A (g4438), .B (g4452), .C (g4443), .D (n_334), .Y(n_5374));
OAI22X1 g61744(.A0 (n_4519), .A1 (n_4956), .B0 (n_512), .B1 (n_9992),.Y (n_4957));
OR4X1 g62628(.A (n_2756), .B (n_11189), .C (n_11188), .D (n_4205), .Y(n_5457));
XOR2X1 g61745(.A (g4608), .B (n_4554), .Y (n_4955));
AND2X1 g61070(.A (n_4756), .B (n_4788), .Y (n_4954));
NAND3X1 g61071(.A (n_4784), .B (n_10853), .C (n_9834), .Y (n_4953));
MX2X1 g62687(.A (n_4893), .B (n_4528), .S0 (n_9000), .Y (n_4952));
MX2X1 g62688(.A (n_5958), .B (n_4526), .S0 (n_9333), .Y (n_4951));
MX2X1 g62692(.A (n_5964), .B (n_4525), .S0 (n_9172), .Y (n_4950));
MX2X1 g62704(.A (n_4948), .B (n_4524), .S0 (n_9172), .Y (n_4949));
MX2X1 g62708(.A (n_4946), .B (n_4523), .S0 (n_9156), .Y (n_4947));
MX2X1 g62712(.A (n_5953), .B (n_4522), .S0 (n_9218), .Y (n_4945));
OAI22X1 g62719(.A0 (n_4530), .A1 (n_9976), .B0 (g2375), .B1 (n_9862),.Y (n_4944));
MX2X1 g62720(.A (n_4942), .B (n_4521), .S0 (n_9553), .Y (n_4943));
OAI22X1 g61841(.A0 (n_4939), .A1 (n_4155), .B0 (n_126), .B1 (n_9651),.Y (n_4940));
DFFSRX1 g736_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g11678), .Q (g_15127), .QN ());
INVX1 g64835(.A (n_4936), .Y (n_5362));
AOI21X1 g64852(.A0 (n_4223), .A1 (n_4032), .B0 (n_8895), .Y (n_4935));
NAND2X1 g62846(.A (n_4546), .B (n_3214), .Y (n_4934));
AOI21X1 g62932(.A0 (g5052), .A1 (n_10078), .B0 (n_4545), .Y (n_4931));
AOI21X1 g61275(.A0 (n_4273), .A1 (n_1713), .B0 (n_4274), .Y (n_4930));
MX2X1 g62964(.A (g5475), .B (n_4163), .S0 (n_9311), .Y (n_4929));
OAI22X1 g62965(.A0 (n_10346), .A1 (n_9599), .B0 (g5481), .B1(n_9992), .Y (n_4928));
MX2X1 g62987(.A (g1779), .B (n_4142), .S0 (n_9000), .Y (n_4927));
MX2X1 g62988(.A (g5821), .B (n_4161), .S0 (n_9091), .Y (n_4926));
OAI22X1 g62989(.A0 (n_4165), .A1 (n_9371), .B0 (g5827), .B1 (n_9698),.Y (n_4925));
MX2X1 g62991(.A (g1772), .B (n_4140), .S0 (n_9311), .Y (n_4924));
MX2X1 g63012(.A (g6167), .B (n_4160), .S0 (n_9664), .Y (n_4923));
OAI22X1 g63013(.A0 (n_10448), .A1 (n_9599), .B0 (g6173), .B1(n_9992), .Y (n_4922));
NAND4X1 g61941(.A (n_3913), .B (n_11079), .C (n_9139), .D (n_284), .Y(n_4921));
XOR2X1 g61139(.A (n_963), .B (n_4150), .Y (n_4920));
XOR2X1 g61141(.A (n_942), .B (n_4151), .Y (n_4919));
MX2X1 g63081(.A (g1913), .B (n_4147), .S0 (n_9992), .Y (n_4918));
MX2X1 g63082(.A (g1906), .B (n_4145), .S0 (n_9834), .Y (n_4917));
MX2X1 g61982(.A (n_640), .B (n_4152), .S0 (n_9167), .Y (n_4915));
AOI21X1 g61429(.A0 (n_4539), .A1 (n_928), .B0 (n_4540), .Y (n_4913));
NAND2X1 g62019(.A (n_4422), .B (g_16404), .Y (n_4912));
NAND4X1 g62023(.A (n_4576), .B (n_4671), .C (n_9209), .D (g_19659),.Y (n_4911));
AOI22X1 g63265(.A0 (n_917), .A1 (n_10378), .B0 (n_10099), .B1(n_4906), .Y (n_4907));
OAI21X1 g63299(.A0 (n_702), .A1 (n_6752), .B0 (n_4184), .Y (n_4905));
AOI21X1 g63300(.A0 (n_10099), .A1 (g2269), .B0 (n_4514), .Y (n_4904));
AOI22X1 g63323(.A0 (n_783), .A1 (n_4108), .B0 (n_4121), .B1 (g1592),.Y (n_4900));
OAI21X1 g63328(.A0 (n_10097), .A1 (n_6025), .B0 (n_4513), .Y(n_4899));
INVX1 g63399(.A (g3329), .Y (n_4898));
INVX1 g63403(.A (g3680), .Y (n_4897));
DFFSRX1 g482_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4553), .Q (g_16475), .QN ());
AND2X1 g63431(.A (n_4615), .B (g5156), .Y (n_4896));
AOI21X1 g63525(.A0 (g13966), .A1 (n_491), .B0 (n_4302), .Y (n_4891));
NAND3X1 g63530(.A (n_4313), .B (g_21806), .C (n_9398), .Y (n_4889));
NAND3X1 g60938(.A (n_4592), .B (g1379), .C (n_9894), .Y (n_4888));
DFFSRX1 g6509_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4547), .Q (g6509), .QN ());
OR2X1 g62239(.A (n_4286), .B (n_4068), .Y (n_4887));
MX2X1 g63616(.A (g3821), .B (n_85), .S0 (n_4885), .Y (n_4886));
MX2X1 g63624(.A (g2197), .B (g2153), .S0 (n_10378), .Y (n_4884));
MX2X1 g63625(.A (g2227), .B (g2197), .S0 (n_10378), .Y (n_4881));
AOI22X1 g63641(.A0 (n_3596), .A1 (n_9461), .B0 (n_4885), .B1(n_4878), .Y (n_4879));
OAI22X1 g63642(.A0 (n_4087), .A1 (n_9772), .B0 (n_3896), .B1(n_9992), .Y (n_4877));
DFFSRX1 g3303_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4512), .Q (g_4050), .QN ());
OAI22X1 g62291(.A0 (n_2567), .A1 (n_5723), .B0 (n_21), .B1 (n_9862),.Y (n_4876));
NAND4X1 g61590(.A (g_15380), .B (n_9992), .C (n_1124), .D (n_4578),.Y (n_4875));
XOR2X1 g62302(.A (g4045), .B (g3990), .Y (n_4874));
OAI22X1 g63794(.A0 (n_4086), .A1 (n_9431), .B0 (g4112), .B1 (n_9521),.Y (n_4870));
OAI22X1 g63795(.A0 (n_4085), .A1 (n_9269), .B0 (g4116), .B1(n_10005), .Y (n_4869));
OAI22X1 g63796(.A0 (n_4084), .A1 (n_9599), .B0 (g4119), .B1 (n_9862),.Y (n_4868));
DFFSRX1 g1018_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4577), .Q (g_16958), .QN ());
NAND4X1 g60945(.A (n_4569), .B (n_4866), .C (n_9359), .D (n_406), .Y(n_4867));
DFFSRX1 g4375_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4283), .Q (g4375), .QN ());
DFFSRX1 g1361_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4298), .Q (g1361), .QN ());
DFFSRX1 g1351_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4573), .Q (g1351), .QN ());
OAI21X1 g61263(.A0 (n_10761), .A1 (n_10097), .B0 (n_4515), .Y(n_4865));
NAND3X1 g64008(.A (n_10373), .B (n_916), .C (n_9894), .Y (n_4864));
DFFSRX1 g6519_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4557), .Q (), .QN (g6519));
DFFSRX1 g6682_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4533), .Q (n_11071), .QN ());
DFFSRX1 g5142_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4561), .Q (), .QN (g5142));
DFFSRX1 g854_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4506), .Q (), .QN (g_22639));
DFFSRX1 g1171_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4290), .Q (g1171), .QN ());
DFFSRX1 g2941_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4574), .Q (g2941), .QN ());
AOI21X1 g61269(.A0 (n_4281), .A1 (n_1702), .B0 (n_4282), .Y (n_4861));
DFFSRX1 g5041_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4563), .Q (g5041), .QN ());
DFFSRX1 g5297_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4538), .Q (g5297), .QN ());
DFFSRX1 g5644_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4537), .Q (g5644), .QN ());
DFFSRX1 g6336_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4534), .Q (g6336), .QN ());
DFFSRX1 g5990_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4535), .Q (g5990), .QN ());
DFFSRX1 g5124_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4550), .Q (g5124), .QN ());
AOI21X1 g61271(.A0 (n_4279), .A1 (n_1703), .B0 (n_4280), .Y (n_4860));
DFFSRX1 g4054_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4518), .Q (g4054), .QN ());
DFFSRX1 g703_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4338), .Q (n_1285), .QN ());
DFFSRX1 g3654_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4510), .Q (g_9298), .QN ());
DFFSRX1 g2886_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4508), .Q (g2886), .QN ());
DFFSRX1 g5406_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4331), .Q (g5406), .QN ());
DFFSRX1 g5022_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4297), .Q (n_6967), .QN ());
AOI21X1 g61272(.A0 (n_4277), .A1 (n_2293), .B0 (n_4278), .Y (n_4859));
MX2X1 g61273(.A (g2311), .B (n_8761), .S0 (n_4125), .Y (n_4858));
MX2X1 g64090(.A (g_22600), .B (g14096), .S0 (n_5582), .Y (n_4857));
AOI21X1 g61274(.A0 (n_4275), .A1 (n_1677), .B0 (n_4276), .Y (n_4856));
AOI21X1 g64083(.A0 (g2902), .A1 (g2907), .B0 (n_4291), .Y (g32185));
AOI21X1 g61277(.A0 (n_4271), .A1 (n_1714), .B0 (n_4272), .Y (n_4854));
AOI21X1 g61278(.A0 (n_4269), .A1 (n_2780), .B0 (n_4270), .Y (n_4853));
MX2X1 g61279(.A (g2445), .B (n_8763), .S0 (n_4123), .Y (n_4852));
AOI21X1 g61280(.A0 (n_4267), .A1 (n_1671), .B0 (n_4268), .Y (n_4851));
MX2X1 g61281(.A (g2563), .B (n_11190), .S0 (n_4117), .Y (n_4850));
MX2X1 g61283(.A (g2571), .B (n_11190), .S0 (n_6746), .Y (n_4849));
MX2X1 g61284(.A (g2575), .B (n_11190), .S0 (n_4113), .Y (n_4847));
MX2X1 g61285(.A (g2579), .B (n_11191), .S0 (n_4119), .Y (n_4846));
MX2X1 g61286(.A (g2583), .B (n_11191), .S0 (n_4111), .Y (n_4845));
NAND3X1 g61729(.A (n_2582), .B (n_4843), .C (n_8757), .Y (n_4844));
DFFSRX1 g4584_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4570), .Q (g4584), .QN ());
NAND3X1 g62601(.A (n_4810), .B (g_12465), .C (n_9698), .Y (n_4842));
NAND3X1 g64355(.A (n_4080), .B (n_4255), .C (n_2590), .Y (n_4841));
NOR2X1 g62622(.A (n_4839), .B (n_8879), .Y (n_4840));
NOR2X1 g61310(.A (n_10761), .B (n_4836), .Y (n_4838));
NOR2X1 g61311(.A (n_10761), .B (n_4834), .Y (n_4835));
NAND4X1 g62670(.A (n_4542), .B (n_4832), .C (n_9359), .D (n_251), .Y(n_4833));
NOR2X1 g61312(.A (n_10761), .B (n_4829), .Y (n_4830));
NOR2X1 g61314(.A (n_10761), .B (n_4827), .Y (n_4828));
MX2X1 g64453(.A (n_10867), .B (n_4248), .S0 (n_9359), .Y (n_4824));
DFFSRX1 g311_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4560), .Q (), .QN (g_16983));
OAI21X1 g64505(.A0 (n_4235), .A1 (n_4042), .B0 (n_10650), .Y(n_4823));
OAI21X1 g64506(.A0 (n_4239), .A1 (n_4043), .B0 (n_10650), .Y(n_4822));
NOR2X1 g60972(.A (n_4180), .B (n_9976), .Y (n_4821));
NAND4X1 g61826(.A (n_1787), .B (n_4045), .C (n_9874), .D (g_14342),.Y (n_4820));
NAND2X1 g62789(.A (n_11079), .B (n_9521), .Y (n_4963));
AND2X1 g62808(.A (n_11079), .B (n_3915), .Y (n_4815));
NAND3X1 g62834(.A (n_10696), .B (n_2985), .C (n_3985), .Y (n_4813));
INVX1 g64836(.A (g2748), .Y (n_4936));
AOI21X1 g64851(.A0 (n_3863), .A1 (n_4035), .B0 (n_8895), .Y (n_4812));
INVX1 g62839(.A (n_4810), .Y (n_4811));
NAND3X1 g62851(.A (n_4541), .B (g_20159), .C (n_9894), .Y (n_4809));
MX2X1 g62910(.A (n_4805), .B (g_17426), .S0 (n_3177), .Y (n_4806));
AOI21X1 g64979(.A0 (n_326), .A1 (n_3868), .B0 (n_4237), .Y (n_4804));
AOI21X1 g64980(.A0 (n_317), .A1 (n_3868), .B0 (n_4238), .Y (n_4803));
MX2X1 g62941(.A (g5128), .B (n_3983), .S0 (n_9091), .Y (n_4800));
OAI22X1 g62942(.A0 (n_3993), .A1 (n_9772), .B0 (g5134), .B1 (n_9501),.Y (n_4799));
AOI21X1 g61377(.A0 (n_10988), .A1 (g1246), .B0 (n_10989), .Y(n_4798));
MX2X1 g62966(.A (g5485), .B (n_3974), .S0 (n_9172), .Y (n_4797));
DFFSRX1 g5703_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4198), .Q (n_10657), .QN ());
MX2X1 g62990(.A (g5831), .B (n_3973), .S0 (n_8955), .Y (n_4796));
NAND4X1 g61133(.A (n_4765), .B (n_4764), .C (n_4791), .D (n_2529), .Y(n_4795));
MX2X1 g61385(.A (g1246), .B (n_515), .S0 (n_9311), .Y (n_4794));
NAND4X1 g61134(.A (n_4762), .B (n_4761), .C (n_4791), .D (n_2556), .Y(n_4792));
DFFSRX1 g5033_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4200), .Q (g5033), .QN ());
NAND4X1 g61135(.A (n_4758), .B (n_4757), .C (n_4791), .D (n_2280), .Y(n_4790));
MX2X1 g63014(.A (g6177), .B (n_3972), .S0 (n_9000), .Y (n_4789));
NAND4X1 g61136(.A (n_4755), .B (n_4791), .C (n_2244), .D (n_4754), .Y(n_4788));
XOR2X1 g61138(.A (n_952), .B (n_3977), .Y (n_4787));
OAI22X1 g63047(.A0 (n_3992), .A1 (n_9772), .B0 (g6519), .B1 (n_9664),.Y (n_4786));
MX2X1 g63049(.A (g6523), .B (n_3971), .S0 (n_10005), .Y (n_4785));
XOR2X1 g61140(.A (n_967), .B (n_3978), .Y (n_4784));
AOI21X1 g61406(.A0 (n_4220), .A1 (n_1710), .B0 (n_4221), .Y (n_4783));
OAI21X1 g61407(.A0 (n_6953), .A1 (n_7025), .B0 (n_4174), .Y (n_4782));
AOI21X1 g61408(.A0 (n_4218), .A1 (n_1711), .B0 (n_4219), .Y (n_4781));
AOI21X1 g61409(.A0 (n_4216), .A1 (n_2550), .B0 (n_4217), .Y (n_4780));
MX2X1 g61410(.A (g1752), .B (n_6953), .S0 (n_3949), .Y (n_4779));
AOI21X1 g61411(.A0 (n_4214), .A1 (n_1666), .B0 (n_4215), .Y (n_4777));
AOI21X1 g61412(.A0 (n_4211), .A1 (n_1705), .B0 (n_4212), .Y (n_4776));
OAI21X1 g61413(.A0 (n_11039), .A1 (n_10920), .B0 (n_4181), .Y(n_4775));
AOI21X1 g61414(.A0 (n_4209), .A1 (n_1706), .B0 (n_4210), .Y (n_4774));
AOI21X1 g61415(.A0 (n_4207), .A1 (n_2306), .B0 (n_4208), .Y (n_4773));
MX2X1 g61416(.A (g1886), .B (n_11039), .S0 (n_3946), .Y (n_4772));
AOI21X1 g61417(.A0 (n_4203), .A1 (n_1688), .B0 (n_4204), .Y (n_4770));
OAI21X1 g61419(.A0 (n_5057), .A1 (n_7102), .B0 (n_4185), .Y (n_4769));
MX2X1 g61420(.A (g2012), .B (n_5057), .S0 (n_3944), .Y (n_4768));
OAI21X1 g61425(.A0 (n_4743), .A1 (n_10899), .B0 (n_4167), .Y(n_4767));
NAND3X1 g61157(.A (n_4765), .B (n_4764), .C (n_4760), .Y (n_4766));
NAND3X1 g61158(.A (n_4762), .B (n_4761), .C (n_4760), .Y (n_4763));
DFFSRX1 g4438_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4171), .Q (g4438), .QN ());
NAND3X1 g61159(.A (n_4758), .B (n_4757), .C (n_4760), .Y (n_4759));
NAND3X1 g61160(.A (n_4755), .B (n_4760), .C (n_4754), .Y (n_4756));
NOR2X1 g63197(.A (g5073), .B (g5084), .Y (n_4753));
DFFSRX1 g1199_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4257), .Q (g1199), .QN ());
NAND2X1 g63200(.A (n_4159), .B (n_4005), .Y (n_4752));
NAND2X1 g63202(.A (n_4157), .B (n_4002), .Y (n_4751));
NAND2X1 g63204(.A (n_4156), .B (n_4000), .Y (n_4750));
NAND2X1 g63244(.A (n_4154), .B (n_3816), .Y (n_4747));
AOI21X1 g63246(.A0 (n_3411), .A1 (n_10005), .B0 (g5073), .Y (n_4746));
NOR2X1 g61469(.A (n_4743), .B (n_4742), .Y (n_4744));
NOR2X1 g61470(.A (n_4743), .B (n_4740), .Y (n_4741));
NOR2X1 g61472(.A (n_4743), .B (n_4738), .Y (n_4739));
NOR2X1 g61474(.A (n_4743), .B (n_4736), .Y (n_4737));
OAI21X1 g63276(.A0 (n_3776), .A1 (n_9193), .B0 (n_4102), .Y (n_4735));
OAI21X1 g63278(.A0 (n_3780), .A1 (n_9193), .B0 (n_4105), .Y (n_4734));
OAI21X1 g63279(.A0 (n_3777), .A1 (n_9107), .B0 (n_4103), .Y (n_4732));
OAI21X1 g63281(.A0 (n_914), .A1 (n_6685), .B0 (n_4188), .Y (n_4731));
AOI21X1 g63286(.A0 (n_10901), .A1 (g1710), .B0 (n_4173), .Y (n_4730));
AOI22X1 g63303(.A0 (n_903), .A1 (n_10978), .B0 (n_4726), .B1(n_10874), .Y (n_4727));
AOI21X1 g63304(.A0 (n_10874), .A1 (g2671), .B0 (n_4192), .Y (n_4725));
AOI21X1 g63313(.A0 (n_7025), .A1 (g1844), .B0 (n_4189), .Y (n_4723));
AOI21X1 g63315(.A0 (n_10920), .A1 (g1978), .B0 (n_4186), .Y (n_4721));
AOI21X1 g63318(.A0 (n_7102), .A1 (g2112), .B0 (n_4182), .Y (n_4719));
AOI21X1 g63322(.A0 (n_8628), .A1 (g2403), .B0 (n_4178), .Y (n_4717));
AOI21X1 g63324(.A0 (n_8633), .A1 (g2537), .B0 (n_4176), .Y (n_4716));
OAI21X1 g63326(.A0 (n_10899), .A1 (n_6027), .B0 (n_4172), .Y(n_4715));
NAND3X1 g62102(.A (n_2778), .B (n_3904), .C (n_3819), .Y (n_4714));
MX2X1 g63341(.A (n_5961), .B (n_864), .S0 (n_10097), .Y (n_4713));
XOR2X1 g63348(.A (n_6020), .B (n_10873), .Y (n_4712));
XOR2X1 g63349(.A (n_5978), .B (n_3956), .Y (n_4711));
XOR2X1 g63350(.A (n_5975), .B (n_10921), .Y (n_4710));
XOR2X1 g63351(.A (n_6017), .B (n_3953), .Y (n_4709));
XOR2X1 g63352(.A (n_5972), .B (n_3952), .Y (n_4708));
XOR2X1 g63353(.A (n_5969), .B (n_3951), .Y (n_4707));
OAI22X1 g62112(.A0 (n_4050), .A1 (n_4956), .B0 (n_3624), .B1(n_9698), .Y (n_4706));
MX2X1 g63361(.A (g3347), .B (n_3933), .S0 (n_9172), .Y (n_4705));
MX2X1 g63366(.A (g3698), .B (n_3934), .S0 (n_9311), .Y (n_4704));
DFFSRX1 g6049_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4196), .Q (n_11198), .QN ());
DFFSRX1 g3329_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16686), .Q (g3329), .QN ());
DFFSRX1 g3680_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16722), .Q (g3680), .QN ());
DFFSRX1 g1399_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4226), .Q (g19357), .QN ());
NAND3X1 g63482(.A (n_937), .B (n_3929), .C (n_10385), .Y (n_4700));
AOI21X1 g63494(.A0 (n_10372), .A1 (n_4301), .B0 (g2153), .Y (n_4699));
NAND3X1 g63503(.A (n_845), .B (n_3922), .C (n_9351), .Y (n_4695));
NAND2X1 g63507(.A (n_6539), .B (n_10626), .Y (n_4693));
NAND4X1 g61022(.A (n_4638), .B (n_4637), .C (n_4679), .D (n_2535), .Y(n_4690));
AOI22X1 g63548(.A0 (n_615), .A1 (n_3929), .B0 (n_10944), .B1 (g3129),.Y (n_4689));
AOI22X1 g63552(.A0 (n_638), .A1 (n_3922), .B0 (n_4447), .B1 (g3480),.Y (n_4688));
NAND3X1 g60937(.A (n_3911), .B (n_2301), .C (n_4070), .Y (n_4684));
NAND4X1 g63560(.A (n_4682), .B (g3582), .C (g13881), .D (n_10894), .Y(n_4683));
NAND4X1 g61023(.A (n_4633), .B (n_4632), .C (n_4679), .D (n_2538), .Y(n_4680));
NAND4X1 g61024(.A (n_4629), .B (n_4628), .C (n_4679), .D (n_2485), .Y(n_4678));
NAND4X1 g61025(.A (n_4618), .B (n_4679), .C (n_4617), .D (n_3383), .Y(n_4677));
MX2X1 g63629(.A (g1636), .B (g1592), .S0 (n_4108), .Y (n_4676));
MX2X1 g63630(.A (n_4120), .B (g1636), .S0 (n_4108), .Y (n_4673));
NOR3X1 g62253(.A (n_4671), .B (g_19659), .C (n_10078), .Y (n_4672));
MX2X1 g63655(.A (g5236), .B (n_4668), .S0 (n_1205), .Y (n_4670));
MX2X1 g63656(.A (g5252), .B (n_4668), .S0 (n_1225), .Y (n_4669));
MX2X1 g63657(.A (g5264), .B (n_4668), .S0 (n_1465), .Y (n_4667));
MX2X1 g63666(.A (g5583), .B (n_4668), .S0 (n_995), .Y (n_4666));
MX2X1 g63668(.A (g5599), .B (n_4668), .S0 (n_1155), .Y (n_4665));
OAI21X1 g62273(.A0 (n_2584), .A1 (n_3690), .B0 (n_4082), .Y (n_4663));
MX2X1 g63680(.A (g5929), .B (n_4668), .S0 (n_1195), .Y (n_4662));
MX2X1 g63684(.A (g5957), .B (n_4668), .S0 (n_1146), .Y (n_4661));
MX2X1 g63692(.A (g6275), .B (n_4668), .S0 (n_1159), .Y (n_4660));
MX2X1 g63696(.A (g6299), .B (n_4668), .S0 (n_1469), .Y (n_4659));
MX2X1 g63697(.A (g6303), .B (n_4668), .S0 (n_1144), .Y (n_4658));
MX2X1 g63698(.A (g6307), .B (n_4668), .S0 (n_1467), .Y (n_4657));
MX2X1 g63709(.A (g5260), .B (n_4668), .S0 (n_1228), .Y (n_4656));
DFFSRX1 g843_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4250), .Q (g_13278), .QN ());
MX2X1 g63748(.A (g3945), .B (n_4668), .S0 (n_1182), .Y (n_4655));
MX2X1 g63749(.A (g3953), .B (n_4668), .S0 (n_1176), .Y (n_4654));
MX2X1 g63753(.A (g6637), .B (n_4668), .S0 (n_1423), .Y (n_4653));
MX2X1 g63755(.A (g6645), .B (n_4668), .S0 (n_1428), .Y (n_4652));
XOR2X1 g63766(.A (n_2686), .B (n_3929), .Y (n_4651));
XOR2X1 g63767(.A (n_2699), .B (n_3922), .Y (n_4650));
MX2X1 g63782(.A (g2040), .B (g1996), .S0 (n_6758), .Y (n_4649));
MX2X1 g63783(.A (g2070), .B (g2040), .S0 (n_6758), .Y (n_4647));
MX2X1 g63784(.A (g2599), .B (g2555), .S0 (n_10978), .Y (n_4645));
AOI22X1 g62326(.A0 (n_4067), .A1 (n_9359), .B0 (n_659), .B1 (n_9693),.Y (n_4642));
MX2X1 g63785(.A (g2629), .B (g2599), .S0 (n_10978), .Y (n_4640));
NAND3X1 g61039(.A (n_4638), .B (n_4637), .C (n_4631), .Y (n_4639));
MX2X1 g63808(.A (n_10568), .B (n_3905), .S0 (n_9000), .Y (n_4636));
NAND3X1 g61040(.A (n_4633), .B (n_4632), .C (n_4631), .Y (n_4634));
NAND3X1 g61041(.A (n_4629), .B (n_4628), .C (n_4631), .Y (n_4630));
NAND2X1 g61637(.A (n_3755), .B (n_4090), .Y (n_4627));
NAND2X1 g61638(.A (n_3753), .B (n_4092), .Y (n_4626));
DFFSRX1 g4027_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13906), .Q (g16748), .QN ());
NAND3X1 g63869(.A (n_4265), .B (n_4055), .C (n_3903), .Y (n_4625));
NAND3X1 g63870(.A (n_4072), .B (n_4066), .C (n_3736), .Y (n_4624));
NAND3X1 g63871(.A (n_4074), .B (n_4065), .C (n_3735), .Y (n_4623));
NAND3X1 g63872(.A (n_4073), .B (n_4056), .C (n_3734), .Y (n_4622));
NAND3X1 g63873(.A (n_4071), .B (n_4060), .C (n_3733), .Y (n_4621));
NAND3X1 g63874(.A (n_4264), .B (n_4062), .C (n_3902), .Y (n_4620));
NAND3X1 g61043(.A (n_4618), .B (n_4631), .C (n_4617), .Y (n_4619));
INVX1 g63908(.A (n_4615), .Y (n_4616));
NAND3X1 g63932(.A (n_6754), .B (g2084), .C (n_9558), .Y (n_4614));
NAND3X1 g63967(.A (n_10982), .B (n_902), .C (n_9811), .Y (n_4611));
DFFSRX1 g1500_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4233), .Q (g7946), .QN ());
NAND4X1 g64052(.A (g3917), .B (n_5402), .C (g16955), .D (n_6808), .Y(n_4607));
DFFSRX1 g4776_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4227), .Q (g4776), .QN ());
DFFSRX1 g4966_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4201), .Q (g4966), .QN ());
DFFSRX1 g832_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4148), .Q (g_19414), .QN ());
DFFSRX1 g4785_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4136), .Q (g4785), .QN ());
DFFSRX1 g4322_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4081), .Q (n_662), .QN ());
DFFSRX1 g4899_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4083), .Q (g4899), .QN ());
NAND4X1 g64042(.A (g3925), .B (n_3894), .C (g16955), .D (n_8917), .Y(n_4605));
DFFSRX1 g5357_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4199), .Q (n_8807), .QN ());
DFFSRX1 g6741_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4193), .Q (g6741), .QN ());
OAI21X1 g61270(.A0 (n_8761), .A1 (n_8628), .B0 (n_4179), .Y (n_4603));
DFFSRX1 g6395_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4194), .Q (g6395), .QN ());
DFFSRX1 g699_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4137), .Q (g_14265), .QN ());
DFFSRX1 g847_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4135), .Q (g_12791), .QN ());
DFFSRX1 g392_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4110), .Q (g_20268), .QN ());
NAND3X1 g60953(.A (n_4030), .B (n_11220), .C (n_1442), .Y (n_4600));
NAND4X1 g62648(.A (n_4260), .B (n_3442), .C (n_3026), .D (n_3022), .Y(g28030));
DFFSRX1 g4369_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4263), .Q (), .QN (g4369));
NAND3X1 g60955(.A (n_4568), .B (g1373), .C (n_9811), .Y (n_4598));
DFFSRX1 g881_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14096), .Q (g14125), .QN ());
OAI21X1 g61276(.A0 (n_8763), .A1 (n_8633), .B0 (n_4177), .Y (n_4597));
OAI21X1 g61282(.A0 (n_11191), .A1 (n_10874), .B0 (n_4175), .Y(n_4594));
INVX1 g60956(.A (n_4592), .Y (n_4593));
OAI21X1 g60958(.A0 (n_367), .A1 (n_9425), .B0 (n_4246), .Y (n_4591));
NOR2X1 g62576(.A (n_4253), .B (g4704), .Y (n_4590));
NAND3X1 g62598(.A (n_4054), .B (n_2528), .C (n_4028), .Y (n_4589));
NAND2X1 g62609(.A (n_4254), .B (n_3846), .Y (n_4587));
AOI22X1 g60960(.A0 (n_4017), .A1 (n_2586), .B0 (g1542), .B1 (n_9903),.Y (n_4586));
NOR2X1 g62654(.A (n_3243), .B (g4045), .Y (n_4585));
NOR2X1 g61313(.A (n_10761), .B (n_4583), .Y (n_4584));
NOR2X1 g61325(.A (n_940), .B (n_4582), .Y (n_4968));
DFFSRX1 g4975_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4266), .Q (n_11129), .QN ());
NAND2X1 g61795(.A (n_8757), .B (g4608), .Y (n_4581));
DFFSRX1 g2856_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4048), .Q (), .QN (g2856));
OAI21X1 g61834(.A0 (n_4045), .A1 (g_14342), .B0 (n_4578), .Y(n_4579));
NAND3X1 g62807(.A (n_3843), .B (n_2286), .C (n_3824), .Y (n_4577));
INVX1 g62816(.A (n_5723), .Y (n_4576));
DFFSRX1 g2748_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4044), .Q (g2748), .QN ());
OAI21X1 g62840(.A0 (n_4053), .A1 (g_20159), .B0 (n_4202), .Y(n_4810));
NOR2X1 g60978(.A (n_4031), .B (n_4284), .Y (n_4575));
OAI21X1 g62897(.A0 (g2927), .A1 (n_9311), .B0 (n_4029), .Y (n_4574));
OAI21X1 g60980(.A0 (n_10245), .A1 (n_9333), .B0 (n_3995), .Y(n_4573));
NAND4X1 g62918(.A (n_10700), .B (n_3984), .C (n_9359), .D (g5057), .Y(n_4572));
AOI21X1 g62920(.A0 (n_3001), .A1 (n_521), .B0 (n_4022), .Y (n_8879));
OAI22X1 g62927(.A0 (n_3625), .A1 (n_4956), .B0 (n_448), .B1 (n_9862),.Y (n_4570));
INVX1 g60981(.A (n_4568), .Y (n_4569));
MX2X1 g62933(.A (n_3836), .B (g5698), .S0 (n_10660), .Y (n_4567));
MX2X1 g62934(.A (n_3835), .B (g6044), .S0 (n_11201), .Y (n_4566));
MX2X1 g62935(.A (n_3834), .B (g6390), .S0 (g6395), .Y (n_4565));
MX2X1 g62936(.A (n_3833), .B (g6736), .S0 (n_523), .Y (n_4564));
MX2X1 g62939(.A (g5037), .B (n_3825), .S0 (n_9091), .Y (n_4563));
AOI21X1 g61370(.A0 (n_3838), .A1 (n_4558), .B0 (n_3837), .Y (n_4562));
MX2X1 g62943(.A (g5138), .B (n_3809), .S0 (n_8955), .Y (n_4561));
MX2X1 g65047(.A (g6744), .B (g_13901), .S0 (n_9599), .Y (n_4560));
AOI21X1 g61376(.A0 (n_3832), .A1 (n_4558), .B0 (n_3831), .Y (n_4559));
DFFSRX1 g401_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3966), .Q (g_19233), .QN ());
INVX1 g65194(.A (n_7097), .Y (g11678));
MX2X1 g63046(.A (g6513), .B (n_3815), .S0 (n_9359), .Y (n_4557));
AOI21X1 g65434(.A0 (n_4231), .A1 (n_326), .B0 (n_4037), .Y (n_4556));
AOI21X1 g65435(.A0 (n_4231), .A1 (n_317), .B0 (n_4033), .Y (n_4555));
INVX1 g61968(.A (n_8758), .Y (n_4554));
DFFSRX1 g6736_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4011), .Q (g6736), .QN ());
MX2X1 g63142(.A (g_8896), .B (n_3823), .S0 (n_9256), .Y (n_4553));
DFFSRX1 g1389_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3970), .Q (g1389), .QN ());
NAND2X1 g63198(.A (n_3982), .B (n_3830), .Y (n_4550));
DFFSRX1 g1008_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4013), .Q (g_15838), .QN ());
NAND2X1 g63207(.A (n_3813), .B (n_3997), .Y (n_4547));
NAND2X1 g63223(.A (n_9129), .B (g18881), .Y (n_4546));
NOR3X1 g63245(.A (n_9505), .B (g5057), .C (n_10700), .Y (n_4545));
INVX1 g63266(.A (n_4541), .Y (n_4542));
NOR2X1 g61473(.A (n_4743), .B (n_4539), .Y (n_4540));
OAI21X1 g63272(.A0 (n_3792), .A1 (n_9129), .B0 (n_3937), .Y (n_4538));
OAI21X1 g63273(.A0 (n_3788), .A1 (n_9599), .B0 (n_4040), .Y (n_4537));
OAI21X1 g63274(.A0 (n_3786), .A1 (n_9672), .B0 (n_3706), .Y (n_4535));
OAI21X1 g63275(.A0 (n_3785), .A1 (n_9107), .B0 (n_3936), .Y (n_4534));
OAI21X1 g63277(.A0 (n_3781), .A1 (n_9443), .B0 (n_4059), .Y (n_4533));
AOI22X1 g63284(.A0 (n_905), .A1 (n_10857), .B0 (n_4531), .B1(n_8633), .Y (n_4532));
AOI22X1 g63301(.A0 (n_912), .A1 (n_10675), .B0 (n_4529), .B1(n_8628), .Y (n_4530));
MX2X1 g63333(.A (n_4893), .B (n_4527), .S0 (n_10899), .Y (n_4528));
MX2X1 g63334(.A (n_5958), .B (n_716), .S0 (n_10874), .Y (n_4526));
MX2X1 g63337(.A (n_5964), .B (n_856), .S0 (n_10899), .Y (n_4525));
MX2X1 g63338(.A (n_4948), .B (n_854), .S0 (n_7025), .Y (n_4524));
MX2X1 g63339(.A (n_4946), .B (n_871), .S0 (n_10920), .Y (n_4523));
MX2X1 g63340(.A (n_5953), .B (n_862), .S0 (n_7102), .Y (n_4522));
MX2X1 g63342(.A (n_4942), .B (n_846), .S0 (n_8628), .Y (n_4521));
MX2X1 g63344(.A (n_5229), .B (n_714), .S0 (n_8633), .Y (n_4520));
XOR2X1 g62113(.A (g4601), .B (n_8885), .Y (n_4519));
MX2X1 g63367(.A (g4049), .B (n_3770), .S0 (n_9311), .Y (n_4518));
AOI21X1 g63490(.A0 (n_6759), .A1 (n_3943), .B0 (g1996), .Y (n_4516));
NAND2X1 g63495(.A (n_1518), .B (n_10097), .Y (n_4515));
NOR2X1 g63497(.A (n_10099), .B (n_8755), .Y (n_4514));
NAND2X1 g63500(.A (n_10097), .B (n_6025), .Y (n_4513));
AOI21X1 g63523(.A0 (g13895), .A1 (n_464), .B0 (n_3942), .Y (n_4512));
AOI21X1 g63524(.A0 (g13926), .A1 (n_11088), .B0 (n_3941), .Y(n_4510));
OAI21X1 g63541(.A0 (g2878), .A1 (n_9992), .B0 (n_3955), .Y (n_4508));
DFFSRX1 g1536_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3932), .Q (g1536), .QN ());
MX2X1 g63571(.A (n_4497), .B (g5244), .S0 (n_1401), .Y (n_4507));
NOR2X1 g62207(.A (n_3906), .B (n_9836), .Y (n_4506));
MX2X1 g63572(.A (n_4499), .B (g5248), .S0 (n_1404), .Y (n_4504));
MX2X1 g63573(.A (n_4494), .B (g5256), .S0 (n_1463), .Y (n_4503));
MX2X1 g63575(.A (n_4494), .B (g5563), .S0 (n_1761), .Y (n_4502));
MX2X1 g63576(.A (n_4499), .B (g5575), .S0 (n_1322), .Y (n_4501));
MX2X1 g63577(.A (n_4499), .B (g5579), .S0 (n_1413), .Y (n_4500));
MX2X1 g63578(.A (n_4497), .B (g5591), .S0 (n_1397), .Y (n_4498));
MX2X1 g63579(.A (n_4482), .B (g5595), .S0 (n_1408), .Y (n_4496));
MX2X1 g63580(.A (n_4494), .B (g5603), .S0 (n_1477), .Y (n_4495));
MX2X1 g63581(.A (n_4494), .B (g5216), .S0 (n_1738), .Y (n_4493));
MX2X1 g63583(.A (n_4499), .B (g5909), .S0 (n_1728), .Y (n_4492));
MX2X1 g63584(.A (n_4482), .B (g5921), .S0 (n_1108), .Y (n_4490));
MX2X1 g63585(.A (n_4499), .B (g5925), .S0 (n_1114), .Y (n_4489));
MX2X1 g63586(.A (n_4494), .B (g5937), .S0 (n_1120), .Y (n_4488));
MX2X1 g63587(.A (n_4499), .B (g5941), .S0 (n_1104), .Y (n_4487));
MX2X1 g63588(.A (n_4494), .B (g5949), .S0 (n_1452), .Y (n_4486));
MX2X1 g63590(.A (g3119), .B (n_0), .S0 (n_10944), .Y (n_4485));
MX2X1 g63591(.A (n_4482), .B (g6255), .S0 (n_1721), .Y (n_4483));
MX2X1 g63592(.A (n_4494), .B (g6267), .S0 (n_1128), .Y (n_4481));
MX2X1 g63593(.A (n_4499), .B (g6271), .S0 (n_1107), .Y (n_4479));
MX2X1 g63594(.A (n_4497), .B (g6283), .S0 (n_1127), .Y (n_4478));
MX2X1 g63595(.A (n_4482), .B (g6287), .S0 (n_1106), .Y (n_4477));
MX2X1 g63596(.A (n_4494), .B (g3207), .S0 (n_1748), .Y (n_4475));
MX2X1 g63598(.A (n_4482), .B (g3219), .S0 (n_1102), .Y (n_4474));
MX2X1 g63599(.A (n_4499), .B (g3223), .S0 (n_1105), .Y (n_4473));
MX2X1 g63600(.A (n_4482), .B (g3235), .S0 (n_1121), .Y (n_4472));
MX2X1 g63601(.A (n_4482), .B (g3239), .S0 (n_1123), .Y (n_4471));
MX2X1 g63602(.A (n_4494), .B (g6613), .S0 (n_1122), .Y (n_4470));
MX2X1 g63603(.A (n_4497), .B (g3247), .S0 (n_1418), .Y (n_4469));
MX2X1 g63604(.A (n_4497), .B (g6601), .S0 (n_1730), .Y (n_4468));
MX2X1 g63605(.A (n_4494), .B (g6641), .S0 (n_1415), .Y (n_4467));
MX2X1 g63607(.A (n_4497), .B (g3558), .S0 (n_1749), .Y (n_4466));
MX2X1 g63608(.A (n_4499), .B (g3570), .S0 (n_1119), .Y (n_4465));
MX2X1 g63609(.A (n_4494), .B (g3574), .S0 (n_1118), .Y (n_4464));
MX2X1 g63610(.A (n_4494), .B (g3586), .S0 (n_1117), .Y (n_4462));
MX2X1 g63611(.A (n_4482), .B (g3590), .S0 (n_1116), .Y (n_4461));
MX2X1 g63612(.A (n_4494), .B (g3598), .S0 (n_1447), .Y (n_4460));
MX2X1 g63613(.A (n_4482), .B (g5232), .S0 (n_1400), .Y (n_4459));
MX2X1 g63615(.A (n_4482), .B (g5228), .S0 (n_1398), .Y (n_4458));
MX2X1 g63617(.A (n_4499), .B (g3909), .S0 (n_1740), .Y (n_4457));
MX2X1 g63618(.A (n_4497), .B (g3921), .S0 (n_1112), .Y (n_4456));
MX2X1 g63619(.A (n_4494), .B (g3925), .S0 (n_1111), .Y (n_4455));
MX2X1 g63620(.A (n_4494), .B (g3937), .S0 (n_1130), .Y (n_4454));
MX2X1 g63621(.A (n_4482), .B (g3941), .S0 (n_1110), .Y (n_4453));
MX2X1 g63622(.A (n_4482), .B (g3949), .S0 (n_1435), .Y (n_4452));
MX2X1 g63626(.A (n_4497), .B (g6633), .S0 (n_1392), .Y (n_4451));
MX2X1 g63627(.A (n_4494), .B (g6295), .S0 (n_1433), .Y (n_4450));
MX2X1 g63628(.A (n_4482), .B (g6629), .S0 (n_1393), .Y (n_4449));
MX2X1 g63631(.A (g3470), .B (n_60), .S0 (n_4447), .Y (n_4448));
MX2X1 g63632(.A (n_4482), .B (g6617), .S0 (n_1103), .Y (n_4446));
AOI22X1 g63637(.A0 (n_3609), .A1 (n_9443), .B0 (n_10944), .B1(n_901), .Y (n_4445));
AOI22X1 g63639(.A0 (n_3601), .A1 (n_10078), .B0 (n_4447), .B1(n_2019), .Y (n_4444));
MX2X1 g63649(.A (n_4497), .B (g5196), .S0 (n_1775), .Y (n_4442));
MX2X1 g63650(.A (n_4499), .B (g5200), .S0 (n_1764), .Y (n_4441));
MX2X1 g63651(.A (n_4482), .B (g5204), .S0 (n_1481), .Y (n_4440));
MX2X1 g63652(.A (n_4499), .B (g5208), .S0 (n_1605), .Y (n_4439));
MX2X1 g63653(.A (n_4499), .B (g5220), .S0 (n_1178), .Y (n_4438));
MX2X1 g63654(.A (n_4482), .B (g5224), .S0 (n_1438), .Y (n_4437));
MX2X1 g63658(.A (n_4497), .B (g6235), .S0 (n_1779), .Y (n_4436));
MX2X1 g63659(.A (g5272), .B (n_4497), .S0 (g26801), .Y (n_4434));
MX2X1 g63660(.A (n_4497), .B (g5543), .S0 (n_1773), .Y (n_4433));
MX2X1 g63661(.A (n_4497), .B (g5547), .S0 (n_1778), .Y (n_4432));
MX2X1 g63662(.A (n_4499), .B (g5551), .S0 (n_1425), .Y (n_4431));
MX2X1 g63663(.A (n_4499), .B (g5559), .S0 (n_1131), .Y (n_4430));
MX2X1 g63664(.A (n_4499), .B (g5567), .S0 (n_1235), .Y (n_4429));
MX2X1 g63665(.A (n_4482), .B (g5571), .S0 (n_1466), .Y (n_4428));
MX2X1 g63667(.A (n_4482), .B (g5587), .S0 (n_1424), .Y (n_4427));
MX2X1 g63669(.A (g5607), .B (n_4424), .S0 (n_1187), .Y (n_4426));
MX2X1 g63670(.A (g5611), .B (n_4424), .S0 (n_1223), .Y (n_4425));
MX2X1 g63671(.A (g5615), .B (n_4424), .S0 (n_1239), .Y (n_4423));
OAI21X1 g62272(.A0 (n_3885), .A1 (n_1285), .B0 (n_3184), .Y (n_4422));
MX2X1 g63672(.A (n_4482), .B (g5619), .S0 (n_4329), .Y (n_4421));
MX2X1 g63673(.A (n_4497), .B (g5889), .S0 (n_1722), .Y (n_4420));
MX2X1 g63674(.A (n_4482), .B (g5893), .S0 (n_1726), .Y (n_4419));
MX2X1 g63675(.A (n_4482), .B (g5897), .S0 (n_1437), .Y (n_4418));
MX2X1 g63676(.A (n_4494), .B (g5901), .S0 (n_1755), .Y (n_4417));
MX2X1 g63677(.A (n_4499), .B (g5905), .S0 (n_1170), .Y (n_4416));
MX2X1 g63678(.A (n_4499), .B (g5913), .S0 (n_999), .Y (n_4415));
MX2X1 g63679(.A (n_4499), .B (g5917), .S0 (n_1456), .Y (n_4414));
MX2X1 g63681(.A (n_4499), .B (g5933), .S0 (n_1431), .Y (n_4413));
MX2X1 g63682(.A (g6621), .B (n_4424), .S0 (n_1152), .Y (n_4412));
MX2X1 g63683(.A (g5945), .B (n_4497), .S0 (n_1247), .Y (n_4411));
MX2X1 g63685(.A (g5961), .B (n_4497), .S0 (n_910), .Y (n_4410));
MX2X1 g63686(.A (n_4482), .B (g5965), .S0 (n_4327), .Y (n_4409));
MX2X1 g63687(.A (n_4494), .B (g6243), .S0 (n_1419), .Y (n_4408));
MX2X1 g63688(.A (n_4482), .B (g6247), .S0 (n_1771), .Y (n_4407));
MX2X1 g63689(.A (n_4482), .B (g6251), .S0 (n_1215), .Y (n_4406));
MX2X1 g63690(.A (n_4497), .B (g6259), .S0 (n_1153), .Y (n_4405));
MX2X1 g63691(.A (n_4482), .B (g6263), .S0 (n_1472), .Y (n_4404));
MX2X1 g63693(.A (g5953), .B (n_4424), .S0 (n_1460), .Y (n_4403));
MX2X1 g63694(.A (n_4494), .B (g6279), .S0 (n_1470), .Y (n_4402));
MX2X1 g63695(.A (g6291), .B (n_4424), .S0 (n_1150), .Y (n_4401));
MX2X1 g63699(.A (g5268), .B (n_4424), .S0 (n_1232), .Y (n_4400));
MX2X1 g63700(.A (n_4494), .B (g6311), .S0 (n_4324), .Y (n_4399));
MX2X1 g63701(.A (n_4497), .B (g3187), .S0 (n_1769), .Y (n_4398));
MX2X1 g63702(.A (n_4499), .B (g3191), .S0 (n_1759), .Y (n_4397));
MX2X1 g63703(.A (n_4499), .B (g3195), .S0 (n_1427), .Y (n_4396));
MX2X1 g63704(.A (n_4494), .B (g3199), .S0 (n_1768), .Y (n_4395));
MX2X1 g63705(.A (n_4497), .B (g3211), .S0 (n_1136), .Y (n_4394));
MX2X1 g63707(.A (n_4499), .B (g3203), .S0 (n_993), .Y (n_4393));
MX2X1 g63706(.A (n_4482), .B (g3215), .S0 (n_1585), .Y (n_4392));
MX2X1 g63708(.A (g3227), .B (n_4424), .S0 (n_1244), .Y (n_4391));
MX2X1 g63710(.A (n_4499), .B (g3231), .S0 (n_1478), .Y (n_4390));
MX2X1 g63711(.A (n_4499), .B (g6593), .S0 (n_1780), .Y (n_4389));
MX2X1 g63712(.A (n_4497), .B (g6581), .S0 (n_1766), .Y (n_4388));
MX2X1 g63713(.A (g3243), .B (n_4497), .S0 (n_1148), .Y (n_4387));
MX2X1 g63714(.A (g3255), .B (n_4497), .S0 (n_1483), .Y (n_4386));
MX2X1 g63715(.A (g3259), .B (n_4497), .S0 (n_897), .Y (n_4385));
MX2X1 g63716(.A (g6649), .B (n_4424), .S0 (n_1487), .Y (n_4384));
MX2X1 g63717(.A (g6653), .B (n_4424), .S0 (n_1326), .Y (n_4383));
MX2X1 g63718(.A (n_4494), .B (g6657), .S0 (n_4322), .Y (n_4382));
MX2X1 g63719(.A (n_4497), .B (g5240), .S0 (n_1453), .Y (n_4381));
MX2X1 g63720(.A (g3251), .B (n_4497), .S0 (n_1475), .Y (n_4380));
MX2X1 g63721(.A (n_4494), .B (g3538), .S0 (n_1754), .Y (n_4379));
MX2X1 g63722(.A (n_4499), .B (g3542), .S0 (n_1753), .Y (n_4378));
MX2X1 g63723(.A (n_4499), .B (g3546), .S0 (n_1451), .Y (n_4377));
MX2X1 g63724(.A (n_4494), .B (g3550), .S0 (n_1750), .Y (n_4376));
MX2X1 g63725(.A (n_4497), .B (g3554), .S0 (n_1211), .Y (n_4375));
MX2X1 g63726(.A (n_4494), .B (g3562), .S0 (n_1209), .Y (n_4374));
MX2X1 g63727(.A (n_4494), .B (g3566), .S0 (n_1449), .Y (n_4373));
MX2X1 g63728(.A (g3578), .B (n_4424), .S0 (n_1208), .Y (n_4372));
MX2X1 g63729(.A (n_4494), .B (g3582), .S0 (n_1448), .Y (n_4371));
MX2X1 g63730(.A (g3594), .B (n_4424), .S0 (n_1202), .Y (n_4370));
MX2X1 g63731(.A (n_4482), .B (g6609), .S0 (n_1432), .Y (n_4369));
MX2X1 g63732(.A (g3602), .B (n_4424), .S0 (n_1200), .Y (n_4368));
MX2X1 g63733(.A (g3606), .B (n_4424), .S0 (n_1198), .Y (n_4367));
MX2X1 g63734(.A (n_4499), .B (g6589), .S0 (n_1446), .Y (n_4366));
MX2X1 g63735(.A (g3610), .B (n_4424), .S0 (n_931), .Y (n_4365));
MX2X1 g63736(.A (n_4497), .B (g3614), .S0 (n_4320), .Y (n_4364));
MX2X1 g63737(.A (n_4499), .B (g6597), .S0 (n_1217), .Y (n_4363));
MX2X1 g63738(.A (n_4497), .B (g3889), .S0 (n_1746), .Y (n_4362));
MX2X1 g63739(.A (n_4482), .B (g3893), .S0 (n_1745), .Y (n_4361));
MX2X1 g63740(.A (n_4497), .B (g6239), .S0 (n_1724), .Y (n_4360));
MX2X1 g63741(.A (n_4494), .B (g3897), .S0 (n_1441), .Y (n_4359));
MX2X1 g63742(.A (n_4499), .B (g3901), .S0 (n_1741), .Y (n_4358));
MX2X1 g63743(.A (n_4482), .B (g3905), .S0 (n_1192), .Y (n_4357));
MX2X1 g63744(.A (n_4482), .B (g3913), .S0 (n_1189), .Y (n_4356));
MX2X1 g63745(.A (n_4494), .B (g3917), .S0 (n_1439), .Y (n_4355));
MX2X1 g63746(.A (g3929), .B (n_4424), .S0 (n_1186), .Y (n_4354));
MX2X1 g63747(.A (n_4482), .B (g3933), .S0 (n_1436), .Y (n_4353));
MX2X1 g63750(.A (g3957), .B (n_4497), .S0 (n_1174), .Y (n_4352));
MX2X1 g63751(.A (g3961), .B (n_4497), .S0 (n_921), .Y (n_4351));
MX2X1 g63752(.A (n_4499), .B (g3965), .S0 (n_4314), .Y (n_4350));
MX2X1 g63754(.A (n_4499), .B (g6605), .S0 (n_1167), .Y (n_4349));
MX2X1 g63756(.A (n_4494), .B (g3263), .S0 (n_4316), .Y (n_4348));
MX2X1 g63758(.A (n_4482), .B (g5212), .S0 (n_1164), .Y (n_4347));
MX2X1 g63759(.A (n_4494), .B (g6585), .S0 (n_1719), .Y (n_4346));
MX2X1 g63760(.A (n_4497), .B (g5555), .S0 (n_1716), .Y (n_4345));
MX2X1 g63761(.A (n_4494), .B (g6625), .S0 (n_1416), .Y (n_4344));
MX2X1 g63773(.A (g2465), .B (g2421), .S0 (n_10853), .Y (n_4343));
MX2X1 g63774(.A (n_4339), .B (g2465), .S0 (n_10853), .Y (n_4340));
MX2X1 g63778(.A (g_12791), .B (n_3745), .S0 (n_9992), .Y (n_4338));
MX2X1 g63779(.A (g2331), .B (g2287), .S0 (n_10671), .Y (n_4336));
MX2X1 g63780(.A (g2361), .B (g2331), .S0 (n_10671), .Y (n_4333));
NAND3X1 g63868(.A (n_4076), .B (n_3883), .C (n_3737), .Y (n_4331));
AND2X1 g63909(.A (n_4424), .B (n_1812), .Y (n_4615));
AND2X1 g63914(.A (n_4329), .B (n_4668), .Y (n_4330));
AND2X1 g63917(.A (n_4327), .B (n_4668), .Y (n_4328));
AND2X1 g63922(.A (n_4324), .B (n_4668), .Y (n_4325));
AND2X1 g63923(.A (n_4668), .B (n_4322), .Y (n_4323));
AND2X1 g63929(.A (n_4320), .B (n_4668), .Y (n_4321));
NOR2X1 g63930(.A (n_4304), .B (n_4318), .Y (n_4319));
AND2X1 g63931(.A (n_4316), .B (n_4668), .Y (n_4317));
AND2X1 g63933(.A (n_4314), .B (n_4668), .Y (n_4315));
INVX1 g63940(.A (n_10626), .Y (n_4313));
NAND3X1 g63952(.A (n_10670), .B (n_911), .C (n_9091), .Y (n_10549));
NAND3X1 g63958(.A (n_10852), .B (n_904), .C (n_10005), .Y (n_4308));
NOR2X1 g63971(.A (n_670), .B (n_4304), .Y (n_4306));
NOR2X1 g63973(.A (n_290), .B (n_4304), .Y (n_4305));
NOR2X1 g63974(.A (n_667), .B (n_4304), .Y (n_4303));
NAND4X1 g64001(.A (n_3907), .B (n_3371), .C (n_10063), .D (n_3486),.Y (n_4302));
NAND3X1 g64002(.A (n_4299), .B (n_4301), .C (g2153), .Y (n_4836));
NAND3X1 g64004(.A (n_10372), .B (g2197), .C (n_259), .Y (n_4834));
NAND3X1 g64005(.A (n_4299), .B (g2227), .C (g2153), .Y (n_4829));
DFFSRX1 g817_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4010), .Q (g_16792), .QN ());
NAND3X1 g64007(.A (n_4299), .B (n_4301), .C (g2227), .Y (n_4827));
DFFSRX1 g1576_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3969), .Q (g10527), .QN ());
NAND3X1 g60952(.A (n_3702), .B (n_2779), .C (n_3848), .Y (n_4298));
DFFSRX1 g4709_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3979), .Q (g4709), .QN ());
DFFSRX1 g969_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4069), .Q (g_13091), .QN ());
DFFSRX1 g5698_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4015), .Q (g5698), .QN ());
DFFSRX1 g6044_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4014), .Q (g6044), .QN ());
DFFSRX1 g6390_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4012), .Q (g6390), .QN ());
DFFSRX1 g5352_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4016), .Q (g5352), .QN ());
DFFSRX1 g1056_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4008), .Q (g19334), .QN ());
DFFSRX1 g4176_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4009), .Q (g4176), .QN ());
DFFSRX1 g4191_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3991), .Q (g11447), .QN ());
DFFSRX1 g528_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3981), .Q (g_8896), .QN ());
DFFSRX1 g837_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3968), .Q (g_15740), .QN ());
DFFSRX1 g405_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3964), .Q (n_11163), .QN ());
DFFSRX1 g424_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3963), .Q (g_21778), .QN ());
DFFSRX1 g429_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3962), .Q (g_17065), .QN ());
DFFSRX1 g433_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3960), .Q (g_16677), .QN ());
DFFSRX1 g437_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3959), .Q (g_21720), .QN ());
DFFSRX1 g441_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3958), .Q (g_13758), .QN ());
DFFSRX1 g475_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3957), .Q (g_19289), .QN ());
DFFSRX1 g417_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3947), .Q (n_640), .QN ());
DFFSRX1 g2719_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_4034), .Q (n_8898), .QN ());
NAND3X1 g64135(.A (n_4046), .B (n_2589), .C (n_3882), .Y (n_4297));
INVX1 g64188(.A (n_6754), .Y (n_4296));
OAI21X1 g60957(.A0 (n_3910), .A1 (g1373), .B0 (n_10427), .Y (n_4592));
INVX1 g64222(.A (n_4885), .Y (n_4293));
NAND3X1 g64279(.A (n_3878), .B (n_637), .C (n_3879), .Y (n_4291));
AOI21X1 g62583(.A0 (n_3856), .A1 (n_2310), .B0 (n_9772), .Y (n_4290));
MX2X1 g64407(.A (n_11106), .B (g14217), .S0 (n_5582), .Y (n_4288));
OAI22X1 g62656(.A0 (n_3492), .A1 (n_3192), .B0 (g4366), .B1 (n_9874),.Y (n_4286));
AOI22X1 g60961(.A0 (n_4284), .A1 (n_10196), .B0 (n_1179), .B1(g7946), .Y (n_4285));
NAND2X1 g61316(.A (n_2619), .B (n_4170), .Y (n_4283));
NOR2X1 g61317(.A (n_8761), .B (n_4281), .Y (n_4282));
NOR2X1 g61318(.A (n_8762), .B (n_4279), .Y (n_4280));
NOR2X1 g61319(.A (n_8762), .B (n_4277), .Y (n_4278));
NOR2X1 g61320(.A (n_8762), .B (n_4275), .Y (n_4276));
NOR2X1 g61321(.A (n_8763), .B (n_4273), .Y (n_4274));
NOR2X1 g61322(.A (n_8764), .B (n_4271), .Y (n_4272));
NOR2X1 g61323(.A (n_8764), .B (n_4269), .Y (n_4270));
NOR2X1 g61324(.A (n_8764), .B (n_4267), .Y (n_4268));
XOR2X1 g61083(.A (g1300), .B (n_11025), .Y (n_4618));
MX2X1 g62727(.A (n_684), .B (n_3677), .S0 (n_9218), .Y (n_4266));
DFFSRX1 g4045_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3847), .Q (), .QN (g4045));
NAND4X1 g64714(.A (g5802), .B (n_9627), .C (g9617), .D (g_7062), .Y(n_4265));
NAND4X1 g64728(.A (g3451), .B (n_9521), .C (g8279), .D (g_5313), .Y(n_4264));
MX2X1 g64778(.A (g4459), .B (g4473), .S0 (n_9091), .Y (n_4263));
AND2X1 g62805(.A (n_327), .B (g4366), .Y (n_4262));
CLKBUFX1 g62817(.A (n_7145), .Y (n_5723));
AOI21X1 g62836(.A0 (n_3287), .A1 (n_2747), .B0 (n_3852), .Y (n_4260));
OAI21X1 g62898(.A0 (n_10644), .A1 (n_9681), .B0 (n_3851), .Y(n_4257));
OR2X1 g64931(.A (g5109), .B (n_9398), .Y (n_4255));
AOI22X1 g62903(.A0 (n_3659), .A1 (n_2585), .B0 (g1199), .B1 (n_9628),.Y (n_4254));
OAI22X1 g62911(.A0 (n_10830), .A1 (g5348), .B0 (n_1058), .B1 (g5352),.Y (n_4253));
NAND4X1 g62913(.A (n_3661), .B (n_4024), .C (n_9811), .D (g_18793),.Y (n_4252));
AOI22X1 g62916(.A0 (n_10621), .A1 (g5348), .B0 (g5352), .B1 (g25114),.Y (n_4251));
OAI21X1 g62923(.A0 (n_708), .A1 (n_9311), .B0 (n_3858), .Y (n_4250));
INVX1 g60982(.A (n_10427), .Y (n_4568));
INVX1 g65050(.A (n_4247), .Y (n_4248));
NAND4X1 g60985(.A (n_4242), .B (n_9209), .C (n_4241), .D (n_2593), .Y(n_4246));
AOI21X1 g61381(.A0 (n_10323), .A1 (g1246), .B0 (n_10321), .Y(n_4582));
NAND4X1 g60987(.A (n_4242), .B (n_4241), .C (n_9558), .D (n_16), .Y(n_4243));
NOR2X1 g65269(.A (g2819), .B (n_3868), .Y (n_4239));
NOR2X1 g65272(.A (g2807), .B (n_3868), .Y (n_4238));
NOR2X1 g65273(.A (g2775), .B (n_3868), .Y (n_4237));
NAND2X1 g65298(.A (g_13901), .B (n_9717), .Y (n_5573));
NOR2X1 g65350(.A (g2787), .B (n_3868), .Y (n_4235));
OAI22X1 g60989(.A0 (n_3692), .A1 (n_9193), .B0 (n_2474), .B1(n_9992), .Y (n_4233));
DFFSRX1 g5016_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3808), .Q (g5016), .QN ());
MX2X1 g65433(.A (g2787), .B (g2783), .S0 (n_4231), .Y (n_4232));
MX2X1 g65436(.A (g2819), .B (g2815), .S0 (n_4231), .Y (n_4230));
AOI21X1 g60990(.A0 (n_2773), .A1 (n_3849), .B0 (n_3861), .Y(n_11220));
NAND3X1 g61959(.A (n_2520), .B (n_3652), .C (n_3717), .Y (n_4227));
MX2X1 g60991(.A (g1333), .B (n_3629), .S0 (n_9091), .Y (n_4226));
MX2X1 g65491(.A (g2079), .B (g1945), .S0 (n_4231), .Y (n_4225));
MX2X1 g65492(.A (g2638), .B (g2504), .S0 (n_4231), .Y (n_4224));
NAND2X1 g65934(.A (g2370), .B (n_3679), .Y (n_4223));
AND2X1 g63194(.A (n_3828), .B (n_1285), .Y (n_11079));
NOR2X1 g61451(.A (n_6953), .B (n_4220), .Y (n_4221));
NOR2X1 g61452(.A (n_6954), .B (n_4218), .Y (n_4219));
NOR2X1 g61455(.A (n_6954), .B (n_4216), .Y (n_4217));
NOR2X1 g61456(.A (n_6954), .B (n_4214), .Y (n_4215));
NAND2X1 g63224(.A (n_3821), .B (n_1576), .Y (n_4213));
NOR2X1 g61458(.A (n_11039), .B (n_4211), .Y (n_4212));
NOR2X1 g61459(.A (n_11040), .B (n_4209), .Y (n_4210));
NOR2X1 g61460(.A (n_11040), .B (n_4207), .Y (n_4208));
NOR2X1 g63235(.A (n_3817), .B (n_2163), .Y (n_4206));
NAND3X1 g63236(.A (n_3826), .B (n_2988), .C (n_2423), .Y (n_4205));
NOR2X1 g61461(.A (n_11040), .B (n_4203), .Y (n_4204));
DFFSRX1 g1157_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3795), .Q (g7916), .QN ());
INVX1 g63267(.A (n_4202), .Y (n_4541));
NAND3X1 g62104(.A (n_2798), .B (n_3564), .C (n_3683), .Y (n_4201));
DFFSRX1 g2917_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3766), .Q (), .QN (g2917));
MX2X1 g63347(.A (g5029), .B (n_3637), .S0 (n_9797), .Y (n_4200));
MX2X1 g63354(.A (g5352), .B (n_3631), .S0 (n_8955), .Y (n_4199));
MX2X1 g63355(.A (g5698), .B (n_3633), .S0 (n_9240), .Y (n_4198));
MX2X1 g63356(.A (g6044), .B (n_3634), .S0 (n_9234), .Y (n_4196));
MX2X1 g63357(.A (g6390), .B (n_3627), .S0 (n_9834), .Y (n_4194));
MX2X1 g63362(.A (g6736), .B (n_3549), .S0 (n_9750), .Y (n_4193));
DFFSRX1 g5073_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3771), .Q (), .QN (g5073));
NOR2X1 g63430(.A (n_717), .B (n_10874), .Y (n_4192));
NOR2X1 g63442(.A (n_855), .B (n_7025), .Y (n_4189));
NAND2X1 g63443(.A (n_4187), .B (n_10920), .Y (n_4188));
NOR2X1 g63444(.A (n_872), .B (n_10920), .Y (n_4186));
NAND2X1 g63445(.A (n_1514), .B (n_7102), .Y (n_4185));
NAND2X1 g63446(.A (n_4183), .B (n_7102), .Y (n_4184));
NOR2X1 g63447(.A (n_863), .B (n_7102), .Y (n_4182));
NAND2X1 g63448(.A (n_1687), .B (n_10920), .Y (n_4181));
AOI21X1 g61018(.A0 (n_3459), .A1 (n_2177), .B0 (n_3811), .Y (n_4180));
NAND2X1 g63449(.A (n_1676), .B (n_8628), .Y (n_4179));
NOR2X1 g63450(.A (n_847), .B (n_8628), .Y (n_4178));
NAND2X1 g63452(.A (n_1670), .B (n_8633), .Y (n_4177));
NOR2X1 g63456(.A (n_715), .B (n_8633), .Y (n_4176));
NAND2X1 g63458(.A (n_1505), .B (n_10874), .Y (n_4175));
NAND2X1 g63459(.A (n_1665), .B (n_7025), .Y (n_4174));
NOR2X1 g63463(.A (n_857), .B (n_10901), .Y (n_4173));
NAND2X1 g63465(.A (n_10901), .B (n_6027), .Y (n_4172));
INVX1 g63498(.A (n_4170), .Y (n_4171));
AOI21X1 g63502(.A0 (n_10672), .A1 (n_4038), .B0 (g2287), .Y (n_4169));
AOI21X1 g63506(.A0 (n_10854), .A1 (n_3939), .B0 (g2421), .Y (n_4168));
NAND2X1 g63510(.A (n_1509), .B (n_10901), .Y (n_4167));
AOI22X1 g63546(.A0 (n_639), .A1 (n_10473), .B0 (n_10472), .B1(g5831), .Y (n_4165));
DFFSRX1 g2882_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3877), .Q (), .QN (g2882));
MX2X1 g63574(.A (g5475), .B (n_94), .S0 (n_10342), .Y (n_4163));
MX2X1 g63582(.A (g5821), .B (n_65), .S0 (n_10472), .Y (n_4161));
MX2X1 g63589(.A (g6167), .B (n_125), .S0 (n_10444), .Y (n_4160));
AOI21X1 g63634(.A0 (n_3616), .A1 (n_9903), .B0 (n_3803), .Y (n_4159));
AOI21X1 g63635(.A0 (n_3611), .A1 (n_9903), .B0 (n_3802), .Y (n_4157));
AOI21X1 g63636(.A0 (n_3589), .A1 (n_9019), .B0 (n_3801), .Y (n_4156));
OAI21X1 g62260(.A0 (n_3447), .A1 (g_15381), .B0 (n_3448), .Y(n_4155));
AOI21X1 g63647(.A0 (g5041), .A1 (n_9856), .B0 (n_3800), .Y (n_4154));
OAI21X1 g62274(.A0 (n_3715), .A1 (n_3569), .B0 (n_3242), .Y (n_4152));
AOI21X1 g61213(.A0 (n_10289), .A1 (n_4149), .B0 (n_10285), .Y(n_4151));
AOI21X1 g61214(.A0 (n_6951), .A1 (n_4149), .B0 (n_3873), .Y (n_4150));
OAI22X1 g62293(.A0 (n_4939), .A1 (n_3686), .B0 (n_10496), .B1(n_9466), .Y (n_4148));
MX2X1 g63770(.A (g1906), .B (g1862), .S0 (n_6677), .Y (n_4147));
MX2X1 g63771(.A (g1936), .B (g1906), .S0 (n_6677), .Y (n_4145));
MX2X1 g63775(.A (g1772), .B (g1728), .S0 (n_10916), .Y (n_4142));
MX2X1 g63776(.A (n_4139), .B (g1772), .S0 (n_10913), .Y (n_4140));
MX2X1 g63777(.A (g_17934), .B (n_3572), .S0 (n_10005), .Y (n_4137));
MX2X1 g62324(.A (n_10818), .B (n_3708), .S0 (n_9240), .Y (n_4136));
OAI22X1 g63781(.A0 (n_3570), .A1 (n_9976), .B0 (g_22639), .B1(n_9830), .Y (n_4135));
XOR2X1 g61225(.A (g_11413), .B (n_4134), .Y (n_4765));
XOR2X1 g61226(.A (g_16456), .B (n_4134), .Y (n_4762));
XOR2X1 g61227(.A (g_20563), .B (n_4134), .Y (n_4758));
XOR2X1 g61228(.A (g_18869), .B (n_4134), .Y (n_4755));
DFFSRX1 g3676_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13881), .Q (g16722), .QN ());
DFFSRX1 g3325_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13865), .Q (g16686), .QN ());
NAND3X1 g63919(.A (n_10912), .B (g1816), .C (n_9698), .Y (n_4133));
NAND3X1 g63928(.A (n_6685), .B (g1950), .C (n_9448), .Y (n_4131));
OR2X1 g63946(.A (n_11094), .B (g_15691), .Y (n_4126));
NOR2X1 g63948(.A (n_4124), .B (n_10674), .Y (n_4125));
NOR2X1 g63954(.A (n_4122), .B (n_10856), .Y (n_4123));
NAND2X1 g63955(.A (n_4108), .B (n_4120), .Y (n_4121));
NOR2X1 g63965(.A (n_6666), .B (n_4118), .Y (n_4119));
NOR2X1 g63975(.A (n_618), .B (n_6666), .Y (n_4117));
NOR2X1 g63977(.A (n_342), .B (n_6666), .Y (n_4113));
NOR2X1 g63978(.A (n_624), .B (n_6666), .Y (n_4111));
NAND3X1 g63999(.A (n_3567), .B (n_2256), .C (n_3551), .Y (n_4110));
OR2X1 g64006(.A (n_10380), .B (n_4109), .Y (n_4583));
DFFSRX1 g4311_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3798), .Q (g4311), .QN ());
NAND3X1 g64018(.A (n_4108), .B (g1592), .C (n_347), .Y (n_4742));
NAND3X1 g64019(.A (n_4108), .B (g1636), .C (n_629), .Y (n_4740));
NAND3X1 g64020(.A (n_4108), .B (g1592), .C (n_4120), .Y (n_4738));
NAND2X1 g64023(.A (n_4108), .B (g25259), .Y (n_4736));
DFFSRX1 g1211_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3840), .Q (n_8800), .QN ());
DFFSRX1 g4801_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3810), .Q (n_8915), .QN ());
DFFSRX1 g4991_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3738), .Q (g4991), .QN ());
NAND4X1 g64038(.A (g3574), .B (n_10893), .C (g16924), .D (n_6973), .Y(n_4107));
AOI21X1 g64041(.A0 (n_6978), .A1 (n_9019), .B0 (n_3744), .Y (n_4105));
AOI21X1 g64044(.A0 (g4054), .A1 (n_9772), .B0 (n_3742), .Y (n_4103));
AOI21X1 g64045(.A0 (n_7003), .A1 (n_9836), .B0 (n_3746), .Y (n_4102));
NAND4X1 g64049(.A (g3566), .B (n_10895), .C (g16924), .D (n_11128),.Y (n_4101));
DFFSRX1 g1193_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3886), .Q (n_10649), .QN ());
DFFSRX1 g2898_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3839), .Q (), .QN (g2898));
DFFSRX1 g79_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3859), .Q (g20899), .QN ());
DFFSRX1 g2999_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3807), .Q (g2999), .QN ());
DFFSRX1 g4287_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3767), .Q (g9019), .QN ());
DFFSRX1 g5037_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3793), .Q (g5037), .QN ());
DFFSRX1 g2729_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3869), .Q (n_10656), .QN ());
DFFSRX1 g4023_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16955), .Q (g13906), .QN ());
OR2X1 g64141(.A (g3808), .B (n_4096), .Y (n_6049));
NAND4X1 g64216(.A (g3901), .B (n_6787), .C (g14518), .D (n_3894), .Y(n_4098));
NAND2X1 g64223(.A (n_11208), .B (n_4096), .Y (n_4885));
INVX1 g62564(.A (n_6551), .Y (n_4671));
NAND3X1 g61737(.A (n_3891), .B (n_10184), .C (n_4091), .Y (n_4092));
NAND3X1 g61738(.A (n_3893), .B (n_10205), .C (n_4091), .Y (n_4090));
NAND4X1 g64378(.A (n_4988), .B (g3889), .C (g14518), .D (n_5402), .Y(n_4088));
AOI21X1 g64398(.A0 (n_3897), .A1 (n_245), .B0 (n_3898), .Y (n_4087));
AOI21X1 g64399(.A0 (n_3730), .A1 (n_282), .B0 (n_3731), .Y (n_4086));
AOI21X1 g64400(.A0 (n_3728), .A1 (n_360), .B0 (n_3729), .Y (n_4085));
AOI21X1 g64401(.A0 (n_3726), .A1 (n_3135), .B0 (n_3727), .Y (n_4084));
OAI21X1 g62662(.A0 (n_3514), .A1 (n_9371), .B0 (n_3881), .Y (n_4083));
AOI22X1 g62666(.A0 (n_3691), .A1 (n_3857), .B0 (g_13278), .B1(n_9129), .Y (n_4082));
OAI22X1 g62677(.A0 (n_3648), .A1 (n_3797), .B0 (n_327), .B1(n_10005), .Y (n_4081));
DFFSRX1 g878_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14217), .Q (g14096), .QN ());
NAND4X1 g64524(.A (g5109), .B (n_9627), .C (g9497), .D (n_107), .Y(n_4080));
XOR2X1 g61080(.A (g1478), .B (n_11025), .Y (n_4638));
XOR2X1 g61081(.A (g1448), .B (n_11026), .Y (n_4633));
XOR2X1 g61082(.A (g1472), .B (n_11026), .Y (n_4629));
NAND4X1 g64711(.A (g5456), .B (n_9627), .C (g9555), .D (g_5508), .Y(n_4076));
NAND4X1 g64720(.A (g6148), .B (n_9627), .C (g9682), .D (g_14965), .Y(n_4074));
NAND4X1 g64722(.A (g6494), .B (n_9627), .C (g9743), .D (g_3861), .Y(n_4073));
NAND4X1 g64726(.A (g3100), .B (n_9627), .C (g8215), .D (g_6579), .Y(n_4072));
NAND4X1 g64729(.A (g3802), .B (n_9627), .C (g8344), .D (g_5156), .Y(n_4071));
NAND3X1 g60973(.A (n_10429), .B (g1367), .C (n_9717), .Y (n_4070));
NOR2X1 g62791(.A (n_3685), .B (n_9775), .Y (n_4069));
AOI21X1 g62799(.A0 (n_1349), .A1 (n_2471), .B0 (n_3680), .Y (n_4068));
DFFSRX1 g1061_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3703), .Q (n_8509), .QN ());
NAND2X1 g62826(.A (n_3681), .B (n_3822), .Y (n_4067));
NOR2X1 g64854(.A (n_3697), .B (n_8557), .Y (n_5703));
OR2X1 g64861(.A (g3100), .B (n_9398), .Y (n_4066));
OR2X1 g64866(.A (g6148), .B (n_9398), .Y (n_4065));
OR2X1 g64874(.A (g3451), .B (n_10687), .Y (n_4062));
OR2X1 g64880(.A (g3802), .B (n_9091), .Y (n_4060));
AOI22X1 g64037(.A0 (n_2018), .A1 (n_3547), .B0 (n_523), .B1 (n_9693),.Y (n_4059));
NOR2X1 g64896(.A (n_3695), .B (n_8557), .Y (n_5701));
OR2X1 g64911(.A (g6494), .B (n_9398), .Y (n_4056));
OR2X1 g64913(.A (g5802), .B (n_9398), .Y (n_4055));
OR4X1 g62899(.A (n_11080), .B (n_4053), .C (n_9856), .D (g_22306), .Y(n_4054));
XOR2X1 g62928(.A (g4593), .B (n_10395), .Y (n_4050));
AOI21X1 g65011(.A0 (g4473), .A1 (n_2861), .B0 (g4459), .Y (n_4049));
MX2X1 g62938(.A (g2848), .B (n_3500), .S0 (n_8955), .Y (n_4048));
NAND4X1 g65041(.A (g5112), .B (n_9521), .C (g_11037), .D (g9553), .Y(n_4046));
AOI21X1 g65051(.A0 (g4164), .A1 (g4253), .B0 (n_3701), .Y (n_4247));
DFFSRX1 g4455_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g4456), .Q (), .QN (g4455));
DFFSRX1 g802_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12184), .Q (g_17653), .QN ());
NAND2X1 g61916(.A (n_4045), .B (g_14342), .Y (n_4578));
DFFSRX1 g728_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3671), .Q (g_12433), .QN ());
AND2X1 g65267(.A (n_11012), .B (n_10078), .Y (n_4044));
NOR2X1 g65289(.A (g2815), .B (g2724), .Y (n_4043));
NOR2X1 g65297(.A (g2783), .B (g2724), .Y (n_4042));
AOI22X1 g64033(.A0 (n_2007), .A1 (n_10948), .B0 (n_10660), .B1(n_10078), .Y (n_4040));
NAND3X1 g64010(.A (n_10672), .B (n_4038), .C (g2287), .Y (n_4281));
DFFSRX1 g518_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3723), .Q (g_14843), .QN ());
NOR2X1 g65747(.A (n_4231), .B (g2775), .Y (n_4037));
NAND2X1 g65781(.A (g1677), .B (n_4231), .Y (n_4035));
NAND2X1 g65853(.A (n_4231), .B (n_9952), .Y (n_4034));
NOR2X1 g65923(.A (g2715), .B (g2807), .Y (n_4033));
NAND2X1 g65936(.A (g2236), .B (n_4231), .Y (n_4032));
INVX1 g61003(.A (n_4030), .Y (n_4031));
OAI21X1 g63193(.A0 (n_3479), .A1 (g4153), .B0 (n_9627), .Y (n_4029));
NAND3X1 g63209(.A (n_11080), .B (g_22306), .C (n_9698), .Y (n_4028));
NAND3X1 g63210(.A (n_4024), .B (n_3660), .C (n_9651), .Y (n_4025));
NAND2X1 g63225(.A (n_3656), .B (n_1434), .Y (n_4022));
NOR2X1 g63227(.A (g5694), .B (n_10660), .Y (n_4021));
NOR2X1 g63229(.A (g6040), .B (n_11201), .Y (n_4020));
NOR2X1 g63230(.A (g6386), .B (g6395), .Y (n_4019));
NOR2X1 g63237(.A (g6732), .B (n_523), .Y (n_4018));
NOR2X1 g61007(.A (n_3778), .B (n_2172), .Y (n_4017));
AND2X1 g63247(.A (n_3172), .B (g5348), .Y (n_4016));
NOR2X1 g63251(.A (n_2882), .B (g5694), .Y (n_4015));
NOR2X1 g63253(.A (n_2613), .B (g6040), .Y (n_4014));
OAI21X1 g63255(.A0 (n_2150), .A1 (n_9978), .B0 (n_3653), .Y (n_4013));
NOR2X1 g63257(.A (n_2607), .B (g6386), .Y (n_4012));
NOR2X1 g63259(.A (n_2872), .B (g6732), .Y (n_4011));
AOI21X1 g63268(.A0 (n_2987), .A1 (n_286), .B0 (n_11081), .Y (n_4202));
DFFSRX1 g1418_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3647), .Q (g17320), .QN ());
DFFSRX1 g1384_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3666), .Q (g1384), .QN ());
OAI22X1 g63327(.A0 (n_4939), .A1 (n_3432), .B0 (n_2583), .B1(n_9627), .Y (n_4010));
MX2X1 g63346(.A (g4172), .B (n_3480), .S0 (n_9091), .Y (n_4009));
MX2X1 g63365(.A (g_15287), .B (n_3521), .S0 (n_9359), .Y (n_4008));
DFFSRX1 g66_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3636), .Q (g18881), .QN ());
AOI21X1 g63470(.A0 (n_10915), .A1 (n_3789), .B0 (g1728), .Y (n_4006));
NAND3X1 g63473(.A (n_1097), .B (n_10347), .C (n_10063), .Y (n_4005));
NAND3X1 g63478(.A (n_1098), .B (n_10473), .C (n_9209), .Y (n_4002));
NAND3X1 g63481(.A (n_1269), .B (n_10445), .C (n_9359), .Y (n_4000));
AOI21X1 g63483(.A0 (n_6676), .A1 (n_3782), .B0 (g1862), .Y (n_3998));
NAND3X1 g63485(.A (n_1099), .B (n_3455), .C (n_10385), .Y (n_3997));
NAND3X1 g63488(.A (n_3640), .B (n_1285), .C (n_11056), .Y (n_4805));
NAND2X1 g63499(.A (g4423), .B (n_10385), .Y (n_4170));
NAND2X1 g63505(.A (g4423), .B (n_9952), .Y (n_3996));
AOI22X1 g61021(.A0 (n_3460), .A1 (n_9627), .B0 (n_3372), .B1(n_3459), .Y (n_3995));
AOI22X1 g63542(.A0 (n_540), .A1 (n_7242), .B0 (n_7245), .B1 (g5138),.Y (n_3993));
DFFSRX1 g753_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3700), .Q (g_22034), .QN ());
AOI22X1 g63549(.A0 (n_600), .A1 (n_3455), .B0 (n_3814), .B1 (g6523),.Y (n_3992));
OAI22X1 g63555(.A0 (n_2748), .A1 (n_9193), .B0 (n_3410), .B1(n_9627), .Y (n_3991));
NAND4X1 g63557(.A (n_2145), .B (n_2144), .C (n_3269), .D (n_2332), .Y(n_3990));
NAND4X1 g63566(.A (n_2128), .B (n_2126), .C (n_3266), .D (n_2029), .Y(n_11189));
NAND4X1 g63569(.A (n_7018), .B (n_3984), .C (g5052), .D (n_10697), .Y(n_3985));
MX2X1 g63570(.A (g5128), .B (n_168), .S0 (n_7245), .Y (n_3983));
AOI21X1 g63633(.A0 (n_3618), .A1 (n_9193), .B0 (n_3642), .Y (n_3982));
MX2X1 g63648(.A (n_10813), .B (n_3449), .S0 (n_8955), .Y (n_3981));
OAI21X1 g62267(.A0 (n_3537), .A1 (n_9599), .B0 (n_3709), .Y (n_3979));
AOI21X1 g61215(.A0 (n_11211), .A1 (g1589), .B0 (n_3870), .Y (n_3978));
AOI21X1 g61220(.A0 (n_10763), .A1 (g1589), .B0 (n_10762), .Y(n_3977));
XOR2X1 g63763(.A (n_3011), .B (n_10347), .Y (n_3974));
XOR2X1 g63764(.A (n_2684), .B (n_10473), .Y (n_3973));
XOR2X1 g63765(.A (n_2704), .B (n_10445), .Y (n_3972));
XOR2X1 g63768(.A (n_3007), .B (n_3455), .Y (n_3971));
NAND3X1 g61037(.A (n_3369), .B (n_2555), .C (n_3523), .Y (n_3970));
MX2X1 g61223(.A (g1589), .B (n_649), .S0 (n_8955), .Y (n_3969));
MX2X1 g63791(.A (n_1285), .B (n_3429), .S0 (n_8955), .Y (n_3968));
MX2X1 g63792(.A (g_17065), .B (n_3424), .S0 (n_8955), .Y (n_3966));
MX2X1 g63793(.A (n_3550), .B (n_3423), .S0 (n_9156), .Y (n_3964));
MX2X1 g63797(.A (g_19113), .B (n_3422), .S0 (n_9091), .Y (n_3963));
MX2X1 g63799(.A (g_16677), .B (n_3420), .S0 (n_9000), .Y (n_3962));
MX2X1 g63800(.A (g_21720), .B (n_3418), .S0 (n_9000), .Y (n_3960));
MX2X1 g63801(.A (g_13758), .B (n_3417), .S0 (n_9000), .Y (n_3959));
MX2X1 g63802(.A (g_19289), .B (n_3416), .S0 (n_9311), .Y (n_3958));
MX2X1 g63807(.A (g_21778), .B (n_3415), .S0 (n_9797), .Y (n_3957));
INVX1 g63880(.A (n_7025), .Y (n_3956));
OR2X1 g63882(.A (n_3615), .B (n_9775), .Y (n_3955));
INVX1 g63887(.A (n_7102), .Y (n_3953));
INVX1 g63890(.A (n_8628), .Y (n_3952));
INVX1 g63897(.A (n_8633), .Y (n_3951));
NOR2X1 g63915(.A (n_3948), .B (n_10917), .Y (n_3949));
NAND2X1 g63925(.A (n_4424), .B (n_9358), .Y (n_5007));
NOR2X1 g63938(.A (n_3557), .B (n_9193), .Y (n_3947));
NOR2X1 g63956(.A (n_3574), .B (n_3945), .Y (n_3946));
NOR3X1 g63972(.A (n_6752), .B (n_3943), .C (g2070), .Y (n_3944));
NAND4X1 g63983(.A (n_3561), .B (n_2918), .C (n_10063), .D (n_3065),.Y (n_3942));
NAND4X1 g63994(.A (n_3560), .B (n_2917), .C (n_9750), .D (n_3062), .Y(n_3941));
DFFSRX1 g1345_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3689), .Q (g1345), .QN ());
NAND3X1 g64011(.A (n_10672), .B (g2331), .C (n_386), .Y (n_4279));
NAND3X1 g64012(.A (n_10675), .B (g2361), .C (g2287), .Y (n_4277));
NAND3X1 g64013(.A (n_10672), .B (n_4038), .C (g2361), .Y (n_4275));
NAND3X1 g64014(.A (n_10854), .B (n_3939), .C (g2421), .Y (n_4273));
NAND3X1 g64015(.A (n_10854), .B (g2465), .C (n_437), .Y (n_4271));
NAND3X1 g64016(.A (n_10857), .B (n_4339), .C (g2421), .Y (n_4269));
NAND3X1 g64017(.A (n_10854), .B (n_3939), .C (n_4339), .Y (n_4267));
DFFSRX1 g661_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3673), .Q (g_20073), .QN ());
DFFSRX1 g1129_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3585), .Q (g_20563), .QN ());
DFFSRX1 g4669_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3620), .Q (g4669), .QN ());
OR2X1 g64022(.A (n_3938), .B (n_5471), .Y (n_4539));
DFFSRX1 g4859_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3725), .Q (n_11216), .QN ());
AOI22X1 g64032(.A0 (n_2588), .A1 (n_3399), .B0 (n_8806), .B1(n_9193), .Y (n_3937));
AOI22X1 g64036(.A0 (n_2015), .A1 (n_3626), .B0 (g6395), .B1(n_10078), .Y (n_3936));
DFFSRX1 g4793_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3721), .Q (g4793), .QN ());
DFFSRX1 g650_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3675), .Q (g_18795), .QN ());
DFFSRX1 g655_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3674), .Q (g_22038), .QN ());
DFFSRX1 g681_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3670), .Q (g_17934), .QN ());
DFFSRX1 g718_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3672), .Q (g_18238), .QN ());
DFFSRX1 g4983_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3688), .Q (g4983), .QN ());
DFFSRX1 g1002_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3662), .Q (g_19911), .QN ());
DFFSRX1 g4633_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3655), .Q (g4633), .QN ());
DFFSRX1 g1046_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3638), .Q (g_18739), .QN ());
DFFSRX1 g4888_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3622), .Q (g4888), .QN ());
DFFSRX1 g499_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3621), .Q (g_19789), .QN ());
OAI21X1 g64072(.A0 (n_3779), .A1 (n_6978), .B0 (n_3598), .Y (n_3934));
DFFSRX1 g370_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3555), .Q (g_5029), .QN ());
DFFSRX1 g1448_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3591), .Q (g1448), .QN ());
DFFSRX1 g5029_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3577), .Q (g5029), .QN ());
DFFSRX1 g504_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3554), .Q (g_18996), .QN ());
DFFSRX1 g4836_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3722), .Q (g34034), .QN ());
DFFSRX1 g513_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3552), .Q (g_22021), .QN ());
DFFSRX1 g2975_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3724), .Q (g2975), .QN ());
DFFSRX1 g4621_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3546), .Q (g4621), .QN ());
DFFSRX1 g5535_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3712), .Q (g5535), .QN ());
DFFSRX1 g6573_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3711), .Q (g6573), .QN ());
DFFSRX1 g3530_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3710), .Q (g3530), .QN ());
OAI21X1 g64080(.A0 (n_3775), .A1 (n_7003), .B0 (n_3592), .Y (n_3933));
NAND2X1 g60954(.A (n_3658), .B (n_3716), .Y (n_3932));
INVX1 g64177(.A (n_10944), .Y (n_3929));
INVX2 g64187(.A (n_6759), .Y (n_4304));
INVX2 g64199(.A (n_3925), .Y (n_4668));
INVX1 g64240(.A (n_4447), .Y (n_3922));
OAI21X1 g62599(.A0 (n_3915), .A1 (n_3914), .B0 (n_3913), .Y (n_3916));
INVX1 g64330(.A (n_10380), .Y (n_4299));
OR4X1 g60959(.A (n_10429), .B (n_3910), .C (n_9856), .D (g1367), .Y(n_3911));
OAI21X1 g64397(.A0 (g16693), .A1 (g14518), .B0 (n_3535), .Y (n_3907));
AOI21X1 g62650(.A0 (n_3718), .A1 (n_28), .B0 (n_11032), .Y (n_3906));
MX2X1 g64408(.A (g_21318), .B (g14201), .S0 (n_5582), .Y (n_3905));
NAND4X1 g62673(.A (n_3646), .B (n_6577), .C (n_10687), .D (g4332), .Y(n_3904));
NAND3X1 g64532(.A (g5752), .B (n_9521), .C (g_7062), .Y (n_3903));
NAND3X1 g64582(.A (g3401), .B (n_9521), .C (g_5313), .Y (n_3902));
INVX1 g64596(.A (n_3900), .Y (n_6364));
NAND3X1 g64664(.A (n_3732), .B (g3965), .C (n_8917), .Y (n_11219));
NOR2X1 g64679(.A (n_3897), .B (n_3896), .Y (n_3898));
NAND4X1 g64732(.A (g3905), .B (n_3894), .C (g16693), .D (n_6808), .Y(n_3895));
AOI21X1 g61821(.A0 (n_1885), .A1 (n_2845), .B0 (n_3775), .Y (n_3893));
AOI21X1 g61822(.A0 (n_1884), .A1 (n_2844), .B0 (n_3779), .Y (n_3891));
DFFSRX1 g875_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14201), .Q (g14217), .QN ());
NAND2X1 g62833(.A (n_3321), .B (n_3516), .Y (n_3886));
INVX1 g62837(.A (n_11031), .Y (n_3885));
OR2X1 g64855(.A (g5456), .B (n_9091), .Y (n_3883));
NAND3X1 g64930(.A (n_6967), .B (n_9553), .C (g_11037), .Y (n_3882));
AOI22X1 g62909(.A0 (n_3331), .A1 (n_10184), .B0 (n_11134), .B1(n_9107), .Y (n_3881));
AOI22X1 g65024(.A0 (g2960), .A1 (n_3356), .B0 (g2970), .B1 (g2975),.Y (n_3879));
AOI22X1 g65032(.A0 (g2922), .A1 (n_3357), .B0 (g2912), .B1 (n_3463),.Y (n_3878));
MX2X1 g62940(.A (n_3501), .B (n_3330), .S0 (n_9167), .Y (n_3877));
DFFSRX1 g1395_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3407), .Q (g1395), .QN ());
DFFSRX1 g4659_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3412), .Q (g4659), .QN ());
DFFSRX1 g5109_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9497), .Q (), .QN (g5109));
NAND2X1 g65266(.A (n_3868), .B (n_9019), .Y (n_3869));
DFFSRX1 g4358_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3414), .Q (n_1627), .QN ());
NOR2X1 g65336(.A (n_10650), .B (n_3868), .Y (n_3866));
NAND2X1 g65810(.A (g1811), .B (n_3679), .Y (n_3863));
DFFSRX1 g4366_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3494), .Q (), .QN (g4366));
INVX1 g61439(.A (g1246), .Y (n_4558));
OR2X1 g61004(.A (n_3860), .B (g7946), .Y (n_4030));
NOR2X1 g61005(.A (n_3860), .B (n_10196), .Y (n_3861));
OAI21X1 g63212(.A0 (n_2425), .A1 (n_10115), .B0 (n_3488), .Y(n_3859));
NAND2X1 g63214(.A (n_3517), .B (n_3857), .Y (n_3858));
NOR2X1 g63234(.A (n_8836), .B (n_3855), .Y (n_3856));
NOR2X1 g63240(.A (n_8836), .B (n_8832), .Y (n_3854));
NAND4X1 g63261(.A (n_3050), .B (n_3302), .C (n_3049), .D (n_3032), .Y(n_3852));
NAND4X1 g63271(.A (n_3845), .B (n_10063), .C (n_3844), .D (n_2428),.Y (n_3851));
NOR2X1 g61009(.A (n_3860), .B (n_3849), .Y (n_4284));
NAND3X1 g61010(.A (n_3484), .B (g1361), .C (n_9811), .Y (n_3848));
OAI21X1 g63283(.A0 (n_3894), .A1 (n_9940), .B0 (n_3487), .Y (n_3847));
NAND4X1 g63285(.A (n_3845), .B (n_3844), .C (n_9279), .D (n_40), .Y(n_3846));
DFFSRX1 g4933_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3468), .Q (g4933), .QN ());
NAND4X1 g63314(.A (n_4832), .B (n_6767), .C (n_9279), .D (n_416), .Y(n_3843));
AOI21X1 g63332(.A0 (g1183), .A1 (n_8837), .B0 (n_3505), .Y (n_3841));
NAND3X1 g62101(.A (n_2278), .B (n_2711), .C (n_3327), .Y (n_3840));
OAI21X1 g63345(.A0 (g2864), .A1 (n_9894), .B0 (n_3503), .Y (n_3839));
AOI21X1 g61499(.A0 (n_3838), .A1 (g1242), .B0 (n_3837), .Y (n_5057));
INVX1 g63374(.A (g5694), .Y (n_3836));
INVX1 g63376(.A (g6040), .Y (n_3835));
INVX1 g63378(.A (g6386), .Y (n_3834));
INVX1 g63380(.A (g6732), .Y (n_3833));
NAND3X1 g63460(.A (n_1101), .B (n_7243), .C (n_9894), .Y (n_3830));
OR2X1 g63487(.A (n_10532), .B (n_3639), .Y (n_3828));
NOR2X1 g63511(.A (n_2755), .B (n_3478), .Y (n_3826));
NAND3X1 g63517(.A (n_10768), .B (n_2638), .C (n_3264), .Y (n_3825));
NAND3X1 g63521(.A (n_3482), .B (g_16958), .C (n_9493), .Y (n_3824));
NAND3X1 g63533(.A (n_3426), .B (n_3822), .C (n_3438), .Y (n_3823));
AOI22X1 g63536(.A0 (n_3260), .A1 (n_8676), .B0 (n_599), .B1 (n_3259),.Y (n_3821));
NAND4X1 g63562(.A (n_6577), .B (n_3645), .C (n_662), .D (n_3213), .Y(n_3819));
NAND4X1 g63564(.A (n_1849), .B (n_3278), .C (n_1858), .D (n_1574), .Y(n_3817));
NAND4X1 g63568(.A (n_10770), .B (n_3984), .C (n_9359), .D (g5046), .Y(n_3816));
MX2X1 g63597(.A (g6513), .B (n_158), .S0 (n_3814), .Y (n_3815));
AOI22X1 g63638(.A0 (n_3604), .A1 (n_9772), .B0 (n_3814), .B1(n_3812), .Y (n_3813));
DFFSRX1 g5881_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3532), .Q (g5881), .QN ());
AOI21X1 g61033(.A0 (n_3366), .A1 (n_2178), .B0 (n_3459), .Y (n_3811));
OAI22X1 g62298(.A0 (n_3346), .A1 (n_3720), .B0 (n_8637), .B1(n_9830), .Y (n_3810));
XOR2X1 g63762(.A (n_2718), .B (n_7242), .Y (n_3809));
DFFSRX1 g5499_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3408), .Q (g5499), .QN ());
MX2X1 g63809(.A (n_6967), .B (n_3271), .S0 (n_9234), .Y (n_3808));
AOI21X1 g63883(.A0 (g2932), .A1 (n_27), .B0 (n_9976), .Y (n_3807));
NOR2X1 g63912(.A (n_10347), .B (n_6399), .Y (n_3803));
NOR2X1 g63916(.A (n_10473), .B (n_6398), .Y (n_3802));
NOR2X1 g63920(.A (n_10445), .B (n_6406), .Y (n_3801));
NOR3X1 g63921(.A (n_10078), .B (g5046), .C (n_10770), .Y (n_3800));
NOR2X1 g63939(.A (n_3538), .B (n_3797), .Y (n_3798));
NAND2X1 g63953(.A (n_4843), .B (n_9493), .Y (n_4956));
MX2X1 g61652(.A (g_20614), .B (n_10752), .S0 (n_9750), .Y (n_3795));
NAND2X1 g63966(.A (n_3427), .B (n_3017), .Y (n_3793));
AOI21X1 g63980(.A0 (n_3244), .A1 (n_11037), .B0 (n_10621), .Y(n_3792));
NAND3X1 g63981(.A (n_10915), .B (n_3789), .C (g1728), .Y (n_4220));
NAND3X1 g63982(.A (n_10915), .B (g1772), .C (n_446), .Y (n_4218));
NAND3X1 g63984(.A (n_10915), .B (n_4139), .C (g1728), .Y (n_4216));
AOI21X1 g63985(.A0 (n_10947), .A1 (n_4982), .B0 (n_7150), .Y(n_3788));
AOI21X1 g63986(.A0 (n_3612), .A1 (n_4980), .B0 (n_10506), .Y(n_3786));
AOI21X1 g63987(.A0 (n_3784), .A1 (n_4978), .B0 (n_3277), .Y (n_3785));
NAND3X1 g63988(.A (n_6676), .B (n_3782), .C (g1862), .Y (n_4211));
NAND3X1 g63989(.A (n_6676), .B (g1936), .C (g1862), .Y (n_4207));
AOI21X1 g63990(.A0 (n_3605), .A1 (n_11070), .B0 (n_3275), .Y(n_3781));
NAND3X1 g63991(.A (n_6676), .B (n_3782), .C (g1936), .Y (n_4203));
NAND3X1 g63992(.A (n_6676), .B (g1906), .C (n_328), .Y (n_4209));
AOI21X1 g63993(.A0 (n_3779), .A1 (g3639), .B0 (n_1273), .Y (n_3780));
INVX1 g61047(.A (n_3778), .Y (n_4242));
AOI21X1 g64000(.A0 (n_6243), .A1 (g3990), .B0 (n_6787), .Y (n_3777));
AOI21X1 g64003(.A0 (n_3775), .A1 (n_10834), .B0 (n_8586), .Y(n_3776));
NAND3X1 g64009(.A (n_10915), .B (n_3789), .C (n_4139), .Y (n_4214));
DFFSRX1 g1404_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3483), .Q (g1404), .QN ());
DFFSRX1 g1105_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3454), .Q (g_16456), .QN ());
DFFSRX1 g956_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3458), .Q (g_18869), .QN ());
DFFSRX1 g4664_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3520), .Q (g4664), .QN ());
NAND3X1 g64031(.A (n_3440), .B (n_659), .C (n_9398), .Y (n_3774));
DFFSRX1 g1554_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3508), .Q (g1554), .QN ());
DFFSRX1 g4854_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3507), .Q (g4854), .QN ());
DFFSRX1 g4849_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3529), .Q (g4849), .QN ());
DFFSRX1 g3343_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3512), .Q (), .QN (g3343));
DFFSRX1 g3694_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3511), .Q (), .QN (g3694));
MX2X1 g64062(.A (g5069), .B (n_2044), .S0 (n_9448), .Y (n_3771));
DFFSRX1 g645_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3496), .Q (g_22464), .QN ());
DFFSRX1 g4653_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3490), .Q (g4653), .QN ());
DFFSRX1 g4064_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3481), .Q (g4064), .QN ());
DFFSRX1 g2848_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3473), .Q (g2848), .QN ());
DFFSRX1 g4743_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3470), .Q (g4743), .QN ());
DFFSRX1 g4754_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3469), .Q (g4754), .QN ());
DFFSRX1 g4698_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3471), .Q (g4698), .QN ());
DFFSRX1 g4843_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3475), .Q (g4843), .QN ());
DFFSRX1 g4765_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3510), .Q (g4765), .QN ());
DFFSRX1 g4955_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3465), .Q (g4955), .QN ());
DFFSRX1 g4944_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3466), .Q (g4944), .QN ());
DFFSRX1 g5313_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3437), .Q (g_4409), .QN ());
DFFSRX1 g5659_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3436), .Q (g_3381), .QN ());
DFFSRX1 g6005_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3435), .Q (n_11050), .QN ());
DFFSRX1 g6351_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3434), .Q (g_6165), .QN ());
DFFSRX1 g1300_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3461), .Q (g1300), .QN ());
DFFSRX1 g6697_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3433), .Q (g_8864), .QN ());
DFFSRX1 g667_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3413), .Q (g_10278), .QN ());
DFFSRX1 g3494_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3402), .Q (g3494), .QN ());
DFFSRX1 g6537_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3403), .Q (g6537), .QN ());
DFFSRX1 g3845_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3400), .Q (g3845), .QN ());
XOR2X1 g64076(.A (n_3769), .B (n_6243), .Y (n_3770));
DFFSRX1 g3143_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3404), .Q (g3143), .QN ());
DFFSRX1 g6191_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3395), .Q (g6191), .QN ());
DFFSRX1 g5188_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3534), .Q (g5188), .QN ());
DFFSRX1 g6227_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3531), .Q (g6227), .QN ());
OAI22X1 g64078(.A0 (n_1557), .A1 (n_9599), .B0 (g4284), .B1 (n_9811),.Y (n_3767));
DFFSRX1 g3179_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3533), .Q (g3179), .QN ());
DFFSRX1 g3881_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3530), .Q (g3881), .QN ());
DFFSRX1 g4467_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3518), .Q (g4467), .QN ());
OAI21X1 g64091(.A0 (n_3765), .A1 (n_9311), .B0 (n_3464), .Y (n_3766));
DFFSRX1 g3672_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16924), .Q (g13881), .QN ());
DFFSRX1 g3321_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16874), .Q (g13865), .QN ());
OR2X1 g64137(.A (g3106), .B (n_10943), .Y (n_6051));
OR2X1 g64148(.A (g3457), .B (n_3758), .Y (n_6052));
NAND2X1 g64170(.A (n_3543), .B (n_2653), .Y (n_3764));
NAND4X1 g64184(.A (g3550), .B (n_4682), .C (g14451), .D (n_10883), .Y(n_3761));
INVX1 g64200(.A (n_4424), .Y (n_3925));
BUFX3 g64203(.A (n_4424), .Y (n_4494));
BUFX3 g64204(.A (n_4424), .Y (n_4499));
BUFX3 g64205(.A (n_4424), .Y (n_4482));
BUFX3 g64209(.A (n_4424), .Y (n_4497));
NAND2X1 g64241(.A (n_2996), .B (n_3758), .Y (n_4447));
NAND3X1 g64271(.A (n_3775), .B (g4939), .C (n_9664), .Y (n_3755));
NAND3X1 g64272(.A (n_3779), .B (g4950), .C (n_9717), .Y (n_3753));
NAND3X1 g64273(.A (n_6243), .B (g4961), .C (n_10063), .Y (n_3752));
NOR2X1 g64317(.A (n_2014), .B (n_3775), .Y (n_3746));
INVX1 g64320(.A (n_3571), .Y (n_3745));
NOR2X1 g64325(.A (n_2016), .B (n_3779), .Y (n_3744));
NOR2X1 g64337(.A (n_2009), .B (n_6243), .Y (n_3742));
INVX4 g64345(.A (n_5471), .Y (n_4108));
NAND4X1 g64377(.A (n_10576), .B (g3538), .C (g14451), .D (n_10894),.Y (n_3740));
OAI22X1 g62680(.A0 (n_3314), .A1 (n_3687), .B0 (n_598), .B1 (n_9627),.Y (n_3738));
DFFSRX1 g4019_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14518), .Q (g16955), .QN ());
NAND3X1 g64529(.A (g5406), .B (n_9091), .C (g_5508), .Y (n_3737));
NAND3X1 g64535(.A (g3050), .B (n_9091), .C (g_6579), .Y (n_3736));
NAND3X1 g64543(.A (g6098), .B (n_9521), .C (g_14965), .Y (n_3735));
NAND3X1 g64545(.A (g6444), .B (n_9553), .C (g_3861), .Y (n_3734));
NAND3X1 g64558(.A (g3752), .B (n_9521), .C (g_5156), .Y (n_3733));
DFFSRX1 g5845_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3406), .Q (g5845), .QN ());
AND2X1 g64565(.A (n_3732), .B (n_8917), .Y (n_4096));
NOR2X1 g64577(.A (n_3730), .B (n_3896), .Y (n_3731));
NOR2X1 g64578(.A (n_3728), .B (n_3896), .Y (n_3729));
NOR2X1 g64581(.A (n_3726), .B (n_3896), .Y (n_3727));
INVX1 g64597(.A (n_6005), .Y (n_3900));
CLKBUFX1 g64598(.A (n_6005), .Y (n_6334));
NAND3X1 g61796(.A (n_2809), .B (n_2234), .C (n_3074), .Y (n_3725));
DFFSRX1 g1559_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3255), .Q (n_10113), .QN ());
OAI21X1 g64691(.A0 (g2965), .A1 (n_9311), .B0 (n_3377), .Y (n_3724));
OAI21X1 g64697(.A0 (n_2884), .A1 (n_2497), .B0 (n_3370), .Y (n_3723));
INVX1 g64760(.A (n_3540), .Y (n_3722));
NAND2X1 g62810(.A (n_3915), .B (n_3914), .Y (n_3913));
NOR2X1 g62823(.A (n_3257), .B (n_3720), .Y (n_3721));
NAND4X1 g62849(.A (n_3351), .B (n_8913), .C (n_10013), .D (n_10823),.Y (n_3717));
NAND3X1 g60979(.A (n_10005), .B (n_3059), .C (n_2252), .Y (n_3716));
XOR2X1 g62905(.A (n_640), .B (n_3713), .Y (n_3715));
OAI21X1 g64972(.A0 (n_1388), .A1 (n_9443), .B0 (n_3360), .Y (n_3712));
OAI21X1 g64974(.A0 (n_1375), .A1 (n_9903), .B0 (n_3361), .Y (n_3711));
OAI21X1 g64976(.A0 (n_1369), .A1 (n_9129), .B0 (n_3362), .Y (n_3710));
AOI21X1 g62929(.A0 (n_3707), .A1 (n_9836), .B0 (n_3352), .Y (n_3709));
OAI21X1 g62930(.A0 (n_3651), .A1 (n_3707), .B0 (n_3350), .Y (n_3708));
DFFSRX1 g1489_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3382), .Q (g1489), .QN ());
DFFSRX1 g1216_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3263), .Q (n_10120), .QN ());
AOI22X1 g64035(.A0 (n_2011), .A1 (n_5459), .B0 (n_11201), .B1(n_9193), .Y (n_3706));
INVX1 g65122(.A (g_7062), .Y (g9680));
INVX1 g65130(.A (g_5313), .Y (g8342));
DFFSRX1 g3451_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8279), .Q (), .QN (g3451));
DFFSRX1 g5802_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9617), .Q (), .QN (g5802));
DFFSRX1 g3802_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8344), .Q (), .QN (g3802));
DFFSRX1 g4459_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3353), .Q (g4459), .QN ());
DFFSRX1 g6494_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9743), .Q (), .QN (g6494));
OAI22X1 g61386(.A0 (n_3075), .A1 (n_1985), .B0 (n_129), .B1 (n_9466),.Y (n_3703));
DFFSRX1 g3100_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8215), .Q (), .QN (g3100));
DFFSRX1 g6148_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9682), .Q (), .QN (g6148));
NAND4X1 g60988(.A (n_6735), .B (n_4866), .C (n_9359), .D (n_297), .Y(n_3702));
NOR2X1 g65349(.A (g4145), .B (g4253), .Y (n_3701));
DFFSRX1 g6727_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3292), .Q (n_11186), .QN ());
MX2X1 g63083(.A (g_18793), .B (n_3058), .S0 (n_9218), .Y (n_3700));
DFFSRX1 g3698_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3261), .Q (g3698), .QN ());
DFFSRX1 g2741_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3344), .Q (n_11013), .QN ());
DFFSRX1 g4456_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3341), .Q (g4456), .QN ());
DFFSRX1 g799_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3336), .Q (g12184), .QN ());
INVX1 g65715(.A (n_3697), .Y (n_5704));
NOR2X1 g65755(.A (n_3679), .B (n_8895), .Y (n_5705));
INVX1 g65867(.A (n_3695), .Y (n_5702));
DFFSRX1 g1246_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3345), .Q (g1246), .QN ());
NOR2X1 g63192(.A (n_3325), .B (n_2437), .Y (n_3693));
XOR2X1 g61053(.A (n_1591), .B (n_3628), .Y (n_3692));
AND2X1 g63213(.A (n_3690), .B (g_10715), .Y (n_3691));
NAND3X1 g61006(.A (n_3312), .B (n_2268), .C (n_2875), .Y (n_3689));
NOR2X1 g63241(.A (n_3381), .B (n_3687), .Y (n_3688));
OAI21X1 g63260(.A0 (n_3431), .A1 (g_19414), .B0 (n_3334), .Y(n_3686));
AOI21X1 g63262(.A0 (n_3323), .A1 (n_1540), .B0 (n_3324), .Y (n_3685));
NAND4X1 g63270(.A (n_3329), .B (n_10188), .C (n_9894), .D (n_551), .Y(n_3683));
AOI21X1 g63302(.A0 (n_3234), .A1 (n_3439), .B0 (n_1417), .Y (n_3681));
AOI22X1 g63320(.A0 (n_2304), .A1 (n_3491), .B0 (n_1734), .B1(n_9627), .Y (n_3680));
INVX1 g66266(.A (n_3679), .Y (n_4231));
OAI21X1 g63331(.A0 (n_3563), .A1 (n_11134), .B0 (n_3328), .Y(n_3677));
MX2X1 g63358(.A (g_14265), .B (n_3175), .S0 (n_9000), .Y (n_3675));
MX2X1 g63359(.A (g_18795), .B (n_3043), .S0 (n_8955), .Y (n_3674));
MX2X1 g63360(.A (n_10103), .B (n_3038), .S0 (n_8955), .Y (n_3673));
MX2X1 g63363(.A (n_3042), .B (n_3040), .S0 (n_8955), .Y (n_3672));
MX2X1 g63364(.A (g_20073), .B (n_3041), .S0 (n_9279), .Y (n_3671));
MX2X1 g63369(.A (g_22464), .B (n_3034), .S0 (n_9156), .Y (n_3670));
DFFSRX1 g5348_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3300), .Q (g5348), .QN ());
DFFSRX1 g5694_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3319), .Q (), .QN (g5694));
DFFSRX1 g6040_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3299), .Q (), .QN (g6040));
DFFSRX1 g6386_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3298), .Q (), .QN (g6386));
DFFSRX1 g6732_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3296), .Q (), .QN (g6732));
NAND3X1 g61052(.A (n_3373), .B (n_2283), .C (n_3187), .Y (n_3666));
AOI21X1 g61515(.A0 (n_10323), .A1 (g23683), .B0 (n_10321), .Y(n_4743));
NAND3X1 g63479(.A (n_3305), .B (n_2285), .C (n_2885), .Y (n_3662));
NAND3X1 g63489(.A (n_3661), .B (n_3660), .C (g_18793), .Y (n_4024));
NOR2X1 g63493(.A (n_3477), .B (n_2043), .Y (n_3659));
AOI22X1 g61020(.A0 (n_2253), .A1 (n_10330), .B0 (g1532), .B1(n_9772), .Y (n_3658));
AOI22X1 g63537(.A0 (n_3014), .A1 (n_8639), .B0 (n_607), .B1 (n_3013),.Y (n_3656));
NAND3X1 g63539(.A (n_2746), .B (n_2545), .C (n_3027), .Y (n_3655));
OR2X1 g63550(.A (n_3309), .B (n_3915), .Y (n_3654));
AOI22X1 g63559(.A0 (n_3029), .A1 (n_9501), .B0 (n_2657), .B1(n_3323), .Y (n_3653));
DFFSRX1 g385_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3320), .Q (g_20951), .QN ());
NAND4X1 g62251(.A (n_3333), .B (n_3651), .C (n_9834), .D (n_10818),.Y (n_3652));
XOR2X1 g63644(.A (n_662), .B (n_3258), .Y (n_3648));
NOR2X1 g61038(.A (n_3288), .B (n_961), .Y (n_3647));
DFFSRX1 g4423_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g10306), .Q (g4423), .QN ());
NAND2X1 g63889(.A (n_3645), .B (n_662), .Y (n_3646));
NOR2X1 g63907(.A (n_7243), .B (n_3641), .Y (n_3642));
INVX1 g63950(.A (n_3639), .Y (n_3640));
NAND2X1 g63970(.A (n_3247), .B (n_3015), .Y (n_3638));
NAND3X1 g63979(.A (n_6970), .B (n_2364), .C (n_3218), .Y (n_3637));
INVX1 g61048(.A (n_3860), .Y (n_3778));
DFFSRX1 g4294_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3359), .Q (g10122), .QN ());
DFFSRX1 g1306_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3348), .Q (g1306), .QN ());
DFFSRX1 g1052_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3347), .Q (g_18488), .QN ());
OAI21X1 g64040(.A0 (n_227), .A1 (n_9681), .B0 (n_3285), .Y (n_3636));
DFFSRX1 g5689_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3322), .Q (g5689), .QN ());
DFFSRX1 g996_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3317), .Q (g_20614), .QN ());
DFFSRX1 g1146_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3308), .Q (g_18902), .QN ());
DFFSRX1 g1135_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3279), .Q (g_11413), .QN ());
DFFSRX1 g3347_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3262), .Q (g3347), .QN ());
DFFSRX1 g4349_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3355), .Q (g4349), .QN ());
DFFSRX1 g1075_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3303), .Q (g17291), .QN ());
DFFSRX1 g5343_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3315), .Q (g5343), .QN ());
XOR2X1 g64065(.A (n_11201), .B (n_5459), .Y (n_3634));
DFFSRX1 g6381_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3313), .Q (g6381), .QN ());
DFFSRX1 g6035_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3301), .Q (g6035), .QN ());
DFFSRX1 g1041_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3273), .Q (n_2458), .QN ());
XOR2X1 g64066(.A (n_10660), .B (n_10948), .Y (n_3633));
DFFSRX1 g4646_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3274), .Q (g34026), .QN ());
DFFSRX1 g5152_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3290), .Q (g5152), .QN ());
DFFSRX1 g278_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3289), .Q (g_13838), .QN ());
XOR2X1 g64069(.A (n_8806), .B (g28753), .Y (n_3631));
DFFSRX1 g3111_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3254), .Q (g3111), .QN ());
DFFSRX1 g1472_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3283), .Q (g1472), .QN ());
DFFSRX1 g1478_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3282), .Q (g1478), .QN ());
DFFSRX1 g4628_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3270), .Q (g4628), .QN ());
XOR2X1 g61054(.A (g1333), .B (n_3628), .Y (n_3629));
DFFSRX1 g550_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3358), .Q (g_18015), .QN ());
XOR2X1 g64081(.A (n_3626), .B (g6395), .Y (n_3627));
DFFSRX1 g2763_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3335), .Q (g2763), .QN ());
DFFSRX1 g4057_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3337), .Q (g4057), .QN ());
DFFSRX1 g4087_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3339), .Q (g4087), .QN ());
DFFSRX1 g4141_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3340), .Q (g4141), .QN ());
DFFSRX1 g4417_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3343), .Q (g4417), .QN ());
XOR2X1 g64094(.A (n_3624), .B (n_10398), .Y (n_3625));
NOR2X1 g65313(.A (g3003), .B (n_9453), .Y (g21727));
MX2X1 g64101(.A (g4894), .B (n_3217), .S0 (n_9218), .Y (n_3622));
NOR2X1 g64134(.A (n_3389), .B (n_9775), .Y (n_3621));
NAND3X1 g61709(.A (n_2868), .B (n_2604), .C (n_3153), .Y (n_3620));
NOR2X1 g64161(.A (g2886), .B (g2946), .Y (n_3615));
NOR2X1 g64167(.A (g2946), .B (g2955), .Y (n_3614));
NAND3X1 g64168(.A (n_3612), .B (n_3611), .C (n_9894), .Y (n_3613));
NAND3X1 g64180(.A (n_3605), .B (n_3604), .C (n_9698), .Y (n_3606));
NAND2X1 g64182(.A (n_3775), .B (n_64), .Y (n_3603));
NAND2X2 g64210(.A (g4284), .B (n_10871), .Y (n_4424));
NAND2X1 g64212(.A (n_3779), .B (n_1818), .Y (n_3599));
NAND2X1 g64214(.A (n_3779), .B (n_6978), .Y (n_3598));
NAND2X1 g64227(.A (n_6243), .B (n_151), .Y (n_3593));
NAND2X1 g64228(.A (n_3775), .B (n_7003), .Y (n_3592));
NAND3X1 g64229(.A (n_3241), .B (n_2539), .C (n_2920), .Y (n_3591));
NAND3X1 g64234(.A (n_3784), .B (n_3589), .C (n_9811), .Y (n_3590));
NAND3X1 g64248(.A (n_8707), .B (g4704), .C (n_9448), .Y (n_3588));
NAND3X1 g61725(.A (n_3221), .B (n_2281), .C (n_3170), .Y (n_3585));
NAND3X1 g64252(.A (n_10947), .B (g4749), .C (n_9834), .Y (n_3582));
NAND3X1 g64254(.A (n_3612), .B (g4760), .C (n_9627), .Y (n_3581));
NAND3X1 g64255(.A (n_3784), .B (g4771), .C (n_10063), .Y (n_3580));
NAND3X1 g64270(.A (n_3605), .B (g4894), .C (n_9750), .Y (n_3578));
NAND2X1 g64280(.A (n_3189), .B (n_3387), .Y (n_3577));
INVX1 g62580(.A (n_3448), .Y (n_4045));
INVX1 g64303(.A (n_6676), .Y (n_3574));
INVX1 g64318(.A (n_3441), .Y (n_3572));
AOI21X1 g64321(.A0 (n_3569), .A1 (n_1285), .B0 (n_3390), .Y (n_3571));
AOI21X1 g64322(.A0 (n_3569), .A1 (g_12791), .B0 (n_3566), .Y(n_3570));
NAND3X1 g64329(.A (n_3566), .B (n_456), .C (n_9425), .Y (n_3567));
INVX2 g64347(.A (n_10270), .Y (n_5471));
NAND4X1 g62644(.A (n_3307), .B (n_3563), .C (n_9209), .D (n_684), .Y(n_3564));
OAI21X1 g64395(.A0 (g16624), .A1 (g14421), .B0 (n_3210), .Y (n_3561));
OAI21X1 g64396(.A0 (g16656), .A1 (g14451), .B0 (n_3209), .Y (n_3560));
INVX1 g61302(.A (g1589), .Y (n_4149));
MX2X1 g64406(.A (n_10568), .B (g14189), .S0 (n_5582), .Y (n_3559));
AOI22X1 g64417(.A0 (n_3003), .A1 (g_21576), .B0 (n_3569), .B1(n_640), .Y (n_3557));
MX2X1 g64447(.A (n_11113), .B (n_3185), .S0 (n_10005), .Y (n_3555));
NOR2X1 g61315(.A (g_6701), .B (n_6705), .Y (n_4134));
MX2X1 g64461(.A (n_3388), .B (n_3178), .S0 (n_9333), .Y (n_3554));
NAND2X1 g64527(.A (n_3368), .B (n_3216), .Y (n_3552));
NAND3X1 g64567(.A (n_3569), .B (n_3550), .C (n_9466), .Y (n_3551));
XOR2X1 g64077(.A (n_523), .B (n_3547), .Y (n_3549));
NOR2X1 g64599(.A (g4581), .B (n_10376), .Y (n_6005));
NAND2X1 g64602(.A (n_3182), .B (n_3349), .Y (n_3546));
NAND3X1 g64658(.A (n_10940), .B (g3263), .C (n_10941), .Y (n_3543));
NAND3X1 g64683(.A (n_3398), .B (g3614), .C (n_6973), .Y (n_3542));
NAND4X1 g64739(.A (g3554), .B (n_10889), .C (g16656), .D (n_11128),.Y (n_3541));
NAND4X1 g64761(.A (n_1578), .B (n_3073), .C (n_9398), .D (n_477), .Y(n_3540));
XOR2X1 g64789(.A (g4311), .B (n_10396), .Y (n_3538));
INVX1 g64811(.A (g4581), .Y (n_5711));
DFFSRX1 g4000_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16693), .Q (g14518), .QN ());
AOI21X1 g62847(.A0 (n_3651), .A1 (n_10226), .B0 (n_8694), .Y(n_3537));
AND2X1 g64881(.A (n_5402), .B (g16693), .Y (n_3732));
NAND2X1 g64969(.A (g16693), .B (g16659), .Y (n_3535));
OAI21X1 g64971(.A0 (n_1390), .A1 (n_9129), .B0 (n_3160), .Y (n_3534));
OAI21X1 g64973(.A0 (n_1373), .A1 (n_9193), .B0 (n_3154), .Y (n_3533));
OAI21X1 g64975(.A0 (n_1384), .A1 (n_10952), .B0 (n_3158), .Y(n_3532));
OAI21X1 g64977(.A0 (n_1380), .A1 (n_9193), .B0 (n_3157), .Y (n_3531));
OAI21X1 g64978(.A0 (n_1366), .A1 (n_9628), .B0 (n_3156), .Y (n_3530));
OAI22X1 g62931(.A0 (n_3506), .A1 (n_2587), .B0 (n_1274), .B1(n_9651), .Y (n_3529));
INVX1 g65118(.A (g_5156), .Y (g8398));
INVX1 g65120(.A (g_6579), .Y (g8277));
DFFSRX1 g5798_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3120), .Q (), .QN (g_7062));
INVX1 g65124(.A (g_5508), .Y (g9615));
INVX1 g65126(.A (g_14965), .Y (g9741));
INVX1 g65128(.A (g_3861), .Y (g9817));
DFFSRX1 g3447_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3112), .Q (), .QN (g_5313));
NAND3X1 g61130(.A (n_3124), .B (g1389), .C (n_9811), .Y (n_3523));
DFFSRX1 g5456_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9555), .Q (), .QN (g5456));
DFFSRX1 g869_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14189), .Q (g14201), .QN ());
NAND2X1 g65326(.A (g_13255), .B (g_13901), .Y (n_3522));
DFFSRX1 g4489_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3116), .Q (g4489), .QN ());
OAI21X1 g64071(.A0 (n_10751), .A1 (g_15287), .B0 (n_3033), .Y(n_3521));
OAI22X1 g61962(.A0 (n_3489), .A1 (n_2161), .B0 (n_143), .B1 (n_9862),.Y (n_3520));
DFFSRX1 g1152_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3018), .Q (n_2429), .QN ());
INVX1 g65561(.A (g_11037), .Y (g9497));
INVX1 g65574(.A (g2724), .Y (n_3868));
INVX1 g65585(.A (g4145), .Y (n_3896));
NAND2X1 g65701(.A (n_1353), .B (n_3072), .Y (n_3518));
OR2X1 g65716(.A (g2715), .B (n_8898), .Y (n_3697));
XOR2X1 g64070(.A (g_13278), .B (n_3291), .Y (n_3517));
NAND2X1 g65868(.A (g2715), .B (n_8895), .Y (n_3695));
NAND3X1 g63243(.A (n_10005), .B (n_2757), .C (n_10647), .Y (n_3516));
DFFSRX1 g5105_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3122), .Q (g9553), .QN ());
DFFSRX1 g460_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3052), .Q (g_6131), .QN ());
AOI21X1 g63269(.A0 (n_3563), .A1 (n_741), .B0 (n_10296), .Y (n_3514));
OAI21X1 g63280(.A0 (n_7383), .A1 (n_9333), .B0 (n_3066), .Y (n_3512));
OAI21X1 g63282(.A0 (n_10889), .A1 (n_9797), .B0 (n_3063), .Y(n_3511));
MX2X1 g64100(.A (g4771), .B (n_2959), .S0 (n_9000), .Y (n_3510));
NAND3X1 g62103(.A (n_2800), .B (n_2697), .C (n_2764), .Y (n_3508));
OAI22X1 g62114(.A0 (n_3506), .A1 (n_2926), .B0 (n_165), .B1 (n_9992),.Y (n_3507));
NOR2X1 g63426(.A (n_8835), .B (n_8768), .Y (n_3505));
OAI21X1 g63440(.A0 (n_3502), .A1 (n_3501), .B0 (n_9279), .Y (n_3503));
OR2X1 g63474(.A (n_3499), .B (n_3497), .Y (n_3500));
NOR2X1 g63477(.A (n_2677), .B (n_3497), .Y (n_3498));
DFFSRX1 g4239_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3077), .Q (g4239), .QN ());
AOI21X1 g63484(.A0 (n_2751), .A1 (n_2744), .B0 (n_9976), .Y (n_3496));
NOR2X1 g63509(.A (n_8835), .B (n_8837), .Y (n_3855));
AOI21X1 g63526(.A0 (n_1783), .A1 (n_3493), .B0 (n_9836), .Y (n_3494));
AOI21X1 g63527(.A0 (n_7260), .A1 (g4349), .B0 (n_3491), .Y (n_3492));
OAI22X1 g63538(.A0 (n_3489), .A1 (n_1308), .B0 (g4688), .B1 (n_9830),.Y (n_3490));
AOI22X1 g63551(.A0 (n_2519), .A1 (n_10115), .B0 (g_12433), .B1(n_9693), .Y (n_3488));
DFFSRX1 g182_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3055), .Q (g_22379), .QN ());
DFFSRX1 g452_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3053), .Q (g_19241), .QN ());
DFFSRX1 g546_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3138), .Q (g_14587), .QN ());
OAI21X1 g63623(.A0 (n_3486), .A1 (n_3894), .B0 (n_2239), .Y (n_3487));
DFFSRX1 g4492_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3114), .Q (g4492), .QN ());
DFFSRX1 g4153_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3136), .Q (g4153), .QN ());
DFFSRX1 g168_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3057), .Q (g_20837), .QN ());
DFFSRX1 g3869_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3141), .Q (n_1191), .QN ());
DFFSRX1 g2984_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3139), .Q (g2984), .QN ());
INVX1 g61035(.A (n_6735), .Y (n_3484));
OAI22X1 g61222(.A0 (n_2672), .A1 (n_2562), .B0 (n_26), .B1 (n_9651),.Y (n_3483));
DFFSRX1 g538_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3133), .Q (g_21651), .QN ());
INVX1 g63926(.A (n_6767), .Y (n_3482));
NAND2X1 g63936(.A (g4072), .B (n_9952), .Y (n_3481));
NAND2X1 g63937(.A (g4072), .B (n_43), .Y (n_3480));
NAND2X1 g63947(.A (g4072), .B (n_98), .Y (n_3479));
NAND3X1 g63951(.A (n_3028), .B (n_83), .C (g_14265), .Y (n_3639));
DFFSRX1 g4273_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3131), .Q (g4273), .QN ());
OAI33X1 g63962(.A0 (n_1137), .A1 (n_2642), .A2 (n_546), .B0(n_10180), .B1 (n_1100), .B2 (n_75), .Y (n_3478));
INVX1 g63996(.A (n_3477), .Y (n_3845));
NAND2X2 g61049(.A (n_1444), .B (n_10330), .Y (n_3860));
DFFSRX1 g1339_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3167), .Q (), .QN (g1339));
DFFSRX1 g6167_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3010), .Q (g6167), .QN ());
OAI22X1 g64024(.A0 (n_3506), .A1 (n_1827), .B0 (g4878), .B1(n_10063), .Y (n_3475));
DFFSRX1 g86_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3143), .Q (g20557), .QN ());
NAND4X1 g64059(.A (n_2378), .B (n_2965), .C (n_2025), .D (n_2027), .Y(n_11188));
DFFSRX1 g174_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3056), .Q (g_21806), .QN ());
DFFSRX1 g5495_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3012), .Q (), .QN (g5495));
DFFSRX1 g6533_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3008), .Q (), .QN (g6533));
DFFSRX1 g962_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3005), .Q (g_15758), .QN ());
DFFSRX1 g4643_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3212), .Q (n_276), .QN ());
DFFSRX1 g5176_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3147), .Q (n_1177), .QN ());
DFFSRX1 g5523_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3146), .Q (n_1234), .QN ());
DFFSRX1 g5869_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3140), .Q (n_1169), .QN ());
DFFSRX1 g6561_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3144), .Q (n_1216), .QN ());
DFFSRX1 g3167_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3145), .Q (n_1135), .QN ());
DFFSRX1 g3518_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3142), .Q (n_1210), .QN ());
DFFSRX1 g215_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3137), .Q (g8291), .QN ());
DFFSRX1 g4172_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3132), .Q (g4172), .QN ());
DFFSRX1 g4486_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3119), .Q (g4486), .QN ());
DFFSRX1 g2912_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3105), .Q (g2912), .QN ());
DFFSRX1 g2868_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3096), .Q (g2868), .QN ());
DFFSRX1 g2936_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3090), .Q (g2936), .QN ());
DFFSRX1 g1779_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3097), .Q (g1779), .QN ());
DFFSRX1 g1798_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3111), .Q (g1798), .QN ());
DFFSRX1 g1913_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3106), .Q (g1913), .QN ());
DFFSRX1 g1932_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3080), .Q (g1932), .QN ());
DFFSRX1 g136_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3102), .Q (g21292), .QN ());
DFFSRX1 g365_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3127), .Q (g8719), .QN ());
DFFSRX1 g2047_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3099), .Q (g2047), .QN ());
DFFSRX1 g2066_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3098), .Q (g2066), .QN ());
DFFSRX1 g4146_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3095), .Q (g4146), .QN ());
DFFSRX1 g2204_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3103), .Q (g2204), .QN ());
DFFSRX1 g2223_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3108), .Q (g2223), .QN ());
DFFSRX1 g4249_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3094), .Q (g4249), .QN ());
DFFSRX1 g2922_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3081), .Q (g2922), .QN ());
DFFSRX1 g2338_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3091), .Q (g2338), .QN ());
DFFSRX1 g2357_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3085), .Q (g2357), .QN ());
DFFSRX1 g4639_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3130), .Q (n_7247), .QN ());
DFFSRX1 g4717_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3088), .Q (g4717), .QN ());
DFFSRX1 g1664_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3086), .Q (g1664), .QN ());
DFFSRX1 g2472_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3084), .Q (g2472), .QN ());
DFFSRX1 g2491_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3082), .Q (g2491), .QN ());
DFFSRX1 g4907_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3092), .Q (g4907), .QN ());
DFFSRX1 g2606_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3079), .Q (g2606), .QN ());
DFFSRX1 g1644_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3109), .Q (g1644), .QN ());
DFFSRX1 g2625_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3100), .Q (g2625), .QN ());
DFFSRX1 g2994_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3104), .Q (g2994), .QN ());
DFFSRX1 g1291_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3070), .Q (g1291), .QN ());
MX2X1 g64095(.A (g20652), .B (n_2678), .S0 (n_8955), .Y (n_3473));
MX2X1 g64097(.A (g4704), .B (n_2961), .S0 (n_9234), .Y (n_3471));
MX2X1 g64098(.A (g4749), .B (n_2962), .S0 (n_8955), .Y (n_3470));
MX2X1 g64099(.A (g4760), .B (n_2960), .S0 (n_9000), .Y (n_3469));
MX2X1 g64102(.A (g4939), .B (n_2963), .S0 (n_9000), .Y (n_3468));
MX2X1 g64103(.A (g4950), .B (n_2958), .S0 (n_9156), .Y (n_3466));
MX2X1 g64104(.A (g4961), .B (n_2957), .S0 (n_9311), .Y (n_3465));
OAI21X1 g64136(.A0 (n_2942), .A1 (n_3463), .B0 (n_9091), .Y (n_3464));
NAND3X1 g64179(.A (n_2989), .B (n_2243), .C (n_2632), .Y (n_3461));
OAI33X1 g61062(.A0 (n_2841), .A1 (n_3365), .A2 (n_3459), .B0(n_11073), .B1 (n_3459), .B2 (n_10245), .Y (n_3460));
NAND3X1 g61721(.A (n_2979), .B (n_2245), .C (n_2870), .Y (n_3458));
INVX2 g64232(.A (n_3814), .Y (n_3455));
NAND3X1 g61723(.A (n_3222), .B (n_2557), .C (n_2350), .Y (n_3454));
NAND3X1 g64244(.A (n_10398), .B (g4616), .C (g4584), .Y (n_4843));
AOI21X1 g64290(.A0 (n_2641), .A1 (n_2934), .B0 (n_3391), .Y (n_3449));
NAND2X1 g62581(.A (n_3447), .B (g_15381), .Y (n_3448));
NAND4X1 g64307(.A (n_3030), .B (n_1262), .C (n_3021), .D (n_2456), .Y(n_3442));
AOI21X1 g64316(.A0 (n_2983), .A1 (n_10867), .B0 (n_3832), .Y(n_3831));
AOI21X1 g64319(.A0 (n_3569), .A1 (g_14265), .B0 (n_3174), .Y(n_3441));
AOI21X1 g64324(.A0 (n_2670), .A1 (n_10871), .B0 (n_3838), .Y(n_3837));
AOI21X1 g64340(.A0 (n_11033), .A1 (n_10867), .B0 (n_8629), .Y(n_3873));
AOI21X1 g64342(.A0 (n_11036), .A1 (n_10867), .B0 (n_8634), .Y(n_3870));
OAI21X1 g64352(.A0 (n_3425), .A1 (n_3439), .B0 (n_3438), .Y (n_3440));
AOI21X1 g64356(.A0 (g14662), .A1 (n_465), .B0 (n_3228), .Y (n_3437));
AOI21X1 g64357(.A0 (g14694), .A1 (n_409), .B0 (n_3229), .Y (n_3436));
AOI21X1 g64358(.A0 (g14738), .A1 (n_11045), .B0 (n_3226), .Y(n_3435));
AOI21X1 g64359(.A0 (g14779), .A1 (n_660), .B0 (n_3225), .Y (n_3434));
AOI21X1 g64360(.A0 (g14828), .A1 (n_322), .B0 (n_3223), .Y (n_3433));
OR2X1 g64367(.A (n_3004), .B (n_3431), .Y (n_3432));
XOR2X1 g64374(.A (n_3894), .B (n_3486), .Y (n_3430));
OAI22X1 g64375(.A0 (n_1568), .A1 (n_3569), .B0 (n_3003), .B1 (n_708),.Y (n_3429));
AOI21X1 g64404(.A0 (g5033), .A1 (n_9193), .B0 (n_3233), .Y (n_3427));
DFFSRX1 g1589_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3179), .Q (g1589), .QN ());
XOR2X1 g64410(.A (n_659), .B (n_3425), .Y (n_3426));
MX2X1 g64415(.A (g_19233), .B (g_17065), .S0 (n_3003), .Y (n_3424));
MX2X1 g64416(.A (n_11162), .B (n_3550), .S0 (n_3003), .Y (n_3423));
MX2X1 g64418(.A (g_21778), .B (g_19113), .S0 (n_3003), .Y (n_3422));
MX2X1 g64419(.A (g_17065), .B (g_16677), .S0 (n_3003), .Y (n_3420));
MX2X1 g64420(.A (g_16677), .B (g_20208), .S0 (n_3003), .Y (n_3418));
MX2X1 g64421(.A (g_21720), .B (g_13758), .S0 (n_3003), .Y (n_3417));
MX2X1 g64422(.A (g_13758), .B (g_19289), .S0 (n_3003), .Y (n_3416));
MX2X1 g64423(.A (g_19289), .B (n_5663), .S0 (n_3003), .Y (n_3415));
OAI21X1 g62667(.A0 (n_221), .A1 (n_9311), .B0 (n_3193), .Y (n_3414));
MX2X1 g64442(.A (g_17426), .B (n_2891), .S0 (n_9172), .Y (n_3413));
OAI22X1 g62679(.A0 (n_3489), .A1 (n_1989), .B0 (n_294), .B1 (n_9862),.Y (n_3412));
INVX1 g64472(.A (g5069), .Y (n_3411));
INVX1 g64488(.A (g2946), .Y (n_3410));
DFFSRX1 g203_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3176), .Q (), .QN (g_7563));
DFFSRX1 g3317_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14421), .Q (g16874), .QN ());
DFFSRX1 g3668_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14451), .Q (g16924), .QN ());
NOR2X1 g64522(.A (n_3208), .B (n_653), .Y (n_3409));
DFFSRX1 g4722_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_3087), .Q (g4722), .QN ());
OAI21X1 g64531(.A0 (n_2372), .A1 (n_887), .B0 (n_3194), .Y (n_3408));
AOI21X1 g61327(.A0 (n_2060), .A1 (n_26), .B0 (n_3186), .Y (n_3407));
OAI21X1 g64534(.A0 (n_2370), .A1 (n_882), .B0 (n_3207), .Y (n_3406));
OAI21X1 g64544(.A0 (n_2615), .A1 (n_880), .B0 (n_3204), .Y (n_3404));
OAI21X1 g64546(.A0 (n_2366), .A1 (n_888), .B0 (n_3202), .Y (n_3403));
OAI21X1 g64549(.A0 (n_2368), .A1 (n_977), .B0 (n_3201), .Y (n_3402));
OAI21X1 g64566(.A0 (n_2367), .A1 (n_838), .B0 (n_3200), .Y (n_3400));
INVX1 g64571(.A (n_8707), .Y (n_3399));
AND2X1 g64600(.A (n_3398), .B (n_6972), .Y (n_3758));
OAI21X1 g64613(.A0 (n_2365), .A1 (n_881), .B0 (n_3206), .Y (n_3395));
INVX1 g64620(.A (n_3784), .Y (n_3394));
INVX2 g64641(.A (n_3547), .Y (n_3605));
DFFSRX1 g6159_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2712), .Q (g6159), .QN ());
NAND2X1 g64660(.A (n_3425), .B (n_3391), .Y (n_3822));
DFFSRX1 g3155_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2854), .Q (g3155), .QN ());
AOI21X1 g64682(.A0 (n_1090), .A1 (n_1279), .B0 (n_3569), .Y (n_3390));
AOI21X1 g64689(.A0 (n_3177), .A1 (n_3388), .B0 (n_2628), .Y (n_3389));
NAND4X1 g64690(.A (n_1656), .B (n_3984), .C (n_10005), .D (g5029), .Y(n_3387));
NAND4X1 g64048(.A (n_2977), .B (n_2389), .C (n_2344), .D (n_2340), .Y(n_3385));
AOI22X1 g64703(.A0 (n_2610), .A1 (n_3383), .B0 (g1472), .B1 (n_9628),.Y (n_3384));
MX2X1 g64707(.A (n_1629), .B (n_2595), .S0 (n_4617), .Y (n_3382));
AOI22X1 g64787(.A0 (n_2361), .A1 (n_598), .B0 (n_3073), .B1 (n_653),.Y (n_3381));
DFFSRX1 g4581_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2863), .Q (), .QN (g4581));
OAI21X1 g64843(.A0 (n_2575), .A1 (g2975), .B0 (n_9351), .Y (n_3377));
NAND2X1 g64918(.A (n_2880), .B (n_6406), .Y (n_3376));
NAND3X1 g61120(.A (n_3372), .B (n_2), .C (n_11041), .Y (n_3373));
AOI21X1 g65001(.A0 (g16775), .A1 (n_493), .B0 (n_2869), .Y (n_3371));
DFFSRX1 g976_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2846), .Q (g_6701), .QN ());
DFFSRX1 g5170_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2914), .Q (g5170), .QN ());
AOI22X1 g65018(.A0 (n_2215), .A1 (n_3177), .B0 (g_22021), .B1(n_9193), .Y (n_3370));
DFFSRX1 g5527_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2903), .Q (g5527), .QN ());
NAND3X1 g61122(.A (n_3123), .B (n_3364), .C (n_9664), .Y (n_3369));
AOI22X1 g65034(.A0 (n_2496), .A1 (n_3177), .B0 (g_18996), .B1(n_9599), .Y (n_3368));
DFFSRX1 g3119_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2709), .Q (g3119), .QN ());
DFFSRX1 g5128_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2720), .Q (g5128), .QN ());
DFFSRX1 g5857_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2858), .Q (g5857), .QN ());
DFFSRX1 g3798_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2829), .Q (), .QN (g_5156));
DFFSRX1 g3096_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2831), .Q (), .QN (g_6579));
DFFSRX1 g5452_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2839), .Q (), .QN (g_5508));
DFFSRX1 g6144_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2833), .Q (), .QN (g_14965));
DFFSRX1 g6490_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2837), .Q (), .QN (g_3861));
DFFSRX1 g3841_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2693), .Q (), .QN (g3841));
AOI21X1 g61132(.A0 (n_3365), .A1 (n_3364), .B0 (n_2834), .Y (n_3366));
DFFSRX1 g5517_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2913), .Q (g5517), .QN ());
DFFSRX1 g4462_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2955), .Q (g4462), .QN ());
DFFSRX1 g4264_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2949), .Q (g4264), .QN ());
DFFSRX1 g2704_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2827), .Q (g2704), .QN ());
DFFSRX1 g5092_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2954), .Q (g5092), .QN ());
DFFSRX1 g1548_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2947), .Q (g1548), .QN ());
DFFSRX1 g3490_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2700), .Q (), .QN (g3490));
AOI22X1 g61955(.A0 (n_2495), .A1 (n_2878), .B0 (g_20563), .B1(n_9129), .Y (n_3363));
AOI22X1 g65441(.A0 (n_2506), .A1 (n_1751), .B0 (g3522), .B1 (n_9129),.Y (n_3362));
AOI22X1 g65442(.A0 (n_2494), .A1 (n_1718), .B0 (g6565), .B1 (n_9491),.Y (n_3361));
AOI22X1 g65444(.A0 (n_2500), .A1 (n_1777), .B0 (g5527), .B1 (n_9129),.Y (n_3360));
OAI22X1 g65499(.A0 (n_2559), .A1 (g4297), .B0 (n_150), .B1 (n_9992),.Y (n_3359));
OAI21X1 g65529(.A0 (n_32), .A1 (n_9681), .B0 (n_2840), .Y (n_3358));
INVX1 g65534(.A (g2927), .Y (n_3357));
DFFSRX1 g2878_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2775), .Q (), .QN (g2878));
DFFSRX1 g5794_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2766), .Q (g9617), .QN ());
DFFSRX1 g3092_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2776), .Q (g8215), .QN ());
DFFSRX1 g6140_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2765), .Q (g9682), .QN ());
DFFSRX1 g3443_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2769), .Q (g8279), .QN ());
DFFSRX1 g6486_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2772), .Q (g9743), .QN ());
INVX1 g65551(.A (g_13901), .Y (n_3519));
DFFSRX1 g5101_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2777), .Q (), .QN (g_11037));
DFFSRX1 g3794_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2770), .Q (g8344), .QN ());
INVX1 g65567(.A (g2965), .Y (n_3356));
DFFSRX1 g2724_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2796), .Q (g2724), .QN ());
DFFSRX1 g3003_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2789), .Q (), .QN (g3003));
DFFSRX1 g4145_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2788), .Q (g4145), .QN ());
DFFSRX1 g4164_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2793), .Q (), .QN (g4164));
DFFSRX1 g1521_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2774), .Q (g1521), .QN ());
DFFSRX1 g1099_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2725), .Q (g_19172), .QN ());
DFFSRX1 g6187_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2705), .Q (), .QN (g6187));
MX2X1 g63135(.A (n_7260), .B (n_2484), .S0 (n_9501), .Y (n_3355));
DFFSRX1 g3139_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2687), .Q (), .QN (g3139));
DFFSRX1 g1442_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2690), .Q (g1442), .QN ());
DFFSRX1 g5467_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2716), .Q (g5467), .QN ());
DFFSRX1 g3462_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2703), .Q (g3462), .QN ());
NAND2X1 g65986(.A (n_3071), .B (n_2862), .Y (n_3353));
DFFSRX1 g4269_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2759), .Q (g4269), .QN ());
NOR2X1 g63226(.A (n_2580), .B (n_3651), .Y (n_3352));
AND2X1 g63231(.A (n_3651), .B (n_3332), .Y (n_3351));
NAND2X1 g63232(.A (n_3651), .B (n_3707), .Y (n_3350));
NAND2X1 g63233(.A (n_3651), .B (n_9493), .Y (n_3720));
DFFSRX1 g4093_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2787), .Q (g4093), .QN ());
NAND4X1 g66084(.A (n_3181), .B (n_7247), .C (n_9940), .D (n_23), .Y(n_3349));
MX2X1 g61169(.A (g1521), .B (n_2475), .S0 (n_8955), .Y (n_3348));
DFFSRX1 g6505_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2707), .Q (g6505), .QN ());
DFFSRX1 g6215_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2864), .Q (n_1214), .QN ());
DFFSRX1 g37_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2819), .Q (), .QN (g23002));
AOI21X1 g61480(.A0 (n_2192), .A1 (n_129), .B0 (n_2791), .Y (n_3347));
INVX1 g66272(.A (g2715), .Y (n_3679));
XOR2X1 g63329(.A (n_2754), .B (n_8913), .Y (n_3346));
NAND2X1 g61494(.A (n_2488), .B (n_3316), .Y (n_3345));
NOR2X1 g66362(.A (n_11), .B (n_9359), .Y (n_3344));
NOR2X1 g66369(.A (n_5363), .B (n_9453), .Y (n_3343));
DFFSRX1 g5148_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2719), .Q (), .QN (g5148));
DFFSRX1 g4340_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2753), .Q (n_7260), .QN ());
NOR2X1 g66409(.A (n_596), .B (n_9398), .Y (n_3341));
NOR2X1 g66471(.A (n_571), .B (n_9453), .Y (n_3340));
NOR2X1 g66512(.A (n_118), .B (n_9398), .Y (n_3339));
DFFSRX1 g3522_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2894), .Q (g3522), .QN ());
NOR2X1 g66528(.A (n_572), .B (n_9940), .Y (n_3337));
NOR2X1 g66558(.A (n_504), .B (n_9940), .Y (n_3336));
OR2X1 g66644(.A (g2759), .B (n_9359), .Y (n_3335));
INVX1 g63453(.A (n_3447), .Y (n_3334));
NAND2X1 g63455(.A (n_3332), .B (n_8913), .Y (n_3333));
NOR2X1 g63457(.A (n_3563), .B (n_9903), .Y (n_3331));
NAND3X1 g63475(.A (n_3149), .B (n_3148), .C (g2882), .Y (n_3330));
DFFSRX1 g2145_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2814), .Q (g2145), .QN ());
AND2X1 g63513(.A (n_3563), .B (n_2465), .Y (n_3329));
NAND2X1 g63514(.A (n_3563), .B (n_11134), .Y (n_3328));
NAND2X1 g63515(.A (n_3563), .B (n_9553), .Y (n_3687));
NAND4X1 g63519(.A (n_2945), .B (n_1331), .C (n_10119), .D (n_2303),.Y (n_3327));
NAND4X1 g63531(.A (n_2660), .B (n_2209), .C (n_2135), .D (n_1701), .Y(n_3326));
NAND4X1 g63534(.A (n_2986), .B (n_2408), .C (n_2122), .D (n_1698), .Y(n_3325));
AOI21X1 g63540(.A0 (n_2468), .A1 (n_2451), .B0 (n_3323), .Y (n_3324));
OAI22X1 g64064(.A0 (n_2624), .A1 (n_9599), .B0 (n_2645), .B1(n_9811), .Y (n_3322));
AOI22X1 g63554(.A0 (n_2263), .A1 (n_8840), .B0 (g1189), .B1 (n_9193),.Y (n_3321));
OAI21X1 g64043(.A0 (n_719), .A1 (n_9311), .B0 (n_2740), .Y (n_3320));
OAI21X1 g64030(.A0 (n_2734), .A1 (n_9681), .B0 (n_2735), .Y (n_3319));
OAI21X1 g61550(.A0 (n_92), .A1 (n_9978), .B0 (n_3316), .Y (n_3317));
OAI22X1 g64063(.A0 (n_2398), .A1 (n_9269), .B0 (n_2647), .B1(n_9811), .Y (n_3315));
DFFSRX1 g1319_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2739), .Q (g1319), .QN ());
DFFSRX1 g2860_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2822), .Q (g2860), .QN ());
XOR2X1 g63646(.A (n_10188), .B (n_2723), .Y (n_3314));
OAI22X1 g64068(.A0 (n_2392), .A1 (n_9836), .B0 (n_2646), .B1(n_9811), .Y (n_3313));
NAND3X1 g61034(.A (n_6734), .B (n_1043), .C (n_9425), .Y (n_3312));
DFFSRX1 g1205_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2953), .Q (n_10129), .QN ());
DFFSRX1 g4912_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2804), .Q (g4912), .QN ());
DFFSRX1 g4927_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2802), .Q (g4927), .QN ());
DFFSRX1 g2907_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2805), .Q (g2907), .QN ());
DFFSRX1 g5164_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2860), .Q (g5164), .QN ());
NOR2X1 g63866(.A (n_10532), .B (n_3310), .Y (n_3915));
AND2X1 g63867(.A (n_10115), .B (n_3310), .Y (n_3309));
NAND2X1 g61644(.A (n_2879), .B (n_2742), .Y (n_3308));
NAND2X1 g63902(.A (n_2465), .B (n_10188), .Y (n_3307));
NAND3X1 g63918(.A (n_6766), .B (n_1541), .C (n_9940), .Y (n_3305));
NOR2X1 g63934(.A (n_2749), .B (n_957), .Y (n_3303));
AOI21X1 g63969(.A0 (n_1789), .A1 (n_3031), .B0 (n_2741), .Y (n_3302));
DFFSRX1 g862_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2896), .Q (g_22552), .QN ());
OAI22X1 g64067(.A0 (n_2397), .A1 (n_9193), .B0 (n_2642), .B1(n_9311), .Y (n_3301));
INVX1 g63997(.A (n_8835), .Y (n_3477));
DFFSRX1 g2873_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2816), .Q (g2873), .QN ());
DFFSRX1 g4427_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2801), .Q (g4427), .QN ());
OAI21X1 g64025(.A0 (n_1695), .A1 (n_9425), .B0 (n_2736), .Y (n_3300));
OAI21X1 g64027(.A0 (n_2421), .A1 (n_9940), .B0 (n_2733), .Y (n_3299));
OAI21X1 g64028(.A0 (n_11150), .A1 (n_9422), .B0 (n_2730), .Y(n_3298));
OAI21X1 g64029(.A0 (n_11173), .A1 (n_9333), .B0 (n_2727), .Y(n_3296));
DFFSRX1 g1189_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2886), .Q (g1189), .QN ());
DFFSRX1 g3821_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2694), .Q (g3821), .QN ());
DFFSRX1 g5097_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2761), .Q (g5097), .QN ());
DFFSRX1 g1221_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2760), .Q (g1221), .QN ());
DFFSRX1 g1564_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2758), .Q (g1564), .QN ());
DFFSRX1 g5120_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2722), .Q (g5120), .QN ());
DFFSRX1 g5475_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2715), .Q (g5475), .QN ());
DFFSRX1 g5821_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2713), .Q (g5821), .QN ());
DFFSRX1 g5813_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2714), .Q (g5813), .QN ());
DFFSRX1 g6513_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2706), .Q (g6513), .QN ());
DFFSRX1 g3813_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2695), .Q (g3813), .QN ());
DFFSRX1 g209_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2691), .Q (g_18635), .QN ());
DFFSRX1 g4277_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2689), .Q (g8839), .QN ());
DFFSRX1 g1495_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2688), .Q (n_2005), .QN ());
DFFSRX1 g4304_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2682), .Q (g9251), .QN ());
DFFSRX1 g376_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2951), .Q (g_20952), .QN ());
DFFSRX1 g5180_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2904), .Q (g5180), .QN ());
DFFSRX1 g5863_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2906), .Q (g5863), .QN ());
DFFSRX1 g3171_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2897), .Q (g3171), .QN ());
DFFSRX1 g6219_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2898), .Q (g6219), .QN ());
DFFSRX1 g6565_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2888), .Q (g6565), .QN ());
DFFSRX1 g3512_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2910), .Q (g3512), .QN ());
DFFSRX1 g3863_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2907), .Q (g3863), .QN ());
DFFSRX1 g3873_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2892), .Q (g3873), .QN ());
DFFSRX1 g3161_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2909), .Q (g3161), .QN ());
DFFSRX1 g1532_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2889), .Q (g1532), .QN ());
DFFSRX1 g1178_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2887), .Q (g1178), .QN ());
DFFSRX1 g6555_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2911), .Q (g6555), .QN ());
OAI22X1 g64082(.A0 (n_2625), .A1 (n_10078), .B0 (n_2644), .B1(n_10063), .Y (n_3292));
DFFSRX1 g2844_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2821), .Q (g2844), .QN ());
DFFSRX1 g2852_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2826), .Q (g2852), .QN ());
DFFSRX1 g5511_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2856), .Q (g5511), .QN ());
DFFSRX1 g2894_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2820), .Q (g2894), .QN ());
DFFSRX1 g2950_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2824), .Q (g2950), .QN ());
DFFSRX1 g6549_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2843), .Q (g6549), .QN ());
DFFSRX1 g94_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2810), .Q (g20652), .QN ());
DFFSRX1 g3506_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2850), .Q (g3506), .QN ());
DFFSRX1 g2697_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2807), .Q (g2697), .QN ());
DFFSRX1 g2988_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2762), .Q (g2988), .QN ());
DFFSRX1 g3857_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2848), .Q (g3857), .QN ());
DFFSRX1 g2138_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2815), .Q (g2138), .QN ());
DFFSRX1 g4157_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2832), .Q (g4157), .QN ());
DFFSRX1 g4245_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2813), .Q (g4245), .QN ());
DFFSRX1 g4253_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2812), .Q (g4253), .QN ());
DFFSRX1 g2970_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2808), .Q (g2970), .QN ());
DFFSRX1 g2960_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2817), .Q (g2960), .QN ());
DFFSRX1 g4732_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2806), .Q (g4732), .QN ());
DFFSRX1 g4737_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2823), .Q (g4737), .QN ());
DFFSRX1 g4922_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2803), .Q (g4922), .QN ());
DFFSRX1 g4098_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2767), .Q (g4098), .QN ());
DFFSRX1 g947_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2768), .Q (g_22349), .QN ());
DFFSRX1 g4258_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2782), .Q (g4258), .QN ());
DFFSRX1 g4537_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2956), .Q (g10306), .QN ());
NAND2X1 g64149(.A (n_3291), .B (g_13278), .Y (n_3690));
OAI21X1 g64153(.A0 (n_2616), .A1 (n_890), .B0 (n_2974), .Y (n_3290));
NOR2X1 g64155(.A (n_2675), .B (n_6694), .Y (n_3289));
OAI21X1 g61061(.A0 (n_2938), .A1 (n_3183), .B0 (n_10005), .Y(n_3288));
AND2X1 g64158(.A (n_2663), .B (n_3025), .Y (n_3287));
NAND4X1 g64166(.A (g5220), .B (n_10621), .C (n_1695), .D (g5339), .Y(n_3286));
DFFSRX1 g2980_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2915), .Q (g2980), .QN ());
NAND4X1 g64181(.A (n_2673), .B (n_512), .C (n_448), .D (n_262), .Y(n_3285));
NAND2X2 g64233(.A (n_3236), .B (n_2039), .Y (n_3814));
NAND3X1 g64235(.A (n_2666), .B (n_2486), .C (n_2400), .Y (n_3283));
NAND3X1 g64236(.A (n_2665), .B (n_2536), .C (n_2634), .Y (n_3282));
NAND4X1 g64256(.A (g5567), .B (n_7150), .C (n_2208), .D (g5685), .Y(n_3281));
NAND3X1 g61726(.A (n_2972), .B (n_2530), .C (n_2603), .Y (n_3279));
NAND4X1 g64257(.A (g6259), .B (n_3277), .C (n_11150), .D (g6377), .Y(n_3278));
NAND4X1 g64275(.A (g6605), .B (n_3275), .C (n_11173), .D (g6723), .Y(n_3276));
AND2X1 g64278(.A (n_10693), .B (n_2077), .Y (n_3829));
NOR2X1 g64315(.A (n_2664), .B (n_2866), .Y (n_3274));
NAND3X1 g64039(.A (n_2658), .B (n_2548), .C (n_2459), .Y (n_3273));
AOI21X1 g64361(.A0 (n_2679), .A1 (n_10134), .B0 (n_2680), .Y(n_3271));
OAI21X1 g64365(.A0 (n_23), .A1 (n_9422), .B0 (n_2981), .Y (n_3270));
NAND4X1 g64376(.A (n_10831), .B (g5204), .C (g25219), .D (g5339), .Y(n_3269));
NAND4X1 g64382(.A (n_2439), .B (g5551), .C (n_1023), .D (g5685), .Y(n_3268));
NAND4X1 g64383(.A (n_2413), .B (g6243), .C (n_11157), .D (g6377), .Y(n_3267));
NAND4X1 g64384(.A (n_10809), .B (g5897), .C (n_546), .D (g6031), .Y(n_3266));
NAND4X1 g64385(.A (n_2435), .B (g6589), .C (n_11177), .D (g6723), .Y(n_3265));
NAND4X1 g64387(.A (n_2042), .B (n_3984), .C (g5041), .D (n_10771), .Y(n_3264));
OAI21X1 g62646(.A0 (n_307), .A1 (n_9333), .B0 (n_2946), .Y (n_3263));
DFFSRX1 g5841_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2685), .Q (), .QN (g5841));
NOR2X1 g62649(.A (n_2662), .B (g3343), .Y (n_3262));
NOR2X1 g62651(.A (n_2669), .B (g3694), .Y (n_3261));
XOR2X1 g64402(.A (n_2637), .B (n_3259), .Y (n_3260));
DFFSRX1 g5873_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2900), .Q (g5873), .QN ());
DFFSRX1 g3470_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2702), .Q (g3470), .QN ());
INVX1 g64411(.A (n_3258), .Y (n_3645));
AOI22X1 g64414(.A0 (n_2410), .A1 (n_8637), .B0 (n_3152), .B1 (n_644),.Y (n_3257));
OAI21X1 g62658(.A0 (n_1295), .A1 (n_9940), .B0 (n_2939), .Y (n_3255));
MX2X1 g64437(.A (n_3253), .B (n_1802), .S0 (n_9627), .Y (n_3254));
DFFSRX1 g5069_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2905), .Q (g5069), .QN ());
DFFSRX1 g2932_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2902), .Q (), .QN (g2932));
DFFSRX1 g4284_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2890), .Q (), .QN (g4284));
DFFSRX1 g2946_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2895), .Q (g2946), .QN ());
NOR2X1 g64509(.A (n_3569), .B (g_22639), .Y (n_3566));
INVX2 g64537(.A (n_3249), .Y (n_3775));
NAND3X1 g64551(.A (n_2654), .B (n_10664), .C (n_9717), .Y (n_3247));
DFFSRX1 g896_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2948), .Q (g_16404), .QN ());
INVX2 g64569(.A (g28753), .Y (n_3244));
NOR2X1 g64575(.A (n_3486), .B (n_2828), .Y (n_3243));
DFFSRX1 g6209_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2912), .Q (g6209), .QN ());
NAND2X1 g64579(.A (n_3569), .B (g_19113), .Y (n_3242));
NAND3X1 g64580(.A (n_835), .B (n_2609), .C (n_9558), .Y (n_3241));
INVX4 g64587(.A (n_3239), .Y (n_3779));
INVX1 g64634(.A (n_4053), .Y (n_4832));
CLKBUFX1 g64642(.A (n_3236), .Y (n_3547));
NAND2X1 g64645(.A (n_3224), .B (n_659), .Y (n_3234));
NOR3X1 g64648(.A (n_3016), .B (g5037), .C (n_9107), .Y (n_3233));
INVX1 g64650(.A (n_10461), .Y (n_3832));
NAND4X1 g64656(.A (n_1643), .B (n_1084), .C (n_9521), .D (n_2881), .Y(n_3229));
NAND4X1 g64657(.A (n_1642), .B (n_1085), .C (n_9501), .D (n_3171), .Y(n_3228));
NAND4X1 g64659(.A (n_1381), .B (n_842), .C (n_9139), .D (n_2732), .Y(n_3226));
NAND4X1 g64661(.A (n_1641), .B (n_1083), .C (n_9091), .D (n_2729), .Y(n_3225));
NAND2X1 g64686(.A (n_3224), .B (n_3391), .Y (n_3438));
NAND4X1 g64688(.A (n_1640), .B (n_1082), .C (n_9091), .D (n_2871), .Y(n_3223));
NAND3X1 g61809(.A (n_851), .B (n_1996), .C (n_10949), .Y (n_3222));
NAND3X1 g61812(.A (n_722), .B (n_1647), .C (n_10949), .Y (n_3221));
NAND4X1 g64731(.A (n_2447), .B (g3953), .C (g16659), .D (n_4988), .Y(n_3219));
NAND4X1 g64772(.A (n_7010), .B (n_1493), .C (g5033), .D (n_3984), .Y(n_3218));
MX2X1 g64781(.A (g4888), .B (g4894), .S0 (n_2351), .Y (n_3217));
DFFSRX1 g3298_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16624), .Q (g14421), .QN ());
DFFSRX1 g3649_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16656), .Q (g14451), .QN ());
NAND3X1 g64853(.A (n_2883), .B (g_18996), .C (n_9681), .Y (n_3216));
AND2X1 g64892(.A (n_10897), .B (g16656), .Y (n_3398));
NAND2X1 g64898(.A (n_10400), .B (g4311), .Y (n_3258));
NAND3X1 g64903(.A (n_2055), .B (n_3213), .C (n_276), .Y (n_3214));
AND2X1 g64912(.A (n_2614), .B (g4633), .Y (n_3212));
NOR2X1 g64924(.A (n_3641), .B (n_6400), .Y (n_3211));
NAND2X1 g64939(.A (g16624), .B (g16603), .Y (n_3210));
NAND2X1 g64941(.A (g16656), .B (g16627), .Y (n_3209));
NOR2X1 g64964(.A (n_2602), .B (n_10296), .Y (n_3208));
INVX1 g61116(.A (n_3910), .Y (n_4866));
AOI22X1 g64986(.A0 (n_2218), .A1 (n_4327), .B0 (n_1807), .B1(n_9193), .Y (n_3207));
AOI22X1 g64988(.A0 (n_2206), .A1 (n_4324), .B0 (n_2084), .B1(n_9599), .Y (n_3206));
AOI22X1 g64989(.A0 (n_2227), .A1 (n_4316), .B0 (n_1805), .B1(n_9193), .Y (n_3204));
AOI22X1 g64992(.A0 (n_2204), .A1 (n_4322), .B0 (n_1794), .B1(n_10376), .Y (n_3202));
AOI22X1 g64995(.A0 (n_2207), .A1 (n_4320), .B0 (n_1799), .B1(n_9526), .Y (n_3201));
AOI22X1 g64998(.A0 (n_2211), .A1 (n_4314), .B0 (n_1796), .B1(n_9193), .Y (n_3200));
AOI22X1 g65002(.A0 (n_2205), .A1 (n_1422), .B0 (g1442), .B1 (n_9300),.Y (n_3197));
AOI22X1 g65004(.A0 (n_2210), .A1 (n_2008), .B0 (g1478), .B1 (n_9672),.Y (n_3196));
AOI22X1 g65005(.A0 (n_2228), .A1 (n_4329), .B0 (n_1810), .B1(n_9193), .Y (n_3194));
MX2X1 g62926(.A (n_2305), .B (n_3192), .S0 (n_2166), .Y (n_3193));
AOI22X1 g65006(.A0 (n_2216), .A1 (n_1252), .B0 (g1448), .B1 (n_9300),.Y (n_3191));
AOI22X1 g65019(.A0 (n_2276), .A1 (n_1655), .B0 (n_10134), .B1(n_9129), .Y (n_3189));
NAND3X1 g61121(.A (g1384), .B (n_2830), .C (n_9558), .Y (n_3187));
NAND2X1 g61369(.A (n_2671), .B (n_2563), .Y (n_3186));
OAI21X1 g65052(.A0 (n_3184), .A1 (n_10524), .B0 (n_2611), .Y(n_3185));
AND2X1 g61123(.A (n_1503), .B (n_3183), .Y (n_3628));
AOI22X1 g65058(.A0 (n_2316), .A1 (n_3181), .B0 (n_7247), .B1(n_9491), .Y (n_3182));
OAI21X1 g61372(.A0 (g1585), .A1 (n_9797), .B0 (n_3165), .Y (n_3179));
AOI22X1 g65084(.A0 (n_1221), .A1 (n_2577), .B0 (n_3177), .B1(n_10528), .Y (n_3178));
MX2X1 g65107(.A (n_2017), .B (n_2320), .S0 (n_9000), .Y (n_3176));
MX2X1 g64084(.A (g_18795), .B (g_17934), .S0 (n_3174), .Y (n_3175));
DFFSRX1 g3976_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16659), .Q (g16693), .QN ());
OR2X1 g65275(.A (n_3171), .B (n_3121), .Y (n_3172));
NAND3X1 g61927(.A (n_1646), .B (g_20563), .C (n_9698), .Y (n_3170));
OAI21X1 g61399(.A0 (g1579), .A1 (n_9425), .B0 (n_3165), .Y (n_3167));
AOI21X1 g61952(.A0 (g_19172), .A1 (n_9775), .B0 (n_2574), .Y(n_3164));
AOI21X1 g61953(.A0 (g_11413), .A1 (n_9775), .B0 (n_2573), .Y(n_3162));
AOI21X1 g61954(.A0 (g_16456), .A1 (n_9884), .B0 (n_2572), .Y(n_3161));
AOI22X1 g65437(.A0 (n_2233), .A1 (n_1762), .B0 (g5180), .B1 (n_9129),.Y (n_3160));
AOI22X1 g65438(.A0 (n_2223), .A1 (n_1725), .B0 (g5873), .B1(n_10376), .Y (n_3158));
AOI22X1 g65440(.A0 (n_2219), .A1 (n_1723), .B0 (g6219), .B1 (n_9129),.Y (n_3157));
AOI22X1 g65443(.A0 (n_2225), .A1 (n_1743), .B0 (g3873), .B1 (n_9129),.Y (n_3156));
AOI22X1 g65446(.A0 (n_2203), .A1 (n_1758), .B0 (g3171), .B1 (n_9107),.Y (n_3154));
NAND4X1 g61957(.A (n_2867), .B (n_3152), .C (n_9359), .D (g4669), .Y(n_3153));
OR2X1 g63963(.A (n_3149), .B (n_3148), .Y (g26877));
OAI22X1 g65493(.A0 (n_2859), .A1 (n_1464), .B0 (n_621), .B1(n_10063), .Y (n_3147));
OAI22X1 g65494(.A0 (n_2855), .A1 (n_673), .B0 (n_686), .B1 (n_9830),.Y (n_3146));
OAI22X1 g65495(.A0 (n_2853), .A1 (n_1482), .B0 (n_623), .B1 (n_9830),.Y (n_3145));
OAI22X1 g65496(.A0 (n_2842), .A1 (n_1486), .B0 (n_603), .B1 (n_9830),.Y (n_3144));
MX2X1 g63084(.A (g5097), .B (n_2182), .S0 (n_10005), .Y (n_3143));
OAI22X1 g65497(.A0 (n_2849), .A1 (n_463), .B0 (n_664), .B1 (n_9992),.Y (n_3142));
OAI22X1 g65498(.A0 (n_2847), .A1 (n_458), .B0 (n_678), .B1 (n_9830),.Y (n_3141));
OAI22X1 g65501(.A0 (n_2857), .A1 (n_1459), .B0 (n_627), .B1(n_10063), .Y (n_3140));
MX2X1 g65530(.A (n_511), .B (g2980), .S0 (n_9269), .Y (n_3139));
MX2X1 g65531(.A (n_1633), .B (g_21651), .S0 (n_9599), .Y (n_3138));
MX2X1 g65532(.A (n_826), .B (n_6958), .S0 (n_9599), .Y (n_3137));
MX2X1 g65533(.A (n_209), .B (n_3135), .S0 (n_9599), .Y (n_3136));
DFFSRX1 g2927_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2509), .Q (), .QN (g2927));
DFFSRX1 g5448_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2517), .Q (g9555), .QN ());
DFFSRX1 g305_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2507), .Q (g_13901), .QN ());
DFFSRX1 g859_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2501), .Q (g14189), .QN ());
DFFSRX1 g2965_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2499), .Q (), .QN (g2965));
NOR2X1 g65624(.A (n_205), .B (n_9836), .Y (n_3133));
NOR2X1 g65641(.A (n_311), .B (n_9353), .Y (n_3132));
MX2X1 g63134(.A (g4269), .B (n_2181), .S0 (n_9000), .Y (n_3131));
NOR3X1 g65891(.A (n_276), .B (n_7247), .C (n_9505), .Y (n_3130));
NOR3X1 g65901(.A (n_11113), .B (n_9775), .C (g8719), .Y (n_3127));
INVX1 g61165(.A (n_3123), .Y (n_3124));
OAI21X1 g66057(.A0 (n_379), .A1 (n_9425), .B0 (n_3121), .Y (n_3122));
OAI21X1 g66063(.A0 (n_87), .A1 (n_9333), .B0 (n_2612), .Y (n_3120));
OAI21X1 g66066(.A0 (n_93), .A1 (n_9681), .B0 (n_3117), .Y (n_3119));
OAI21X1 g66067(.A0 (n_89), .A1 (n_9681), .B0 (n_3115), .Y (n_3116));
OAI21X1 g66068(.A0 (n_13), .A1 (n_9311), .B0 (n_3113), .Y (n_3114));
OAI21X1 g66078(.A0 (n_59), .A1 (n_9333), .B0 (n_2668), .Y (n_3112));
MX2X1 g66098(.A (g1798), .B (n_5996), .S0 (n_9269), .Y (n_3111));
MX2X1 g66099(.A (g1644), .B (g1592), .S0 (n_9599), .Y (n_3109));
MX2X1 g66105(.A (g2223), .B (n_5941), .S0 (n_9599), .Y (n_3108));
MX2X1 g66107(.A (g1913), .B (g1862), .S0 (n_9672), .Y (n_3106));
MX2X1 g66108(.A (g2912), .B (g2907), .S0 (n_9628), .Y (n_3105));
MX2X1 g66109(.A (g2994), .B (g2999), .S0 (n_9599), .Y (n_3104));
MX2X1 g66110(.A (g2204), .B (g2153), .S0 (n_9672), .Y (n_3103));
MX2X1 g66111(.A (g21292), .B (g_18015), .S0 (n_9269), .Y (n_3102));
MX2X1 g66112(.A (g2625), .B (n_5928), .S0 (n_9599), .Y (n_3100));
MX2X1 g66115(.A (g2047), .B (g1996), .S0 (n_9672), .Y (n_3099));
MX2X1 g66116(.A (g2066), .B (n_5932), .S0 (n_9628), .Y (n_3098));
MX2X1 g66117(.A (g1779), .B (g1728), .S0 (n_9019), .Y (n_3097));
MX2X1 g66122(.A (g2868), .B (g2988), .S0 (n_9599), .Y (n_3096));
MX2X1 g66123(.A (g4146), .B (g4176), .S0 (n_9269), .Y (n_3095));
MX2X1 g66127(.A (g4249), .B (g4253), .S0 (n_9269), .Y (n_3094));
MX2X1 g66130(.A (g4907), .B (g4922), .S0 (n_9599), .Y (n_3092));
MX2X1 g66132(.A (g2338), .B (g2287), .S0 (n_9672), .Y (n_3091));
MX2X1 g66134(.A (g2936), .B (g2922), .S0 (n_9599), .Y (n_3090));
MX2X1 g66135(.A (g4717), .B (g4732), .S0 (n_9269), .Y (n_3088));
MX2X1 g66136(.A (g4722), .B (g4717), .S0 (n_9269), .Y (n_3087));
MX2X1 g66139(.A (g1664), .B (n_5936), .S0 (n_9599), .Y (n_3086));
MX2X1 g66140(.A (g2357), .B (n_5917), .S0 (n_9599), .Y (n_3085));
MX2X1 g66141(.A (g2472), .B (g2421), .S0 (n_9019), .Y (n_3084));
MX2X1 g66142(.A (g2491), .B (n_5921), .S0 (n_9599), .Y (n_3082));
MX2X1 g66144(.A (g2922), .B (g2912), .S0 (n_9269), .Y (n_3081));
MX2X1 g66146(.A (g1932), .B (n_5925), .S0 (n_9599), .Y (n_3080));
MX2X1 g66149(.A (g2606), .B (g2555), .S0 (n_9628), .Y (n_3079));
MX2X1 g66154(.A (n_150), .B (g4273), .S0 (n_9019), .Y (n_3077));
XOR2X1 g61485(.A (n_8508), .B (n_2790), .Y (n_3075));
NAND4X1 g62097(.A (n_2925), .B (n_3073), .C (n_9139), .D (n_11216),.Y (n_3074));
INVX1 g66410(.A (n_3071), .Y (n_3072));
NOR2X1 g66656(.A (n_10956), .B (n_9353), .Y (n_3070));
AND2X1 g63454(.A (n_3431), .B (g_19414), .Y (n_3447));
DFFSRX1 g4917_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2512), .Q (g4917), .QN ());
DFFSRX1 g2890_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2493), .Q (g2890), .QN ());
DFFSRX1 g4108_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2498), .Q (g4108), .QN ());
DFFSRX1 g2759_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2510), .Q (g2759), .QN ());
DFFSRX1 g4082_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2503), .Q (g4082), .QN ());
OAI21X1 g63606(.A0 (n_3065), .A1 (n_7383), .B0 (n_2237), .Y (n_3066));
OAI21X1 g63614(.A0 (n_3062), .A1 (n_10889), .B0 (n_2264), .Y(n_3063));
DFFSRX1 g2735_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2491), .Q (g2735), .QN ());
DFFSRX1 g2715_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_9453), .Q (), .QN (g2715));
OR2X1 g61032(.A (n_4241), .B (g1413), .Y (n_3059));
MX2X1 g63772(.A (g_18793), .B (n_503), .S0 (n_3661), .Y (n_3058));
MX2X1 g63786(.A (g_21806), .B (n_2160), .S0 (n_9469), .Y (n_3057));
MX2X1 g63789(.A (g_22379), .B (n_2159), .S0 (n_9558), .Y (n_3056));
MX2X1 g63790(.A (n_11162), .B (n_2157), .S0 (n_9091), .Y (n_3055));
MX2X1 g63803(.A (g_6131), .B (n_2156), .S0 (n_9172), .Y (n_3053));
MX2X1 g63805(.A (g_20837), .B (n_2155), .S0 (n_9874), .Y (n_3052));
XOR2X1 g63810(.A (n_640), .B (n_2167), .Y (n_3713));
NOR2X1 g63906(.A (n_2743), .B (n_7260), .Y (n_3491));
NAND2X1 g63913(.A (n_3036), .B (n_3035), .Y (n_3497));
NAND4X1 g63968(.A (n_3048), .B (n_965), .C (n_3047), .D (n_2153), .Y(n_3050));
NAND4X1 g63995(.A (n_3048), .B (n_1630), .C (n_3047), .D (n_1263), .Y(n_3049));
NAND4X1 g64046(.A (n_2121), .B (n_1696), .C (n_2038), .D (n_2031), .Y(n_3044));
MX2X1 g64085(.A (n_3042), .B (g_18795), .S0 (n_3174), .Y (n_3043));
MX2X1 g64087(.A (g_12433), .B (g_20073), .S0 (n_3174), .Y (n_3041));
DFFSRX1 g6203_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2579), .Q (g6203), .QN ());
MX2X1 g64088(.A (n_10108), .B (n_3042), .S0 (n_3174), .Y (n_3040));
MX2X1 g64089(.A (g_20073), .B (n_10103), .S0 (n_3174), .Y (n_3038));
DFFSRX1 g4727_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2492), .Q (g4727), .QN ());
DFFSRX1 g2689_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2515), .Q (n_11099), .QN ());
DFFSRX1 g4076_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2502), .Q (g4076), .QN ());
DFFSRX1 g2130_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2504), .Q (g2130), .QN ());
DFFSRX1 g4104_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2514), .Q (g4104), .QN ());
OR2X1 g63949(.A (n_3036), .B (n_3035), .Y (g26876));
DFFSRX1 g4072_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_2454), .Q (), .QN (g4072));
MX2X1 g64086(.A (g_17934), .B (g_22464), .S0 (n_3174), .Y (n_3034));
NAND2X1 g64211(.A (g_15287), .B (n_10751), .Y (n_3033));
NAND3X1 g64213(.A (n_3031), .B (n_3030), .C (n_1250), .Y (n_3032));
NAND2X1 g64226(.A (n_1542), .B (n_2656), .Y (n_3029));
NOR2X1 g64242(.A (n_2453), .B (g_18795), .Y (n_3028));
NAND4X1 g64314(.A (n_2980), .B (n_3181), .C (n_9209), .D (g4633), .Y(n_3027));
NAND4X1 g64326(.A (n_1788), .B (n_3030), .C (n_3025), .D (n_2114), .Y(n_3026));
NAND4X1 g64368(.A (n_3030), .B (n_1266), .C (n_3021), .D (n_2116), .Y(n_3022));
XOR2X1 g64372(.A (n_3065), .B (n_7383), .Y (n_3020));
XOR2X1 g64373(.A (n_3062), .B (n_10889), .Y (n_3019));
MX2X1 g61747(.A (g_18902), .B (n_2346), .S0 (n_10063), .Y (n_3018));
NAND4X1 g64386(.A (n_3016), .B (n_3984), .C (n_10385), .D (g5037), .Y(n_3017));
AOI21X1 g64394(.A0 (n_2458), .A1 (n_9505), .B0 (n_2655), .Y (n_3015));
XOR2X1 g64403(.A (n_2415), .B (n_3013), .Y (n_3014));
XOR2X1 g64409(.A (n_2082), .B (n_2373), .Y (n_3660));
MX2X1 g64430(.A (n_3011), .B (n_1811), .S0 (n_9894), .Y (n_3012));
MX2X1 g64436(.A (g6163), .B (n_2375), .S0 (n_9359), .Y (n_3010));
MX2X1 g64441(.A (n_3007), .B (n_1795), .S0 (n_9553), .Y (n_3008));
MX2X1 g64460(.A (g1178), .B (n_2374), .S0 (n_9333), .Y (n_3005));
NOR2X1 g64508(.A (n_3003), .B (g_16792), .Y (n_3004));
NOR2X1 g64523(.A (n_2629), .B (n_644), .Y (n_3001));
INVX1 g64552(.A (n_7103), .Y (n_3838));
NAND2X1 g64583(.A (n_6577), .B (n_9448), .Y (n_3797));
CLKBUFX1 g64590(.A (n_2996), .Y (n_3239));
INVX1 g64616(.A (n_3612), .Y (n_5459));
INVX1 g64623(.A (n_3784), .Y (n_3626));
NAND3X1 g64630(.A (n_969), .B (n_2053), .C (n_9425), .Y (n_2989));
NAND4X1 g64632(.A (g5957), .B (n_11101), .C (g17715), .D (n_2421), .Y(n_2988));
INVX1 g64635(.A (n_2987), .Y (n_4053));
AND2X1 g64643(.A (n_2409), .B (g34034), .Y (n_3236));
NAND4X1 g64647(.A (g6649), .B (n_2600), .C (g17764), .D (n_11173), .Y(n_2986));
OR2X1 g64649(.A (n_10697), .B (g5052), .Y (n_2985));
NAND4X1 g64684(.A (n_3181), .B (n_10063), .C (n_2980), .D (n_974), .Y(n_2981));
NAND3X1 g61805(.A (n_830), .B (n_2002), .C (n_9425), .Y (n_2979));
NAND4X1 g64701(.A (g5256), .B (g25219), .C (g17639), .D (g25114), .Y(n_2977));
NAND4X1 g64709(.A (n_1163), .B (n_1668), .C (n_1712), .D (n_938), .Y(n_2975));
AOI22X1 g64710(.A0 (n_1813), .A1 (n_10078), .B0 (n_2973), .B1(g5152), .Y (n_2974));
NAND3X1 g61814(.A (n_848), .B (n_1994), .C (n_9209), .Y (n_2972));
NAND4X1 g64721(.A (n_2352), .B (g6295), .C (g17743), .D (n_11157), .Y(n_2971));
NAND4X1 g64723(.A (n_1226), .B (n_1715), .C (n_1672), .D (n_906), .Y(n_2969));
NAND4X1 g64735(.A (n_6806), .B (g3961), .C (g16659), .D (n_6786), .Y(n_2968));
NAND4X1 g64743(.A (n_1162), .B (n_1704), .C (n_1678), .D (n_915), .Y(n_2967));
NAND4X1 g64749(.A (n_2443), .B (g5603), .C (g17678), .D (n_1023), .Y(n_2966));
NAND4X1 g64759(.A (n_10623), .B (g5949), .C (g17715), .D (n_2376), .Y(n_2965));
NAND4X1 g64771(.A (n_2432), .B (g6641), .C (g17764), .D (n_11184), .Y(n_2964));
MX2X1 g64773(.A (g4939), .B (g4933), .S0 (n_2048), .Y (n_2963));
MX2X1 g64774(.A (g4749), .B (g4743), .S0 (n_2051), .Y (n_2962));
MX2X1 g64782(.A (g4698), .B (g4704), .S0 (n_2068), .Y (n_2961));
MX2X1 g64783(.A (g4754), .B (g4760), .S0 (n_2049), .Y (n_2960));
MX2X1 g64784(.A (g4765), .B (g4771), .S0 (n_2069), .Y (n_2959));
MX2X1 g64785(.A (g4944), .B (g4950), .S0 (n_2065), .Y (n_2958));
MX2X1 g64786(.A (g4955), .B (g4961), .S0 (n_2046), .Y (n_2957));
MX2X1 g64790(.A (g4492), .B (n_1563), .S0 (n_9240), .Y (n_2956));
MX2X1 g64791(.A (g4473), .B (n_1354), .S0 (n_9091), .Y (n_2955));
MX2X1 g64792(.A (g5084), .B (n_696), .S0 (n_9091), .Y (n_2954));
MX2X1 g64793(.A (g_18330), .B (n_469), .S0 (n_9834), .Y (n_2953));
MX2X1 g64794(.A (n_10524), .B (n_10535), .S0 (n_9256), .Y (n_2951));
MX2X1 g64795(.A (g4258), .B (n_695), .S0 (n_9172), .Y (n_2949));
MX2X1 g64796(.A (g_22552), .B (n_1095), .S0 (n_9940), .Y (n_2948));
MX2X1 g64797(.A (g1430), .B (n_652), .S0 (n_9894), .Y (n_2947));
NAND4X1 g62835(.A (n_2945), .B (n_9834), .C (n_2710), .D (n_1330), .Y(n_2946));
NAND2X1 g64850(.A (n_2061), .B (n_9398), .Y (n_3506));
NAND3X1 g64859(.A (n_2943), .B (n_4329), .C (n_10013), .Y (n_2944));
NAND2X1 g64860(.A (n_2785), .B (n_2784), .Y (n_2942));
NAND3X1 g64862(.A (n_2940), .B (n_4327), .C (n_9398), .Y (n_2941));
INVX1 g64864(.A (n_3224), .Y (n_3425));
NAND4X1 g62848(.A (n_2938), .B (n_9651), .C (n_2696), .D (n_1327), .Y(n_2939));
NAND3X1 g64867(.A (n_2936), .B (n_4324), .C (n_9466), .Y (n_2937));
NAND2X1 g64868(.A (n_2363), .B (n_2639), .Y (n_2934));
NAND3X1 g64869(.A (n_3253), .B (n_4316), .C (n_10950), .Y (n_2933));
NAND3X1 g64871(.A (n_2930), .B (n_4322), .C (n_9398), .Y (n_2931));
NAND3X1 g64876(.A (n_2928), .B (n_4320), .C (n_10013), .Y (n_2929));
OAI21X1 g62852(.A0 (n_2312), .A1 (g4854), .B0 (n_2925), .Y (n_2926));
NAND3X1 g64885(.A (n_2923), .B (n_4314), .C (n_9139), .Y (n_2924));
INVX2 g64950(.A (n_3003), .Y (n_3569));
NAND3X1 g64958(.A (n_2608), .B (g1448), .C (n_9698), .Y (n_2920));
INVX1 g61117(.A (n_10431), .Y (n_3910));
AOI21X1 g64993(.A0 (g16718), .A1 (n_238), .B0 (n_2348), .Y (n_2918));
AOI21X1 g64997(.A0 (g16744), .A1 (n_242), .B0 (n_2347), .Y (n_2917));
NAND4X1 g65031(.A (g16775), .B (g16659), .C (g11418), .D (g13966), .Y(n_3486));
MX2X1 g65081(.A (g2886), .B (n_992), .S0 (n_9311), .Y (n_2915));
MX2X1 g65086(.A (g5164), .B (n_1650), .S0 (n_9359), .Y (n_2914));
MX2X1 g65087(.A (g5511), .B (n_1649), .S0 (n_9750), .Y (n_2913));
MX2X1 g65088(.A (g6203), .B (n_1017), .S0 (n_9091), .Y (n_2912));
MX2X1 g65090(.A (g6549), .B (n_1396), .S0 (n_9091), .Y (n_2911));
MX2X1 g65091(.A (g3506), .B (n_1115), .S0 (n_9448), .Y (n_2910));
MX2X1 g65092(.A (g3155), .B (n_1109), .S0 (n_9091), .Y (n_2909));
MX2X1 g65094(.A (g3857), .B (n_1113), .S0 (n_9091), .Y (n_2907));
MX2X1 g65096(.A (g5857), .B (n_1002), .S0 (n_9091), .Y (n_2906));
MX2X1 g65097(.A (g5057), .B (n_2045), .S0 (n_9359), .Y (n_2905));
MX2X1 g65098(.A (n_1177), .B (n_1077), .S0 (n_9256), .Y (n_2904));
MX2X1 g65099(.A (n_1234), .B (n_1079), .S0 (n_9000), .Y (n_2903));
MX2X1 g65100(.A (g4308), .B (n_1570), .S0 (n_9834), .Y (n_2902));
MX2X1 g65101(.A (n_1169), .B (n_1069), .S0 (n_9091), .Y (n_2900));
MX2X1 g65102(.A (n_1214), .B (n_1072), .S0 (n_9000), .Y (n_2898));
MX2X1 g65103(.A (n_1135), .B (n_1075), .S0 (n_9750), .Y (n_2897));
MX2X1 g65104(.A (g_16571), .B (n_1081), .S0 (n_9240), .Y (n_2896));
MX2X1 g65105(.A (g4291), .B (n_1556), .S0 (n_9358), .Y (n_2895));
MX2X1 g65106(.A (n_1210), .B (n_1074), .S0 (n_8955), .Y (n_2894));
MX2X1 g65108(.A (n_1191), .B (n_998), .S0 (n_9167), .Y (n_2892));
MX2X1 g65109(.A (g_17426), .B (g_10278), .S0 (n_3177), .Y (n_2891));
MX2X1 g65110(.A (g4281), .B (n_1820), .S0 (n_9091), .Y (n_2890));
MX2X1 g65111(.A (g1306), .B (n_1997), .S0 (n_9000), .Y (n_2889));
MX2X1 g65112(.A (n_1216), .B (n_1071), .S0 (n_9750), .Y (n_2888));
MX2X1 g65113(.A (g1183), .B (n_1991), .S0 (n_9359), .Y (n_2887));
MX2X1 g65114(.A (g_15758), .B (n_1992), .S0 (n_8955), .Y (n_2886));
NAND3X1 g65260(.A (g_19911), .B (n_3323), .C (n_9501), .Y (n_2885));
INVX1 g65264(.A (n_2883), .Y (n_2884));
NOR2X1 g65276(.A (n_2881), .B (n_2838), .Y (n_2882));
NOR2X1 g65278(.A (n_6398), .B (n_2319), .Y (n_2880));
NAND3X1 g61929(.A (g_18902), .B (n_2878), .C (n_9750), .Y (n_2879));
NAND3X1 g65348(.A (g1345), .B (n_3459), .C (n_10063), .Y (n_2875));
NOR2X1 g65371(.A (n_2871), .B (n_2835), .Y (n_2872));
NAND3X1 g61943(.A (n_2003), .B (g_18869), .C (n_9091), .Y (n_2870));
NOR2X1 g65419(.A (g16775), .B (n_2594), .Y (n_2869));
OR4X1 g61951(.A (n_2867), .B (n_2410), .C (n_9129), .D (g4669), .Y(n_2868));
NAND3X1 g65422(.A (n_987), .B (n_986), .C (n_10005), .Y (n_2866));
OAI22X1 g65500(.A0 (n_2578), .A1 (n_1468), .B0 (n_612), .B1(n_10063), .Y (n_2864));
OAI22X1 g65503(.A0 (n_2862), .A1 (g4473), .B0 (n_2861), .B1 (n_9830),.Y (n_2863));
NOR2X1 g65698(.A (n_2859), .B (g5164), .Y (n_2860));
NOR2X1 g65704(.A (n_2857), .B (g5857), .Y (n_2858));
NOR2X1 g65711(.A (n_2855), .B (g5511), .Y (n_2856));
NOR2X1 g65737(.A (n_2853), .B (g3155), .Y (n_2854));
NAND3X1 g65769(.A (g_16404), .B (g_16571), .C (n_9651), .Y (n_2852));
NOR2X1 g65773(.A (n_2849), .B (g3506), .Y (n_2850));
NOR2X1 g65811(.A (n_2847), .B (g3857), .Y (n_2848));
MX2X1 g61435(.A (n_8508), .B (n_1351), .S0 (n_9000), .Y (n_2846));
NOR2X1 g62013(.A (n_2174), .B (g4939), .Y (n_2845));
NOR2X1 g62014(.A (n_2173), .B (g4950), .Y (n_2844));
NOR2X1 g65874(.A (n_2842), .B (g6549), .Y (n_2843));
NAND2X1 g61162(.A (n_10242), .B (n_2176), .Y (n_2841));
OAI21X1 g65951(.A0 (g_18015), .A1 (n_2518), .B0 (n_9351), .Y(n_2840));
OAI21X1 g66005(.A0 (n_144), .A1 (n_9311), .B0 (n_2838), .Y (n_2839));
OAI21X1 g66007(.A0 (n_1), .A1 (n_9422), .B0 (n_2835), .Y (n_2837));
NAND2X1 g61164(.A (n_2180), .B (n_10243), .Y (n_2834));
OAI21X1 g66019(.A0 (n_127), .A1 (n_9422), .B0 (n_2606), .Y (n_2833));
MX2X1 g66124(.A (g4146), .B (g4157), .S0 (n_9240), .Y (n_2832));
OAI21X1 g66029(.A0 (n_39), .A1 (n_9425), .B0 (n_2661), .Y (n_2831));
AOI21X1 g61166(.A0 (n_2), .A1 (n_1275), .B0 (n_2830), .Y (n_3123));
OAI21X1 g66040(.A0 (n_117), .A1 (n_9425), .B0 (n_2828), .Y (n_2829));
OAI22X1 g66096(.A0 (n_10280), .A1 (n_9627), .B0 (n_169), .B1(n_9672), .Y (n_2827));
MX2X1 g66097(.A (g2844), .B (g2852), .S0 (n_9000), .Y (n_2826));
MX2X1 g66101(.A (g2936), .B (g2950), .S0 (n_10005), .Y (n_2824));
MX2X1 g66102(.A (g4722), .B (g4737), .S0 (n_8955), .Y (n_2823));
MX2X1 g66103(.A (g2852), .B (g2860), .S0 (n_9091), .Y (n_2822));
MX2X1 g66106(.A (g2890), .B (g2844), .S0 (n_9000), .Y (n_2821));
MX2X1 g66113(.A (g2860), .B (g2894), .S0 (n_9000), .Y (n_2820));
MX2X1 g66114(.A (g2894), .B (n_22), .S0 (n_9172), .Y (n_2819));
MX2X1 g66118(.A (g2950), .B (g2960), .S0 (n_9311), .Y (n_2817));
MX2X1 g66119(.A (g2868), .B (g2873), .S0 (n_9234), .Y (n_2816));
MX2X1 g66120(.A (g2130), .B (g2138), .S0 (n_9091), .Y (n_2815));
OAI22X1 g66121(.A0 (n_1240), .A1 (n_10385), .B0 (n_308), .B1(n_9903), .Y (n_2814));
MX2X1 g66126(.A (g4249), .B (g4245), .S0 (n_9333), .Y (n_2813));
MX2X1 g66128(.A (g4300), .B (g4253), .S0 (n_9311), .Y (n_2812));
MX2X1 g66129(.A (n_22), .B (g20652), .S0 (n_9834), .Y (n_2810));
OR4X1 g62078(.A (n_2925), .B (n_2361), .C (n_9404), .D (n_11216), .Y(n_2809));
MX2X1 g66133(.A (g2960), .B (g2970), .S0 (n_9167), .Y (n_2808));
MX2X1 g66137(.A (n_11097), .B (g2697), .S0 (n_9091), .Y (n_2807));
MX2X1 g66138(.A (g4727), .B (g4732), .S0 (n_9172), .Y (n_2806));
MX2X1 g66143(.A (g2984), .B (g2907), .S0 (n_9311), .Y (n_2805));
MX2X1 g66145(.A (g4907), .B (g4912), .S0 (n_9834), .Y (n_2804));
MX2X1 g66147(.A (g4917), .B (g4922), .S0 (n_9234), .Y (n_2803));
MX2X1 g66148(.A (g4912), .B (g4927), .S0 (n_9256), .Y (n_2802));
MX2X1 g61486(.A (g4430), .B (n_1315), .S0 (n_8955), .Y (n_2801));
NAND2X1 g66280(.A (n_10112), .B (n_9431), .Y (n_2800));
NAND2X1 g66322(.A (n_10188), .B (n_9371), .Y (n_2798));
NAND2X1 g66323(.A (n_3914), .B (n_9431), .Y (n_2797));
AND2X1 g66398(.A (n_8895), .B (n_9019), .Y (n_2796));
NAND2X1 g66401(.A (n_926), .B (n_9884), .Y (n_2795));
NAND2X1 g66411(.A (n_2861), .B (n_9940), .Y (n_3071));
NAND2X1 g66412(.A (g1367), .B (n_9772), .Y (n_2794));
AND2X1 g66419(.A (g4153), .B (n_9672), .Y (n_2793));
NAND2X1 g61498(.A (n_2790), .B (n_1986), .Y (n_2791));
AND2X1 g66439(.A (g2975), .B (n_9672), .Y (n_2789));
AND2X1 g66443(.A (g4104), .B (n_9672), .Y (n_2788));
AND2X1 g66464(.A (g4087), .B (n_9672), .Y (n_2787));
OR2X1 g64887(.A (n_2785), .B (n_2784), .Y (g28041));
NAND2X1 g66525(.A (g_22306), .B (n_9419), .Y (n_2783));
NOR2X1 g66541(.A (g4258), .B (n_9772), .Y (n_2782));
NAND2X1 g66543(.A (n_2780), .B (n_9836), .Y (n_2781));
NAND2X1 g66549(.A (g1345), .B (n_9505), .Y (n_2779));
NAND2X1 g66557(.A (n_662), .B (n_9952), .Y (n_2778));
AND2X1 g66611(.A (g5188), .B (n_9448), .Y (n_2777));
NOR2X1 g66698(.A (n_553), .B (n_9353), .Y (n_2776));
NAND2X1 g66715(.A (g2882), .B (n_9952), .Y (n_2775));
NAND2X1 g63451(.A (n_2483), .B (n_10818), .Y (n_3651));
MX2X1 g61182(.A (n_2773), .B (n_1869), .S0 (n_8955), .Y (n_2774));
AND2X1 g66753(.A (g6573), .B (n_9698), .Y (n_2772));
AND2X1 g66807(.A (g3881), .B (n_9448), .Y (n_2770));
AND2X1 g66823(.A (g3530), .B (n_9448), .Y (n_2769));
NOR2X1 g66852(.A (n_10557), .B (n_9775), .Y (n_2768));
NAND2X1 g66853(.A (n_955), .B (n_9952), .Y (n_2767));
AND2X1 g66879(.A (g5881), .B (n_9448), .Y (n_2766));
NOR2X1 g66909(.A (n_617), .B (n_9019), .Y (n_2765));
NAND4X1 g63529(.A (n_1597), .B (n_10112), .C (n_9883), .D (n_392), .Y(n_2764));
NAND2X1 g61568(.A (n_9811), .B (g12919), .Y (n_3316));
MX2X1 g66100(.A (g2994), .B (g2988), .S0 (n_9000), .Y (n_2762));
MX2X1 g63787(.A (g5092), .B (n_1590), .S0 (n_10005), .Y (n_2761));
MX2X1 g63788(.A (n_10128), .B (n_1842), .S0 (n_9797), .Y (n_2760));
MX2X1 g63798(.A (g4264), .B (n_1839), .S0 (n_9000), .Y (n_2759));
MX2X1 g63806(.A (g1548), .B (n_1296), .S0 (n_9358), .Y (n_2758));
NAND2X1 g63899(.A (n_2465), .B (n_684), .Y (n_3563));
OR2X1 g63903(.A (n_3844), .B (g_6283), .Y (n_2757));
NAND4X1 g64057(.A (n_2129), .B (n_1669), .C (n_1717), .D (n_1694), .Y(n_2756));
NAND4X1 g64058(.A (n_1846), .B (n_1857), .C (n_1844), .D (n_1699), .Y(n_2755));
INVX1 g64092(.A (n_2754), .Y (n_3332));
MX2X1 g64096(.A (n_276), .B (n_2090), .S0 (n_8955), .Y (n_2753));
OR2X1 g64139(.A (n_3174), .B (n_83), .Y (n_2751));
OAI21X1 g64143(.A0 (n_2945), .A1 (n_10753), .B0 (n_10005), .Y(n_2749));
AOI21X1 g64150(.A0 (n_2110), .A1 (n_344), .B0 (n_643), .Y (n_2748));
NAND3X1 g64165(.A (n_2457), .B (n_2456), .C (n_2747), .Y (n_3502));
OR4X1 g64247(.A (n_2980), .B (n_276), .C (n_9129), .D (g4633), .Y(n_2746));
NAND2X1 g64259(.A (n_3174), .B (g_21576), .Y (n_2744));
INVX1 g64282(.A (n_2743), .Y (n_3493));
NAND2X1 g61730(.A (n_2430), .B (n_10005), .Y (n_2742));
NOR2X1 g64323(.A (n_1632), .B (n_2154), .Y (n_2741));
NAND3X1 g64327(.A (n_1658), .B (n_1887), .C (n_9209), .Y (n_2740));
MX2X1 g61295(.A (g1404), .B (n_1569), .S0 (n_9091), .Y (n_2739));
NAND4X1 g64362(.A (n_1193), .B (n_1689), .C (n_1707), .D (n_932), .Y(n_2738));
OAI21X1 g64388(.A0 (n_3171), .A1 (n_1695), .B0 (n_2302), .Y (n_2736));
OAI21X1 g64389(.A0 (n_2881), .A1 (n_2734), .B0 (n_2241), .Y (n_2735));
OAI21X1 g64390(.A0 (n_2732), .A1 (n_2421), .B0 (n_2289), .Y (n_2733));
OAI21X1 g64391(.A0 (n_2729), .A1 (n_11150), .B0 (n_2277), .Y(n_2730));
OAI21X1 g64392(.A0 (n_2871), .A1 (n_11173), .B0 (n_2274), .Y(n_2727));
MX2X1 g61750(.A (n_2429), .B (n_2032), .S0 (n_9797), .Y (n_2725));
MX2X1 g64425(.A (g5156), .B (n_1792), .S0 (n_9333), .Y (n_2722));
MX2X1 g64426(.A (g5124), .B (n_2087), .S0 (n_9240), .Y (n_2720));
MX2X1 g64427(.A (n_2718), .B (n_1814), .S0 (n_9797), .Y (n_2719));
MX2X1 g64428(.A (n_2943), .B (n_1798), .S0 (n_9000), .Y (n_2716));
MX2X1 g64429(.A (g5471), .B (n_2098), .S0 (n_9091), .Y (n_2715));
MX2X1 g64432(.A (n_2940), .B (n_1809), .S0 (n_9992), .Y (n_2714));
MX2X1 g64433(.A (g5817), .B (n_2097), .S0 (n_9091), .Y (n_2713));
MX2X1 g64435(.A (n_2936), .B (n_2086), .S0 (n_9091), .Y (n_2712));
NAND4X1 g62668(.A (n_2710), .B (n_2945), .C (n_9664), .D (n_8799), .Y(n_2711));
MX2X1 g64438(.A (g3115), .B (n_2092), .S0 (n_9311), .Y (n_2709));
MX2X1 g64439(.A (n_2930), .B (n_1803), .S0 (n_9156), .Y (n_2707));
MX2X1 g64440(.A (g6509), .B (n_2095), .S0 (n_9091), .Y (n_2706));
MX2X1 g64443(.A (n_2704), .B (n_2085), .S0 (n_9000), .Y (n_2705));
MX2X1 g64444(.A (n_2928), .B (n_1801), .S0 (n_9167), .Y (n_2703));
MX2X1 g64445(.A (g3466), .B (n_2091), .S0 (n_9627), .Y (n_2702));
MX2X1 g64446(.A (n_2699), .B (n_1800), .S0 (n_9000), .Y (n_2700));
NAND4X1 g62674(.A (n_2696), .B (n_2938), .C (n_9992), .D (g1554), .Y(n_2697));
MX2X1 g64448(.A (n_2923), .B (n_1843), .S0 (n_9156), .Y (n_2695));
MX2X1 g64449(.A (g3817), .B (n_2093), .S0 (n_9664), .Y (n_2694));
MX2X1 g64450(.A (n_2692), .B (n_1797), .S0 (n_9000), .Y (n_2693));
MX2X1 g64451(.A (g_14535), .B (n_2083), .S0 (n_9218), .Y (n_2691));
MX2X1 g64452(.A (n_2005), .B (n_1793), .S0 (n_9797), .Y (n_2690));
MX2X1 g64454(.A (g4245), .B (n_1821), .S0 (n_9240), .Y (n_2689));
MX2X1 g64455(.A (g1489), .B (n_1804), .S0 (n_9359), .Y (n_2688));
MX2X1 g64456(.A (n_2686), .B (n_1806), .S0 (n_9256), .Y (n_2687));
MX2X1 g64458(.A (n_2684), .B (n_1808), .S0 (n_8955), .Y (n_2685));
AND2X1 g64507(.A (n_10526), .B (g_12791), .Y (n_3291));
NOR2X1 g64510(.A (n_1571), .B (n_9353), .Y (n_2682));
NAND2X1 g64517(.A (n_3152), .B (n_9209), .Y (n_3489));
AOI21X1 g64526(.A0 (n_2679), .A1 (n_3984), .B0 (n_10134), .Y(n_2680));
OR2X1 g64530(.A (n_2426), .B (n_2677), .Y (n_2678));
NAND2X1 g64547(.A (n_6695), .B (n_9627), .Y (n_2675));
NOR2X1 g64548(.A (n_1268), .B (n_2406), .Y (n_2673));
XOR2X1 g61328(.A (g1404), .B (n_2671), .Y (n_2672));
NOR2X1 g64557(.A (n_3062), .B (n_2668), .Y (n_2669));
INVX2 g64563(.A (n_11207), .Y (n_6243));
NAND3X1 g64584(.A (n_981), .B (n_1756), .C (n_9091), .Y (n_2666));
NAND3X1 g64585(.A (n_849), .B (n_2056), .C (n_9558), .Y (n_2665));
AND2X1 g64591(.A (n_2387), .B (g34036), .Y (n_2996));
NAND2X1 g64603(.A (n_3152), .B (n_988), .Y (n_2664));
NOR2X1 g64606(.A (n_2630), .B (n_1549), .Y (n_2663));
NOR2X1 g64626(.A (n_3065), .B (n_2661), .Y (n_2662));
NAND4X1 g64627(.A (g5611), .B (n_2597), .C (g17678), .D (n_2208), .Y(n_2660));
NAND4X1 g64629(.A (g6303), .B (n_2325), .C (g17743), .D (n_11150), .Y(n_2659));
NAND2X1 g64631(.A (n_2118), .B (n_2657), .Y (n_2658));
INVX1 g64636(.A (n_6765), .Y (n_2987));
NAND4X1 g64662(.A (n_777), .B (n_1541), .C (n_1548), .D (n_2452), .Y(n_2656));
NOR2X1 g64663(.A (n_1976), .B (n_2654), .Y (n_2655));
NAND4X1 g64716(.A (n_8586), .B (g3259), .C (g16603), .D (n_8548), .Y(n_2653));
NAND4X1 g64736(.A (n_10879), .B (g3610), .C (g16627), .D (n_4682), .Y(n_2652));
NAND4X1 g64737(.A (n_920), .B (n_1530), .C (n_1521), .D (n_704), .Y(n_2651));
XOR2X1 g64788(.A (g8358), .B (n_1733), .Y (n_2648));
INVX1 g64817(.A (g5339), .Y (n_2647));
INVX1 g64819(.A (g6377), .Y (n_2646));
INVX1 g64828(.A (g5685), .Y (n_2645));
INVX1 g64830(.A (g6723), .Y (n_2644));
INVX1 g64833(.A (g6031), .Y (n_2642));
NAND2X1 g64841(.A (n_2640), .B (g_8896), .Y (n_2641));
NOR2X1 g64865(.A (n_2640), .B (n_2639), .Y (n_3224));
OR2X1 g64873(.A (n_2042), .B (g5041), .Y (n_2638));
NAND2X2 g64906(.A (n_11192), .B (n_11193), .Y (n_3259));
NAND2X1 g64907(.A (n_2034), .B (n_1682), .Y (n_2637));
NAND3X1 g64937(.A (n_2057), .B (g1478), .C (n_9811), .Y (n_2634));
NAND3X1 g64938(.A (n_2054), .B (g1300), .C (n_9558), .Y (n_2632));
BUFX3 g64951(.A (n_10526), .Y (n_3003));
NOR2X1 g64965(.A (n_1975), .B (n_8694), .Y (n_2629));
AOI21X1 g64967(.A0 (n_1363), .A1 (n_10813), .B0 (n_3177), .Y(n_2628));
AND2X1 g64970(.A (n_2070), .B (n_6970), .Y (n_3016));
XOR2X1 g64982(.A (n_2871), .B (n_11171), .Y (n_2625));
XOR2X1 g64985(.A (n_2881), .B (n_2224), .Y (n_2624));
NAND2X1 g61371(.A (g4427), .B (n_9129), .Y (n_2619));
DFFSRX1 g3274_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16603), .Q (g16624), .QN ());
DFFSRX1 g3625_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16627), .Q (g16656), .QN ());
NAND2X1 g65236(.A (g26801), .B (n_9750), .Y (n_2616));
OR2X1 g65241(.A (n_4316), .B (n_9772), .Y (n_2615));
NOR2X1 g65248(.A (n_1576), .B (n_9193), .Y (n_4091));
OAI21X1 g65254(.A0 (n_276), .A1 (n_10402), .B0 (n_9894), .Y (n_2614));
NOR2X1 g65265(.A (n_3177), .B (n_3391), .Y (n_2883));
NOR2X1 g65280(.A (n_2732), .B (n_2612), .Y (n_2613));
NAND2X1 g65292(.A (n_6404), .B (n_6395), .Y (n_6400));
NAND2X1 g65324(.A (n_3184), .B (n_10524), .Y (n_2611));
NOR2X1 g65328(.A (n_4617), .B (n_10078), .Y (n_2610));
INVX1 g65346(.A (n_2608), .Y (n_2609));
NOR2X1 g65351(.A (n_2729), .B (n_2606), .Y (n_2607));
NAND2X1 g66420(.A (g4664), .B (n_9884), .Y (n_2604));
NAND3X1 g61949(.A (n_1993), .B (g_11413), .C (n_9311), .Y (n_2603));
OR2X1 g65430(.A (n_2004), .B (n_10184), .Y (n_2602));
NAND4X1 g65473(.A (g6585), .B (n_2600), .C (g12470), .D (n_11171), .Y(n_2601));
NAND4X1 g65477(.A (g5547), .B (n_2597), .C (g12300), .D (n_1023), .Y(n_2598));
OAI21X1 g65502(.A0 (g1442), .A1 (n_9599), .B0 (n_2006), .Y (n_2595));
NAND2X1 g61149(.A (n_2592), .B (g1542), .Y (n_4241));
OR2X1 g61150(.A (n_2592), .B (g1542), .Y (n_2593));
NAND3X1 g65687(.A (n_1356), .B (n_9811), .C (n_107), .Y (n_2590));
OR2X1 g65690(.A (g5112), .B (n_9398), .Y (n_2589));
NOR2X1 g65700(.A (n_1058), .B (n_9107), .Y (n_2588));
OAI21X1 g64021(.A0 (n_1826), .A1 (g4849), .B0 (n_1875), .Y (n_2587));
AND2X1 g61154(.A (n_6781), .B (n_11042), .Y (n_3183));
NOR2X1 g65803(.A (n_1982), .B (n_16), .Y (n_2586));
NOR2X1 g65823(.A (n_1979), .B (n_40), .Y (n_2585));
NAND2X1 g65876(.A (n_2583), .B (n_3857), .Y (n_2584));
NOR2X1 g65887(.A (n_1971), .B (g4616), .Y (n_2582));
INVX1 g65895(.A (n_2580), .Y (n_2581));
NOR2X1 g65908(.A (n_2578), .B (g6203), .Y (n_2579));
NAND2X1 g65953(.A (n_2481), .B (n_2480), .Y (n_2575));
NAND2X1 g61463(.A (n_9359), .B (g12923), .Y (n_3165));
NOR2X1 g62058(.A (n_1969), .B (n_4764), .Y (n_2574));
NOR2X1 g62064(.A (n_2000), .B (n_4761), .Y (n_2573));
NOR2X1 g62065(.A (n_1977), .B (n_4757), .Y (n_2572));
NAND2X1 g66302(.A (n_2566), .B (n_9466), .Y (n_2567));
NAND2X1 g66306(.A (g4608), .B (n_9431), .Y (n_2564));
INVX1 g66309(.A (n_2562), .Y (n_2563));
NAND2X1 g66318(.A (g5813), .B (n_9775), .Y (n_2560));
OR2X1 g66330(.A (n_9672), .B (g10122), .Y (n_2559));
NAND2X1 g66334(.A (g2227), .B (n_9672), .Y (n_2558));
NAND2X1 g66365(.A (n_2556), .B (n_9107), .Y (n_2557));
NAND2X1 g66374(.A (g1384), .B (n_9505), .Y (n_2555));
NOR2X1 g66393(.A (n_10314), .B (n_10716), .Y (n_2554));
NAND2X1 g66397(.A (n_2550), .B (n_9836), .Y (n_2551));
NAND2X1 g66405(.A (g_12465), .B (n_9976), .Y (n_2548));
NOR2X1 g66406(.A (g_18112), .B (n_10376), .Y (n_2546));
NAND2X1 g66413(.A (g4628), .B (n_9599), .Y (n_2545));
NAND2X1 g66438(.A (g_14342), .B (n_9928), .Y (n_2543));
NAND2X1 g66463(.A (g6159), .B (n_9599), .Y (n_2540));
NAND2X1 g66472(.A (n_2538), .B (n_10952), .Y (n_2539));
NAND2X1 g66482(.A (g2236), .B (n_9300), .Y (n_2537));
NAND2X1 g66495(.A (n_2535), .B (n_9193), .Y (n_2536));
NAND2X1 g66501(.A (n_4339), .B (n_9952), .Y (n_2533));
NAND2X1 g66509(.A (g_19304), .B (n_9300), .Y (n_2531));
NAND2X1 g66510(.A (n_2529), .B (n_9628), .Y (n_2530));
NAND2X1 g66522(.A (g_16958), .B (n_10078), .Y (n_2528));
NAND2X1 g66533(.A (g_20159), .B (n_9836), .Y (n_2526));
NAND2X1 g66540(.A (g2638), .B (n_9300), .Y (n_2524));
NAND2X1 g66555(.A (g1677), .B (n_9505), .Y (n_2523));
NAND2X1 g66561(.A (n_2521), .B (n_10952), .Y (n_2522));
NAND2X1 g66565(.A (n_8913), .B (n_9884), .Y (n_2520));
NOR2X1 g66602(.A (n_9836), .B (n_2518), .Y (n_2519));
AND2X1 g66636(.A (g5535), .B (n_9698), .Y (n_2517));
NAND2X1 g66643(.A (n_9553), .B (g6748), .Y (n_3117));
NAND2X1 g66672(.A (g25219), .B (n_9139), .Y (n_3121));
AND2X1 g66676(.A (n_11097), .B (n_9717), .Y (n_2515));
OR2X1 g66684(.A (g4108), .B (n_9627), .Y (n_2514));
AND2X1 g66695(.A (g4917), .B (n_9501), .Y (n_2512));
OR2X1 g66697(.A (g2756), .B (n_9453), .Y (n_2510));
OR2X1 g66701(.A (n_3463), .B (n_9627), .Y (n_2509));
NAND2X1 g66707(.A (n_9553), .B (g6750), .Y (n_3113));
AND2X1 g66714(.A (n_9501), .B (g6745), .Y (n_2507));
NOR2X1 g66727(.A (n_365), .B (n_9884), .Y (n_2506));
AND2X1 g66744(.A (g2130), .B (n_9717), .Y (n_2504));
OR2X1 g66745(.A (g4141), .B (n_9501), .Y (n_2503));
OR2X1 g66750(.A (g4082), .B (n_9627), .Y (n_2502));
AND2X1 g66751(.A (n_9501), .B (g21176), .Y (n_2501));
NOR2X1 g66763(.A (n_383), .B (n_9107), .Y (n_2500));
OR2X1 g66810(.A (g2955), .B (n_9398), .Y (n_2499));
NAND2X1 g66840(.A (n_9627), .B (g6749), .Y (n_3115));
OR2X1 g66844(.A (g4098), .B (n_9627), .Y (n_2498));
INVX1 g66858(.A (n_2496), .Y (n_2497));
NOR2X1 g66893(.A (g_18200), .B (n_9107), .Y (n_2495));
NOR2X1 g66894(.A (n_261), .B (n_10078), .Y (n_2494));
OR2X1 g66897(.A (g2873), .B (n_9501), .Y (n_2493));
AND2X1 g66903(.A (g4727), .B (n_10005), .Y (n_2492));
OR2X1 g66905(.A (n_10650), .B (n_9501), .Y (n_2491));
NAND2X1 g61530(.A (g23683), .B (n_9772), .Y (n_2488));
NAND2X1 g66544(.A (n_2485), .B (n_9628), .Y (n_2486));
XOR2X1 g64079(.A (n_221), .B (n_2165), .Y (n_2484));
INVX1 g64093(.A (n_2483), .Y (n_2754));
OR2X1 g65969(.A (n_2481), .B (n_2480), .Y (g28042));
NAND2X1 g64151(.A (n_1863), .B (n_10949), .Y (n_3148));
NAND4X1 g64185(.A (n_1567), .B (n_1822), .C (n_11051), .D (n_273), .Y(n_2479));
NAND2X1 g64237(.A (n_1862), .B (n_10687), .Y (n_3036));
NAND2X1 g64253(.A (n_1861), .B (n_10949), .Y (n_3035));
NAND2X1 g64261(.A (n_2152), .B (n_9862), .Y (n_3149));
AOI21X1 g64283(.A0 (n_1429), .A1 (n_1832), .B0 (n_1838), .Y (n_2743));
OAI21X1 g61288(.A0 (n_2062), .A1 (n_2474), .B0 (n_2063), .Y (n_2475));
NAND4X1 g64363(.A (n_925), .B (n_1516), .C (n_1525), .D (n_927), .Y(n_2472));
AOI22X1 g64364(.A0 (n_1791), .A1 (n_448), .B0 (n_797), .B1 (g4311),.Y (n_2471));
NAND4X1 g64366(.A (n_929), .B (n_1511), .C (n_1534), .D (n_894), .Y(n_2469));
AOI21X1 g64393(.A0 (n_10664), .A1 (n_1538), .B0 (n_2151), .Y(n_2468));
NAND4X1 g64405(.A (n_934), .B (n_1507), .C (n_1523), .D (n_895), .Y(n_2466));
INVX1 g64413(.A (n_2465), .Y (n_2723));
NOR2X1 g64511(.A (n_10496), .B (n_10525), .Y (n_3431));
OR2X1 g64513(.A (n_2096), .B (n_10952), .Y (n_2464));
OR2X1 g64514(.A (n_2094), .B (n_9193), .Y (n_2463));
OR2X1 g64516(.A (n_2089), .B (n_9193), .Y (n_2461));
OR2X1 g64518(.A (n_2088), .B (n_9491), .Y (n_2460));
NAND3X1 g64550(.A (n_2458), .B (n_10725), .C (n_10063), .Y (n_2459));
AND2X1 g64554(.A (n_2457), .B (n_2456), .Y (n_3031));
AND2X1 g64576(.A (n_2103), .B (n_10005), .Y (n_2454));
NAND2X1 g64592(.A (n_2107), .B (g_17934), .Y (n_2453));
OR2X1 g64888(.A (n_1736), .B (n_2449), .Y (g26875));
NAND4X1 g64702(.A (n_2447), .B (g3937), .C (g16775), .D (n_8917), .Y(n_2448));
NAND4X1 g64742(.A (n_1494), .B (n_2443), .C (g17711), .D (g5591), .Y(n_2444));
INVX1 g64745(.A (n_2134), .Y (n_2442));
NAND4X1 g64747(.A (n_1494), .B (n_2439), .C (g17580), .D (g5607), .Y(n_2441));
NAND4X1 g64748(.A (n_7150), .B (g5575), .C (g14694), .D (n_1494), .Y(n_2438));
INVX1 g64766(.A (n_2120), .Y (n_2437));
NAND4X1 g64768(.A (n_2433), .B (n_2435), .C (g17688), .D (g6645), .Y(n_2436));
NAND4X1 g64769(.A (n_2433), .B (n_2432), .C (g17778), .D (g6629), .Y(n_2434));
NAND4X1 g64770(.A (n_2433), .B (g6613), .C (g14828), .D (n_3275), .Y(n_2431));
OAI21X1 g61838(.A0 (n_2345), .A1 (n_2429), .B0 (n_1645), .Y (n_2430));
DFFSRX1 g5339_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17639), .Q (g5339), .QN ());
DFFSRX1 g6377_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17743), .Q (g6377), .QN ());
DFFSRX1 g5685_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17678), .Q (g5685), .QN ());
DFFSRX1 g6723_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17764), .Q (g6723), .QN ());
DFFSRX1 g6031_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17715), .Q (g6031), .QN ());
NAND2X1 g64838(.A (n_2427), .B (g1199), .Y (n_3844));
OR2X1 g64839(.A (n_2427), .B (g1199), .Y (n_2428));
NAND2X1 g64842(.A (n_2449), .B (n_38), .Y (n_2426));
OR2X1 g64845(.A (n_891), .B (n_9526), .Y (n_2425));
NAND4X1 g64856(.A (n_2421), .B (g5941), .C (g14673), .D (n_10808), .Y(n_2423));
INVX1 g64857(.A (n_10268), .Y (g27831));
NAND2X1 g66449(.A (g2079), .B (n_9371), .Y (n_2419));
NAND4X1 g64893(.A (n_1785), .B (n_946), .C (g4698), .D (n_10225), .Y(n_2416));
NAND2X1 g64909(.A (n_1680), .B (n_1675), .Y (n_2415));
NAND2X1 g64910(.A (n_1674), .B (n_1681), .Y (n_3013));
NAND4X1 g64917(.A (n_2413), .B (g6287), .C (g14705), .D (n_11150), .Y(n_2414));
INVX1 g64921(.A (n_2410), .Y (n_3152));
NAND4X1 g64927(.A (n_1786), .B (n_11133), .C (g4888), .D (n_740), .Y(n_2409));
NOR2X1 g64928(.A (n_2061), .B (n_598), .Y (n_2465));
NAND4X1 g64929(.A (n_2435), .B (g6633), .C (g14749), .D (n_11173), .Y(n_2408));
OR4X1 g64932(.A (n_1735), .B (g4616), .C (n_9019), .D (g4608), .Y(n_2406));
NAND3X1 g64956(.A (n_2403), .B (n_572), .C (g4057), .Y (n_3728));
NAND3X1 g64957(.A (n_2403), .B (g4064), .C (g4057), .Y (n_3726));
NAND3X1 g64959(.A (n_2403), .B (g4064), .C (n_571), .Y (n_3730));
NAND3X1 g64960(.A (n_1757), .B (g1472), .C (n_9698), .Y (n_2400));
INVX1 g64962(.A (n_2456), .Y (n_2630));
AOI21X1 g64983(.A0 (g_16456), .A1 (n_10557), .B0 (n_10560), .Y(n_2983));
XOR2X1 g64984(.A (n_3171), .B (g25219), .Y (n_2398));
XOR2X1 g64987(.A (n_2732), .B (n_2376), .Y (n_2397));
NAND2X1 g66444(.A (n_365), .B (n_9091), .Y (n_2849));
XOR2X1 g64991(.A (n_11157), .B (n_2729), .Y (n_2392));
AOI21X1 g64996(.A0 (n_10557), .A1 (g_18869), .B0 (n_10560), .Y(n_2670));
NAND4X1 g65022(.A (n_10906), .B (g4765), .C (n_8639), .D (n_8777), .Y(n_2391));
NAND4X1 g65023(.A (g5240), .B (n_10621), .C (g14597), .D (g25219), .Y(n_2389));
NAND4X1 g65026(.A (g6625), .B (n_3275), .C (g14749), .D (n_11184), .Y(n_2388));
NAND4X1 g65027(.A (g16744), .B (g16627), .C (g11388), .D (g13926), .Y(n_3062));
NAND4X1 g65028(.A (g16718), .B (g16603), .C (g_4050), .D (g13895), .Y(n_3065));
NOR2X1 g66441(.A (g4332), .B (n_9884), .Y (n_3213));
NAND4X1 g65033(.A (n_8676), .B (g4944), .C (n_10984), .D (n_10998),.Y (n_2387));
NAND4X1 g65035(.A (n_10905), .B (g4743), .C (n_8639), .D (n_8810), .Y(n_2385));
NAND4X1 g65037(.A (g5587), .B (n_7150), .C (g14635), .D (n_1023), .Y(n_2382));
NAND4X1 g65038(.A (n_8676), .B (g4933), .C (n_10185), .D (n_10984),.Y (n_10181));
NAND4X1 g65039(.A (g6279), .B (n_3277), .C (g14705), .D (n_11157), .Y(n_2379));
NAND4X1 g65040(.A (g5933), .B (n_10506), .C (g14673), .D (n_2376), .Y(n_2378));
OAI21X1 g65046(.A0 (g6167), .A1 (n_4324), .B0 (n_1776), .Y (n_2375));
MX2X1 g65072(.A (g_20614), .B (g_15758), .S0 (n_1491), .Y (n_2374));
XOR2X1 g65082(.A (n_1409), .B (n_650), .Y (n_2373));
OR2X1 g65240(.A (n_4329), .B (n_9772), .Y (n_2372));
OR2X1 g65242(.A (n_4327), .B (n_9772), .Y (n_2370));
OR2X1 g65244(.A (n_4320), .B (n_9772), .Y (n_2368));
OR2X1 g65247(.A (n_4314), .B (n_9772), .Y (n_2367));
OR2X1 g65250(.A (n_4322), .B (n_9772), .Y (n_2366));
OR2X1 g65251(.A (n_4324), .B (n_9772), .Y (n_2365));
OR2X1 g65270(.A (n_1493), .B (g5033), .Y (n_2364));
INVX1 g65282(.A (n_2640), .Y (n_2363));
INVX1 g65308(.A (n_2361), .Y (n_3073));
NAND2X1 g65332(.A (n_6705), .B (n_10687), .Y (n_2785));
OR2X1 g65347(.A (n_2008), .B (n_1729), .Y (n_2608));
NAND2X1 g65364(.A (g4477), .B (n_9836), .Y (n_2356));
NAND2X1 g65374(.A (n_1124), .B (n_9521), .Y (n_4939));
NAND4X1 g65385(.A (n_2443), .B (g5579), .C (g17813), .D (n_2208), .Y(n_2354));
NAND4X1 g65388(.A (n_2352), .B (g6271), .C (g17845), .D (n_11150), .Y(n_2353));
AND2X1 g65399(.A (n_2064), .B (n_1626), .Y (n_2351));
NAND3X1 g61946(.A (n_1995), .B (g_16456), .C (n_9311), .Y (n_2350));
NAND4X1 g65403(.A (n_2432), .B (g6617), .C (g17871), .D (n_11178), .Y(n_2349));
NOR2X1 g65409(.A (g16718), .B (n_2020), .Y (n_2348));
NOR2X1 g65413(.A (g16744), .B (n_2023), .Y (n_2347));
NAND2X1 g61950(.A (n_1644), .B (n_2345), .Y (n_2346));
NAND4X1 g65452(.A (n_10831), .B (g5196), .C (g13039), .D (g25219), .Y(n_2344));
NAND4X1 g65453(.A (n_2413), .B (g6235), .C (g13085), .D (n_11157), .Y(n_2343));
NAND4X1 g65454(.A (g6247), .B (n_3277), .C (g13085), .D (n_11150), .Y(n_2342));
NAND4X1 g65456(.A (g5224), .B (n_2339), .C (g17787), .D (g25219), .Y(n_2340));
NAND4X1 g65459(.A (g6609), .B (n_2600), .C (g17871), .D (n_11177), .Y(n_2338));
NAND4X1 g65460(.A (n_2439), .B (g5543), .C (g13049), .D (n_1023), .Y(n_2336));
NAND4X1 g65461(.A (g6597), .B (n_2600), .C (g17722), .D (n_11173), .Y(n_2334));
NAND4X1 g65462(.A (g5200), .B (n_2339), .C (g12238), .D (g25219), .Y(n_2332));
NAND4X1 g65474(.A (n_2597), .B (g5559), .C (g17604), .D (n_2208), .Y(n_2331));
NAND4X1 g65475(.A (g5555), .B (n_7150), .C (g13049), .D (n_2208), .Y(n_2329));
NAND4X1 g65478(.A (g5571), .B (n_2597), .C (g17813), .D (n_1023), .Y(n_2327));
NAND4X1 g65480(.A (g6251), .B (n_2325), .C (g17685), .D (n_11150), .Y(n_2326));
NAND4X1 g65482(.A (g6263), .B (n_2325), .C (g17845), .D (n_11157), .Y(n_2324));
NAND4X1 g65487(.A (g6593), .B (n_3275), .C (g13099), .D (n_11178), .Y(n_2323));
NAND4X1 g65488(.A (n_2435), .B (g6581), .C (g13099), .D (n_11184), .Y(n_2321));
INVX1 g65597(.A (g16659), .Y (n_2594));
INVX1 g65644(.A (n_3184), .Y (n_2320));
INVX1 g65688(.A (n_6395), .Y (n_2319));
NOR2X1 g65889(.A (n_10402), .B (n_9107), .Y (n_2316));
NAND2X1 g65896(.A (n_8809), .B (n_9351), .Y (n_2580));
INVX1 g65915(.A (n_3177), .Y (n_2577));
NAND2X1 g63196(.A (n_2312), .B (g4854), .Y (n_2925));
NOR2X1 g66376(.A (n_6324), .B (n_10078), .Y (n_2311));
XOR2X1 g66173(.A (n_8768), .B (n_8837), .Y (n_2310));
XOR2X1 g66182(.A (n_10196), .B (n_3849), .Y (n_2309));
NOR2X1 g66281(.A (n_6252), .B (n_10716), .Y (n_2308));
NAND2X1 g66286(.A (n_2306), .B (n_10078), .Y (n_2307));
INVX1 g66288(.A (n_2304), .Y (n_2305));
NOR2X1 g66291(.A (n_8799), .B (n_9193), .Y (n_2303));
NOR2X1 g66295(.A (g5352), .B (n_9107), .Y (n_2302));
NAND2X1 g66296(.A (g1361), .B (n_9628), .Y (n_2301));
NAND2X1 g66298(.A (g6505), .B (n_9599), .Y (n_2298));
NAND2X1 g66310(.A (n_1502), .B (n_9874), .Y (n_2562));
NAND2X1 g66317(.A (n_303), .B (n_9894), .Y (n_2847));
NOR2X1 g66321(.A (g_18308), .B (n_10078), .Y (n_2296));
NAND2X1 g66326(.A (n_2293), .B (n_10078), .Y (n_2294));
NOR2X1 g66327(.A (n_2290), .B (n_9129), .Y (n_2291));
NOR2X1 g66335(.A (g6044), .B (n_10078), .Y (n_2289));
NAND2X1 g66338(.A (g1373), .B (n_9599), .Y (n_2288));
NAND2X1 g66340(.A (g_19911), .B (n_9193), .Y (n_2286));
NAND2X1 g66341(.A (n_10499), .B (n_9353), .Y (n_2285));
NAND2X1 g66344(.A (g2629), .B (n_9775), .Y (n_2284));
NAND2X1 g66348(.A (g1379), .B (n_9353), .Y (n_2283));
NAND2X1 g66349(.A (n_2280), .B (n_9884), .Y (n_2281));
NAND2X1 g66351(.A (n_10119), .B (n_9300), .Y (n_2278));
NOR2X1 g66352(.A (g6390), .B (n_9371), .Y (n_2277));
NOR2X1 g66361(.A (g5029), .B (n_9672), .Y (n_2276));
NOR2X1 g66372(.A (g6736), .B (n_9903), .Y (n_2274));
NAND2X1 g66383(.A (g2070), .B (n_9884), .Y (n_2272));
NAND2X1 g66388(.A (n_383), .B (n_9894), .Y (n_2855));
NOR2X1 g66395(.A (n_6928), .B (n_9903), .Y (n_2271));
NOR2X1 g66396(.A (n_6057), .B (n_9129), .Y (n_2270));
NAND2X1 g66399(.A (g4388), .B (n_9884), .Y (n_2269));
NAND2X1 g66400(.A (n_261), .B (n_9894), .Y (n_2842));
NAND2X1 g66402(.A (n_1275), .B (n_9599), .Y (n_2268));
NAND2X1 g66403(.A (g1936), .B (n_9672), .Y (n_2266));
NOR2X1 g66404(.A (g_12922), .B (n_9129), .Y (n_2265));
NAND2X1 g66408(.A (n_388), .B (n_9883), .Y (n_2859));
NOR2X1 g66426(.A (g3698), .B (n_9903), .Y (n_2264));
NOR2X1 g66436(.A (n_10647), .B (n_9129), .Y (n_2263));
NOR2X1 g66466(.A (g_11293), .B (n_10782), .Y (n_2260));
NAND2X1 g66467(.A (n_2258), .B (n_9628), .Y (n_2259));
NAND2X1 g66468(.A (g_19233), .B (n_9599), .Y (n_2256));
NAND2X1 g66474(.A (g_21576), .B (n_10952), .Y (n_2255));
NAND2X1 g66476(.A (n_933), .B (n_10078), .Y (n_2254));
NOR2X1 g66477(.A (n_2252), .B (n_10782), .Y (n_2253));
NOR2X1 g66496(.A (g_15879), .B (n_9129), .Y (n_2250));
NOR2X1 g66514(.A (g_16311), .B (n_10782), .Y (n_2249));
NOR2X1 g66518(.A (g_16464), .B (n_9129), .Y (n_2248));
NAND2X1 g66524(.A (g2361), .B (n_9836), .Y (n_2247));
NOR2X1 g66534(.A (n_8793), .B (n_9129), .Y (n_2246));
NAND2X1 g66537(.A (n_2244), .B (n_9976), .Y (n_2245));
NAND2X1 g66539(.A (n_3383), .B (n_9193), .Y (n_2243));
NAND2X1 g66542(.A (n_4139), .B (n_9371), .Y (n_2242));
NOR2X1 g66546(.A (g5698), .B (n_10078), .Y (n_2241));
NOR2X1 g66554(.A (g4049), .B (n_10376), .Y (n_2239));
NOR2X1 g66556(.A (g3347), .B (n_9903), .Y (n_2237));
NAND2X1 g66562(.A (n_370), .B (n_9894), .Y (n_2853));
NAND2X1 g66574(.A (g4854), .B (n_9884), .Y (n_2234));
NAND2X1 g66581(.A (n_215), .B (n_9139), .Y (n_2857));
NOR2X1 g66594(.A (n_388), .B (n_9107), .Y (n_2233));
AND2X1 g66609(.A (g2823), .B (n_9091), .Y (n_2231));
NOR2X1 g66610(.A (g2518), .B (n_9693), .Y (n_2230));
NOR2X1 g66612(.A (g2384), .B (n_9903), .Y (n_2229));
AND2X1 g66616(.A (g5499), .B (n_9209), .Y (n_2228));
AND2X1 g66640(.A (g3143), .B (n_9521), .Y (n_2227));
NOR2X1 g66650(.A (n_303), .B (n_9903), .Y (n_2225));
NAND2X1 g66662(.A (n_2224), .B (n_9139), .Y (n_2838));
NOR2X1 g66671(.A (n_215), .B (n_9775), .Y (n_2223));
NOR2X1 g66678(.A (n_10307), .B (n_10078), .Y (n_2221));
NOR2X1 g66679(.A (n_330), .B (n_9884), .Y (n_2219));
AND2X1 g66683(.A (g5845), .B (n_9521), .Y (n_2218));
NOR2X1 g66685(.A (g1467), .B (n_9353), .Y (n_2216));
AND2X1 g66689(.A (n_10813), .B (n_9521), .Y (n_2215));
NAND2X1 g66700(.A (n_11171), .B (n_9883), .Y (n_2835));
NOR2X1 g66706(.A (g1959), .B (n_9693), .Y (n_2212));
AND2X1 g66719(.A (g3845), .B (n_9521), .Y (n_2211));
NOR2X1 g66726(.A (g1454), .B (n_9107), .Y (n_2210));
NAND4X1 g64872(.A (n_2439), .B (g5595), .C (g14635), .D (n_2208), .Y(n_2209));
AND2X1 g66776(.A (g3494), .B (n_9139), .Y (n_2207));
AND2X1 g66790(.A (g6191), .B (n_9311), .Y (n_2206));
NOR2X1 g66812(.A (g1437), .B (n_9353), .Y (n_2205));
NOR2X1 g66859(.A (n_6527), .B (n_9599), .Y (n_2496));
NAND2X1 g66882(.A (n_5402), .B (n_9139), .Y (n_2828));
AND2X1 g66888(.A (g6537), .B (n_9521), .Y (n_2204));
NOR2X1 g66900(.A (n_370), .B (n_10078), .Y (n_2203));
OR2X1 g61528(.A (n_2192), .B (n_129), .Y (n_2790));
XOR2X1 g63640(.A (g20557), .B (n_1581), .Y (n_2182));
XOR2X1 g63643(.A (g4273), .B (n_1583), .Y (n_2181));
NAND2X1 g61201(.A (n_1277), .B (n_11073), .Y (n_2180));
NAND2X1 g61202(.A (n_11073), .B (n_2177), .Y (n_2178));
NAND2X1 g61204(.A (n_11073), .B (n_6782), .Y (n_2176));
INVX1 g61207(.A (n_11041), .Y (n_2830));
INVX1 g62287(.A (n_1883), .Y (n_2174));
INVX1 g62289(.A (n_1882), .Y (n_2173));
INVX1 g61218(.A (n_2592), .Y (n_2172));
AOI21X1 g64681(.A0 (n_1546), .A1 (n_1312), .B0 (n_2111), .Y (g31521));
NOR2X1 g66856(.A (g1825), .B (n_10376), .Y (n_2168));
OAI21X1 g64146(.A0 (n_692), .A1 (n_11162), .B0 (n_1860), .Y (n_2167));
OR2X1 g64147(.A (n_2165), .B (n_221), .Y (n_2166));
NAND2X1 g64258(.A (n_1700), .B (n_1847), .Y (n_2163));
OAI21X1 g62657(.A0 (n_1840), .A1 (g4664), .B0 (n_2867), .Y (n_2161));
MX2X1 g64424(.A (g_21806), .B (g_20837), .S0 (n_6460), .Y (n_2160));
MX2X1 g64431(.A (g_22379), .B (g_21806), .S0 (n_6460), .Y (n_2159));
MX2X1 g64434(.A (g_21576), .B (g_22379), .S0 (n_6460), .Y (n_2157));
MX2X1 g64457(.A (g_6131), .B (g_19241), .S0 (n_6460), .Y (n_2156));
MX2X1 g64459(.A (n_5663), .B (g_6131), .S0 (n_6460), .Y (n_2155));
AND2X1 g64512(.A (n_1817), .B (n_6464), .Y (n_3174));
NAND3X1 g64555(.A (n_2153), .B (n_2457), .C (n_2747), .Y (n_2154));
NOR2X1 g64605(.A (n_2106), .B (n_8637), .Y (n_2483));
NAND4X1 g64633(.A (n_335), .B (n_17), .C (n_943), .D (n_353), .Y(n_2152));
AOI21X1 g64646(.A0 (n_1013), .A1 (n_2150), .B0 (n_1559), .Y (n_2151));
NAND4X1 g64693(.A (n_2133), .B (n_2439), .C (g14694), .D (g5583), .Y(n_2149));
NAND4X1 g64696(.A (n_2119), .B (n_2435), .C (g14828), .D (g6621), .Y(n_2148));
NAND4X1 g64700(.A (n_10877), .B (g3586), .C (g16744), .D (n_6973), .Y(n_2146));
NAND4X1 g64717(.A (n_2143), .B (g5244), .C (g17674), .D (g25114), .Y(n_2145));
NAND4X1 g64718(.A (n_2143), .B (g5228), .C (g14662), .D (n_10621), .Y(n_2144));
NAND4X1 g64724(.A (n_2131), .B (n_2352), .C (g17760), .D (g6283), .Y(n_2141));
NAND4X1 g64725(.A (n_10879), .B (g3594), .C (g16744), .D (n_11128),.Y (n_2140));
NAND4X1 g64727(.A (n_10877), .B (g3570), .C (g13926), .D (n_4682), .Y(n_2138));
NAND4X1 g64730(.A (n_2447), .B (g3921), .C (g13966), .D (n_6787), .Y(n_2137));
NAND4X1 g64744(.A (n_2133), .B (g5615), .C (g17580), .D (n_7150), .Y(n_2135));
NAND4X1 g64746(.A (n_2133), .B (g5599), .C (g17711), .D (n_2597), .Y(n_2134));
NAND4X1 g64752(.A (n_2131), .B (g6267), .C (g14779), .D (n_3277), .Y(n_2132));
NAND4X1 g64753(.A (n_2131), .B (n_2413), .C (g17649), .D (g6299), .Y(n_2130));
NAND4X1 g64754(.A (n_2127), .B (n_10809), .C (g17607), .D (g5953), .Y(n_2129));
NAND4X1 g64755(.A (n_2127), .B (g5921), .C (g14738), .D (n_10506), .Y(n_2128));
NAND4X1 g64756(.A (n_2127), .B (n_10622), .C (g17739), .D (g5937), .Y(n_2126));
NAND4X1 g64764(.A (n_2119), .B (g6653), .C (g17688), .D (n_3275), .Y(n_2122));
NAND4X1 g64765(.A (n_2143), .B (n_10831), .C (g17519), .D (g5260), .Y(n_2121));
NAND4X1 g64767(.A (n_2119), .B (g6637), .C (g17778), .D (n_2600), .Y(n_2120));
NOR2X1 g65294(.A (g26801), .B (n_9856), .Y (n_2973));
NOR2X1 g64875(.A (n_2458), .B (n_10725), .Y (n_2118));
AND2X1 g64877(.A (n_3021), .B (n_2115), .Y (n_3047));
AND2X1 g64884(.A (n_2113), .B (n_2115), .Y (n_2116));
AND2X1 g64886(.A (n_3021), .B (n_2113), .Y (n_2114));
OR2X1 g64894(.A (n_1737), .B (n_2111), .Y (n_3897));
NOR2X1 g64895(.A (n_1552), .B (g8788), .Y (n_2110));
NOR2X1 g64902(.A (n_10551), .B (n_10552), .Y (n_2107));
INVX1 g64922(.A (n_2106), .Y (n_2410));
NAND4X1 g64955(.A (n_1544), .B (g4087), .C (g4076), .D (g4098), .Y(n_2103));
AND2X1 g64963(.A (n_1555), .B (n_2113), .Y (n_2456));
AOI21X1 g64981(.A0 (n_397), .A1 (n_10499), .B0 (n_10725), .Y(n_2654));
INVX1 g65012(.A (n_2100), .Y (n_2101));
XOR2X1 g65042(.A (g1677), .B (n_1248), .Y (n_2099));
OAI21X1 g65043(.A0 (g5475), .A1 (n_4329), .B0 (n_1535), .Y (n_2098));
OAI21X1 g65044(.A0 (g5821), .A1 (n_4327), .B0 (n_1545), .Y (n_2097));
XOR2X1 g65045(.A (g1811), .B (n_1237), .Y (n_2096));
OAI21X1 g65048(.A0 (g6513), .A1 (n_4322), .B0 (n_1553), .Y (n_2095));
XOR2X1 g65049(.A (g1945), .B (n_1231), .Y (n_2094));
OAI21X1 g65053(.A0 (g3821), .A1 (n_4314), .B0 (n_1547), .Y (n_2093));
OAI21X1 g65054(.A0 (g3119), .A1 (n_4316), .B0 (n_1539), .Y (n_2092));
OAI21X1 g65055(.A0 (g3470), .A1 (n_4320), .B0 (n_1551), .Y (n_2091));
XOR2X1 g65056(.A (n_7260), .B (n_6582), .Y (n_2090));
XOR2X1 g65057(.A (g2370), .B (n_1161), .Y (n_2089));
XOR2X1 g65059(.A (g2504), .B (n_1139), .Y (n_2088));
XOR2X1 g65060(.A (g5128), .B (g26801), .Y (n_2087));
MX2X1 g65061(.A (n_2936), .B (g6159), .S0 (n_4324), .Y (n_2086));
MX2X1 g65066(.A (n_2704), .B (n_2084), .S0 (n_4324), .Y (n_2085));
MX2X1 g65077(.A (n_1732), .B (n_6958), .S0 (n_1731), .Y (n_2083));
XOR2X1 g65083(.A (n_10550), .B (n_10568), .Y (n_2082));
XOR2X1 g65089(.A (g2638), .B (n_1014), .Y (n_2081));
XOR2X1 g65093(.A (g2079), .B (n_1304), .Y (n_2080));
XOR2X1 g65095(.A (g2236), .B (n_1168), .Y (n_2079));
NOR2X1 g65235(.A (n_389), .B (n_2077), .Y (n_2078));
NOR2X1 g65239(.A (n_202), .B (n_10475), .Y (n_2072));
NAND2X1 g65256(.A (n_1662), .B (g5033), .Y (n_2070));
AND2X1 g65261(.A (n_2067), .B (n_8694), .Y (n_2069));
AND2X1 g65263(.A (n_2067), .B (n_8777), .Y (n_2068));
NOR2X1 g66777(.A (n_708), .B (n_10078), .Y (n_3857));
OR2X1 g65283(.A (n_11027), .B (n_1652), .Y (n_2640));
AND2X1 g65285(.A (n_10184), .B (n_2064), .Y (n_2065));
NAND2X1 g65299(.A (n_2062), .B (g1306), .Y (n_2063));
INVX1 g65309(.A (n_2061), .Y (n_2361));
OR2X1 g61396(.A (n_2060), .B (n_26), .Y (n_2671));
NAND2X1 g65338(.A (n_10200), .B (n_9651), .Y (n_2784));
INVX1 g65359(.A (n_2056), .Y (n_2057));
NOR2X1 g65367(.A (n_1462), .B (n_7260), .Y (n_2055));
INVX1 g65368(.A (n_2053), .Y (n_2054));
NOR2X1 g65390(.A (n_10527), .B (g_8896), .Y (n_2639));
NAND2X1 g65394(.A (n_8906), .B (n_2067), .Y (n_2051));
AND2X1 g65395(.A (n_2067), .B (n_8809), .Y (n_2049));
NAND2X1 g65400(.A (n_10205), .B (n_2064), .Y (n_2048));
AND2X1 g65401(.A (n_2064), .B (n_10296), .Y (n_2046));
AND2X1 g65404(.A (n_2045), .B (n_2044), .Y (n_3984));
INVX1 g65417(.A (n_2427), .Y (n_2043));
INVX1 g65427(.A (n_10765), .Y (n_2042));
NAND4X1 g65449(.A (g5208), .B (n_10621), .C (g13039), .D (n_1695), .Y(n_2038));
AOI22X1 g65464(.A0 (n_10206), .A1 (g4888), .B0 (g4955), .B1(n_10214), .Y (n_11192));
AOI22X1 g65466(.A0 (g4917), .A1 (n_10214), .B0 (g4912), .B1(n_10206), .Y (n_2034));
MX2X1 g61964(.A (n_2429), .B (g_19172), .S0 (n_2878), .Y (n_2032));
NAND4X1 g65476(.A (g5212), .B (n_2339), .C (g17577), .D (n_1695), .Y(n_2031));
NAND4X1 g65479(.A (g6239), .B (n_2325), .C (g12422), .D (n_11157), .Y(n_2030));
NAND4X1 g65484(.A (g5893), .B (n_11101), .C (g12350), .D (n_546), .Y(n_2029));
NAND4X1 g65485(.A (g5917), .B (n_11101), .C (g17819), .D (n_546), .Y(n_2027));
NAND4X1 g65486(.A (n_10808), .B (g5889), .C (g13068), .D (n_546), .Y(n_2025));
AOI21X1 g65504(.A0 (n_8917), .A1 (g4049), .B0 (n_1479), .Y (n_2024));
NOR2X1 g65689(.A (n_2019), .B (n_4878), .Y (n_6395));
AND2X1 g65727(.A (n_2600), .B (n_9091), .Y (n_2018));
NAND2X1 g65645(.A (n_2001), .B (n_2017), .Y (n_3184));
NAND2X1 g65794(.A (n_11126), .B (n_10687), .Y (n_2016));
AND2X1 g65796(.A (n_2325), .B (n_10687), .Y (n_2015));
NAND2X1 g65798(.A (n_8572), .B (n_9311), .Y (n_2014));
DFFSRX1 g1582_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7946), .Q (g8475), .QN ());
AND2X1 g65838(.A (n_11101), .B (n_9521), .Y (n_2011));
NAND2X1 g65843(.A (n_6808), .B (n_10687), .Y (n_2009));
INVX1 g65847(.A (n_2008), .Y (n_4632));
AND2X1 g65865(.A (n_2597), .B (n_9750), .Y (n_2007));
OR2X1 g65866(.A (n_1628), .B (n_2005), .Y (n_2006));
NOR2X1 g65878(.A (g4927), .B (n_1625), .Y (n_2004));
INVX1 g62034(.A (n_2002), .Y (n_2003));
NAND3X1 g65970(.A (n_2001), .B (n_488), .C (n_10524), .Y (n_3718));
NAND2X1 g66747(.A (n_2556), .B (n_9501), .Y (n_2000));
MX2X1 g66125(.A (g1521), .B (g1532), .S0 (n_3849), .Y (n_1997));
INVX1 g62062(.A (n_1995), .Y (n_1996));
INVX1 g62068(.A (n_1993), .Y (n_1994));
MX2X1 g66104(.A (g1178), .B (g1189), .S0 (n_8837), .Y (n_1992));
MX2X1 g66150(.A (g_20614), .B (g1178), .S0 (n_8837), .Y (n_1991));
OAI21X1 g63528(.A0 (n_1307), .A1 (g4659), .B0 (n_1329), .Y (n_1989));
NOR2X1 g66289(.A (n_1627), .B (n_9884), .Y (n_2304));
NAND2X1 g66324(.A (n_330), .B (n_9521), .Y (n_2578));
OR2X1 g66360(.A (g4467), .B (n_9628), .Y (n_2862));
INVX1 g66363(.A (n_1985), .Y (n_1986));
OR2X1 g66527(.A (g1306), .B (n_10078), .Y (n_2480));
NAND2X1 g66583(.A (n_8588), .B (n_9351), .Y (n_2661));
NAND2X1 g66585(.A (g1542), .B (n_9521), .Y (n_1982));
NAND2X1 g66589(.A (n_11157), .B (n_9139), .Y (n_2606));
INVX1 g66592(.A (n_5453), .Y (n_1980));
NAND2X1 g66623(.A (g1199), .B (n_9894), .Y (n_1979));
NAND2X1 g66628(.A (n_10894), .B (n_9351), .Y (n_2668));
NOR2X1 g66677(.A (n_10503), .B (n_9526), .Y (n_2657));
NAND2X1 g66680(.A (n_2376), .B (n_9883), .Y (n_2612));
NAND2X1 g66705(.A (n_2280), .B (n_9501), .Y (n_1977));
NAND2X1 g66713(.A (g_18739), .B (n_9139), .Y (n_1976));
OR2X1 g65414(.A (n_1426), .B (n_8809), .Y (n_1975));
NOR2X1 g66749(.A (n_6782), .B (n_9856), .Y (n_3372));
NOR2X1 g66773(.A (g4332), .B (n_662), .Y (n_1972));
NAND2X1 g66785(.A (g4608), .B (n_9627), .Y (n_1971));
NAND2X1 g66826(.A (n_2529), .B (n_9521), .Y (n_1969));
AND2X1 g66829(.A (g2827), .B (n_10687), .Y (n_1968));
OR2X1 g64846(.A (n_10520), .B (n_2017), .Y (n_1887));
AOI21X1 g62278(.A0 (n_11029), .A1 (g3343), .B0 (n_1473), .Y (n_1885));
AOI21X1 g62279(.A0 (n_10576), .A1 (g3694), .B0 (n_1474), .Y (n_1884));
INVX1 g68049(.A (n_2224), .Y (n_2734));
AOI21X1 g62288(.A0 (n_10941), .A1 (g3347), .B0 (n_1311), .Y (n_1883));
AOI21X1 g62290(.A0 (n_6972), .A1 (g3698), .B0 (n_1310), .Y (n_1882));
AND2X1 g61219(.A (n_1443), .B (n_10329), .Y (n_2592));
DFFSRX1 g1239_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7916), .Q (g8416), .QN ());
INVX1 g64144(.A (n_2312), .Y (n_1875));
MX2X1 g61296(.A (n_460), .B (g1521), .S0 (n_3849), .Y (n_1869));
NAND2X1 g66478(.A (g_5342), .B (n_9091), .Y (n_1865));
NAND4X1 g64525(.A (n_235), .B (n_157), .C (n_958), .D (n_194), .Y(n_1863));
NAND4X1 g64594(.A (n_425), .B (n_29), .C (n_950), .D (n_428), .Y(n_1862));
NAND4X1 g64619(.A (n_340), .B (n_5), .C (n_947), .D (n_248), .Y(n_1861));
AOI22X1 g64680(.A0 (n_694), .A1 (g_21720), .B0 (n_693), .B1(g_19233), .Y (n_1860));
NAND4X1 g64692(.A (n_1854), .B (n_10833), .C (g14662), .D (g5236), .Y(n_1859));
NAND4X1 g64694(.A (n_1848), .B (n_2413), .C (g14779), .D (g6275), .Y(n_1858));
NAND4X1 g64695(.A (n_1845), .B (n_10809), .C (g14738), .D (g5929), .Y(n_1857));
NAND4X1 g64712(.A (n_1854), .B (g5252), .C (g17674), .D (n_2339), .Y(n_1855));
NAND4X1 g64713(.A (n_1854), .B (g5268), .C (g17519), .D (n_10621), .Y(n_11194));
NAND4X1 g64715(.A (n_8548), .B (g3227), .C (g13895), .D (n_11029), .Y(n_6948));
NAND4X1 g64733(.A (n_6806), .B (g3929), .C (g13966), .D (n_4988), .Y(n_1851));
NAND4X1 g64738(.A (n_10879), .B (g3578), .C (g13926), .D (n_10576),.Y (n_1850));
NAND4X1 g64750(.A (n_1848), .B (g6291), .C (g17760), .D (n_2325), .Y(n_1849));
NAND4X1 g64751(.A (n_1848), .B (g6307), .C (g17649), .D (n_3277), .Y(n_1847));
NAND4X1 g64757(.A (n_1845), .B (g5945), .C (g17739), .D (n_11101), .Y(n_1846));
NAND4X1 g64758(.A (n_1845), .B (g5961), .C (g17607), .D (n_10508), .Y(n_1844));
MX2X1 g65074(.A (n_2923), .B (g3813), .S0 (n_4314), .Y (n_1843));
XOR2X1 g64775(.A (n_307), .B (n_474), .Y (n_1842));
NAND2X1 g62798(.A (n_1840), .B (g4664), .Y (n_2867));
XOR2X1 g64776(.A (g4269), .B (n_1582), .Y (n_1839));
OAI22X1 g64777(.A0 (n_821), .A1 (n_1831), .B0 (n_747), .B1 (g4593),.Y (n_1838));
NAND3X1 g64889(.A (n_991), .B (n_6762), .C (g7916), .Y (n_1833));
AND2X1 g64900(.A (n_1096), .B (n_1831), .Y (n_1832));
INVX1 g64904(.A (n_10597), .Y (n_1830));
OR2X1 g64923(.A (n_10907), .B (g4688), .Y (n_2106));
OR2X1 g64925(.A (n_1016), .B (n_1826), .Y (n_1827));
AOI22X1 g65465(.A0 (g4933), .A1 (n_10185), .B0 (g4944), .B1(n_10998), .Y (n_11193));
AOI21X1 g64994(.A0 (g_13758), .A1 (n_3550), .B0 (n_1291), .Y(n_1822));
OAI21X1 g65007(.A0 (n_1820), .A1 (g8839), .B0 (n_1278), .Y (n_1821));
XOR2X1 g65013(.A (g4527), .B (n_1562), .Y (n_2100));
AOI21X1 g65014(.A0 (n_1818), .A1 (g34036), .B0 (n_994), .Y (n_1819));
MX2X1 g65020(.A (n_6501), .B (n_924), .S0 (n_11051), .Y (n_1817));
MX2X1 g65062(.A (n_2718), .B (n_1813), .S0 (n_1812), .Y (n_1814));
MX2X1 g65063(.A (n_3011), .B (n_1810), .S0 (n_4329), .Y (n_1811));
MX2X1 g65064(.A (n_2940), .B (g5813), .S0 (n_4327), .Y (n_1809));
MX2X1 g65065(.A (n_2684), .B (n_1807), .S0 (n_4327), .Y (n_1808));
MX2X1 g65067(.A (n_2686), .B (n_1805), .S0 (n_4316), .Y (n_1806));
MX2X1 g65068(.A (n_2005), .B (g1489), .S0 (n_4617), .Y (n_1804));
MX2X1 g65069(.A (n_2930), .B (g6505), .S0 (n_4322), .Y (n_1803));
MX2X1 g65070(.A (n_3253), .B (g3111), .S0 (n_4316), .Y (n_1802));
MX2X1 g65071(.A (n_2928), .B (g3462), .S0 (n_4320), .Y (n_1801));
MX2X1 g65073(.A (n_2699), .B (n_1799), .S0 (n_4320), .Y (n_1800));
MX2X1 g65075(.A (n_2943), .B (g5467), .S0 (n_4329), .Y (n_1798));
MX2X1 g65076(.A (n_2692), .B (n_1796), .S0 (n_4314), .Y (n_1797));
MX2X1 g65078(.A (n_3007), .B (n_1794), .S0 (n_4322), .Y (n_1795));
MX2X1 g65079(.A (g1442), .B (n_2005), .S0 (n_4617), .Y (n_1793));
MX2X1 g65080(.A (g5156), .B (g5120), .S0 (n_1812), .Y (n_1792));
AOI21X1 g65085(.A0 (n_720), .A1 (n_564), .B0 (n_1251), .Y (n_1791));
DFFSRX1 g5335_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14597), .Q (g17639), .QN ());
DFFSRX1 g5681_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14635), .Q (g17678), .QN ());
DFFSRX1 g6027_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14673), .Q (g17715), .QN ());
DFFSRX1 g6373_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14705), .Q (g17743), .QN ());
DFFSRX1 g6719_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14749), .Q (g17764), .QN ());
NOR2X1 g65232(.A (n_3030), .B (n_1250), .Y (n_1789));
NOR2X1 g65233(.A (n_1266), .B (n_1631), .Y (n_1788));
NOR2X1 g65234(.A (n_1405), .B (g_15380), .Y (n_1787));
AND2X1 g65246(.A (n_10984), .B (n_8676), .Y (n_1786));
AND2X1 g65249(.A (n_8639), .B (n_10905), .Y (n_1785));
NAND2X1 g65252(.A (n_6582), .B (n_7260), .Y (n_2165));
NOR2X1 g65253(.A (n_6578), .B (n_1220), .Y (n_1783));
OR2X1 g65255(.A (n_7010), .B (g5033), .Y (n_6970));
NAND2X1 g65257(.A (n_1765), .B (n_1391), .Y (n_1780));
NAND2X1 g65258(.A (n_1770), .B (n_1471), .Y (n_1779));
NAND2X1 g65259(.A (n_1772), .B (n_1777), .Y (n_1778));
NAND2X1 g65262(.A (g6167), .B (n_4324), .Y (n_1776));
NAND2X1 g65268(.A (n_1763), .B (n_1480), .Y (n_1775));
NAND2X1 g65274(.A (n_1772), .B (n_1476), .Y (n_1773));
NAND2X1 g65284(.A (n_1770), .B (n_1377), .Y (n_1771));
NAND2X1 g65286(.A (n_1767), .B (n_1584), .Y (n_1769));
NAND2X1 g65287(.A (n_1767), .B (n_1370), .Y (n_1768));
NAND2X1 g65290(.A (n_1765), .B (n_1445), .Y (n_1766));
NAND2X1 g65291(.A (n_1763), .B (n_1762), .Y (n_1764));
NAND2X1 g65295(.A (n_1772), .B (n_973), .Y (n_1761));
NAND2X1 g65300(.A (n_1767), .B (n_1758), .Y (n_1759));
INVX1 g65302(.A (n_1756), .Y (n_1757));
NAND2X1 g65304(.A (n_1727), .B (n_1382), .Y (n_1755));
OR2X1 g65310(.A (n_10983), .B (g4878), .Y (n_2061));
NAND2X1 g65314(.A (n_1752), .B (n_1450), .Y (n_1754));
NAND2X1 g65316(.A (n_1752), .B (n_1751), .Y (n_1753));
NAND2X1 g65317(.A (n_1752), .B (n_1367), .Y (n_1750));
NAND2X1 g65319(.A (n_1752), .B (n_1206), .Y (n_1749));
NAND2X1 g65322(.A (n_1767), .B (n_1242), .Y (n_1748));
AND2X1 g65325(.A (n_10214), .B (n_8676), .Y (n_1747));
NAND2X1 g65330(.A (n_1744), .B (n_1440), .Y (n_1746));
NAND2X1 g65331(.A (n_1744), .B (n_1743), .Y (n_1745));
NAND2X1 g65334(.A (n_1744), .B (n_1364), .Y (n_1741));
NAND2X1 g65335(.A (n_1744), .B (n_1184), .Y (n_1740));
NAND2X1 g65341(.A (n_1763), .B (n_970), .Y (n_1738));
INVX1 g65342(.A (n_1737), .Y (n_2403));
INVX1 g65344(.A (n_2677), .Y (n_1736));
NAND2X1 g65357(.A (n_918), .B (n_10949), .Y (n_2449));
NAND3X1 g65361(.A (n_1219), .B (n_7260), .C (n_1734), .Y (n_1735));
NOR2X1 g65362(.A (n_1732), .B (n_1731), .Y (n_1733));
NAND2X1 g65363(.A (n_1765), .B (n_590), .Y (n_1730));
NOR2X1 g65369(.A (n_1729), .B (n_1238), .Y (n_2053));
NAND2X1 g65376(.A (n_1727), .B (n_1245), .Y (n_1728));
NAND2X1 g65377(.A (n_1727), .B (n_1725), .Y (n_1726));
NAND2X1 g65378(.A (n_1770), .B (n_1723), .Y (n_1724));
NAND2X1 g65382(.A (n_1727), .B (n_1455), .Y (n_1722));
NAND2X1 g65384(.A (n_1770), .B (n_1264), .Y (n_1721));
NAND2X1 g65387(.A (n_1765), .B (n_1718), .Y (n_1719));
NAND4X1 g65392(.A (n_10623), .B (g5925), .C (g17819), .D (n_423), .Y(n_1717));
NAND2X1 g65398(.A (n_1772), .B (n_1411), .Y (n_1716));
AOI22X1 g65408(.A0 (n_790), .A1 (n_1714), .B0 (n_1713), .B1 (n_808),.Y (n_1715));
AOI22X1 g65410(.A0 (n_805), .A1 (n_1711), .B0 (n_1710), .B1 (n_798),.Y (n_1712));
NAND3X1 g65411(.A (n_10827), .B (n_746), .C (n_8796), .Y (n_1709));
AOI22X1 g65415(.A0 (n_697), .A1 (n_1706), .B0 (n_1705), .B1 (n_778),.Y (n_1707));
AOI22X1 g65421(.A0 (n_707), .A1 (n_1703), .B0 (n_1702), .B1 (n_793),.Y (n_1704));
NAND3X1 g65423(.A (n_2443), .B (n_1484), .C (g5619), .Y (n_1701));
NAND3X1 g65424(.A (n_2352), .B (n_1457), .C (g6311), .Y (n_1700));
NAND3X1 g65425(.A (n_10622), .B (n_1458), .C (g5965), .Y (n_1699));
NAND3X1 g65426(.A (n_2432), .B (n_1461), .C (g6657), .Y (n_1698));
NAND4X1 g65439(.A (g5232), .B (n_1695), .C (g17787), .D (g25114), .Y(n_1696));
NAND4X1 g65447(.A (g5905), .B (n_11101), .C (g17646), .D (n_423), .Y(n_1694));
NAND4X1 g65450(.A (g3542), .B (n_10895), .C (g11388), .D (n_11128),.Y (n_1691));
AOI22X1 g65455(.A0 (n_1062), .A1 (n_1688), .B0 (n_1687), .B1 (n_648),.Y (n_1689));
NAND4X1 g65457(.A (g3893), .B (n_5402), .C (g11418), .D (n_6808), .Y(n_1686));
AOI22X1 g65467(.A0 (g4907), .A1 (n_10185), .B0 (g4922), .B1(n_10998), .Y (n_1682));
AOI22X1 g65468(.A0 (g4743), .A1 (n_8810), .B0 (g4754), .B1 (n_8693),.Y (n_1681));
AOI22X1 g65469(.A0 (g4722), .A1 (n_10227), .B0 (g4727), .B1 (n_8778),.Y (n_1680));
AOI22X1 g65470(.A0 (n_1059), .A1 (n_1677), .B0 (n_1676), .B1 (n_591),.Y (n_1678));
AOI22X1 g65471(.A0 (g4717), .A1 (n_8810), .B0 (g4732), .B1 (n_8693),.Y (n_1675));
AOI22X1 g65472(.A0 (n_10227), .A1 (g4698), .B0 (g4765), .B1 (n_8778),.Y (n_1674));
AOI22X1 g65481(.A0 (n_1064), .A1 (n_1671), .B0 (n_1670), .B1 (n_486),.Y (n_1672));
NAND4X1 g65483(.A (g5901), .B (n_10506), .C (g13068), .D (n_423), .Y(n_1669));
INVX1 g65508(.A (n_2119), .Y (n_2433));
AOI22X1 g65448(.A0 (n_1667), .A1 (n_1666), .B0 (n_1665), .B1 (n_562),.Y (n_1668));
INVX1 g65592(.A (g16627), .Y (n_2023));
INVX1 g65610(.A (g16603), .Y (n_2020));
NAND3X1 g65707(.A (n_11113), .B (n_1352), .C (n_2017), .Y (n_1658));
OR2X1 g65784(.A (g4417), .B (n_5378), .Y (n_1657));
NAND2X1 g65848(.A (n_978), .B (g13272), .Y (n_2008));
INVX1 g65871(.A (n_1655), .Y (n_1656));
CLKBUFX1 g65917(.A (n_1652), .Y (n_3177));
NAND2X1 g65948(.A (n_817), .B (n_822), .Y (n_1650));
NAND2X1 g65961(.A (n_983), .B (n_795), .Y (n_1649));
NOR2X1 g62035(.A (n_2878), .B (n_799), .Y (n_2002));
INVX1 g62040(.A (n_1646), .Y (n_1647));
OR2X1 g62043(.A (n_2878), .B (g_19172), .Y (n_1645));
NAND2X1 g62044(.A (n_2878), .B (n_2429), .Y (n_1644));
OAI21X1 g66013(.A0 (g17604), .A1 (g13049), .B0 (n_1054), .Y (n_1643));
OAI21X1 g66015(.A0 (g17577), .A1 (g13039), .B0 (n_1094), .Y (n_1642));
OAI21X1 g66024(.A0 (g17685), .A1 (g13085), .B0 (n_1046), .Y (n_1641));
OAI21X1 g66042(.A0 (g17722), .A1 (g13099), .B0 (n_1021), .Y (n_1640));
NAND2X1 g62063(.A (n_4761), .B (n_1599), .Y (n_1995));
DFFSRX1 g3969_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16775), .Q (g16659), .QN ());
AND2X1 g65418(.A (n_1188), .B (n_1636), .Y (n_2427));
OR2X1 g66328(.A (g5084), .B (n_9836), .Y (n_5514));
OR2X1 g66364(.A (n_10123), .B (n_10376), .Y (n_1985));
OR2X1 g66462(.A (g_15758), .B (n_9371), .Y (n_2481));
NAND2X1 g66498(.A (n_35), .B (n_11055), .Y (n_1633));
NAND3X1 g64878(.A (n_1554), .B (n_1631), .C (n_1630), .Y (n_1632));
NOR2X1 g66593(.A (n_596), .B (n_9884), .Y (n_5453));
INVX1 g66595(.A (n_1628), .Y (n_1629));
NAND2X1 g66626(.A (n_1627), .B (n_9311), .Y (n_3192));
INVX1 g66631(.A (n_1625), .Y (n_1626));
NAND2X1 g65405(.A (n_1763), .B (n_1402), .Y (n_1605));
OAI21X1 g61588(.A0 (n_705), .A1 (g_15287), .B0 (g12919), .Y (n_2192));
NAND2X1 g62069(.A (n_4764), .B (n_1599), .Y (n_1993));
AND2X1 g63895(.A (n_2938), .B (n_1328), .Y (n_1597));
AND2X1 g64145(.A (n_1826), .B (g4849), .Y (n_2312));
NAND2X1 g64243(.A (n_1300), .B (n_1271), .Y (n_1592));
OR4X1 g65365(.A (g1333), .B (g19357), .C (g13272), .D (n_568), .Y(n_1591));
XOR2X1 g64779(.A (g5097), .B (n_1580), .Y (n_1590));
NOR2X1 g65360(.A (n_1729), .B (n_1422), .Y (n_2056));
CLKBUFX1 g68050(.A (n_1023), .Y (n_2224));
NAND3X1 g64593(.A (n_11217), .B (g3558), .C (n_6973), .Y (n_1587));
NAND3X1 g64628(.A (g3207), .B (n_801), .C (n_10941), .Y (n_1586));
NOR2X1 g65303(.A (n_1252), .B (n_1729), .Y (n_1756));
NAND2X1 g65699(.A (n_1243), .B (n_1584), .Y (n_1585));
AND2X1 g64847(.A (n_1582), .B (g4269), .Y (n_1583));
AND2X1 g64848(.A (n_1580), .B (g5097), .Y (n_1581));
INVX1 g65693(.A (n_1576), .Y (n_2064));
NAND3X1 g64936(.A (n_824), .B (g5216), .C (g25114), .Y (n_1575));
NAND3X1 g64940(.A (n_819), .B (n_2352), .C (g6255), .Y (n_1574));
XOR2X1 g65009(.A (g9251), .B (n_1570), .Y (n_1571));
NAND3X1 g61365(.A (g19357), .B (n_415), .C (n_635), .Y (n_1569));
AOI22X1 g65021(.A0 (n_636), .A1 (g_15740), .B0 (n_588), .B1 (n_708),.Y (n_1568));
AOI22X1 g65025(.A0 (n_1290), .A1 (g_22379), .B0 (n_691), .B1(g_19113), .Y (n_1567));
AND2X1 g65226(.A (n_10984), .B (g4955), .Y (n_1564));
NAND2X1 g65227(.A (n_1562), .B (n_162), .Y (n_1563));
AOI21X1 g65229(.A0 (n_268), .A1 (n_4980), .B0 (g4760), .Y (n_1561));
AOI21X1 g65231(.A0 (n_524), .A1 (n_11070), .B0 (g4894), .Y (n_1560));
XOR2X1 g65008(.A (g9019), .B (n_1556), .Y (n_1557));
AND2X1 g65277(.A (n_1554), .B (n_1631), .Y (n_1555));
NAND2X1 g65281(.A (n_10678), .B (n_10667), .Y (n_2452));
NAND2X1 g65288(.A (g6513), .B (n_4322), .Y (n_1553));
AND2X1 g65296(.A (n_3030), .B (n_1550), .Y (n_2747));
OR4X1 g65301(.A (n_954), .B (g8785), .C (g8783), .D (g8784), .Y(n_1552));
NAND2X1 g65311(.A (g3470), .B (n_4320), .Y (n_1551));
AND2X1 g65312(.A (n_3030), .B (n_1554), .Y (n_3048));
AND2X1 g65315(.A (n_1550), .B (n_1549), .Y (n_3021));
AND2X1 g65318(.A (n_1631), .B (n_3025), .Y (n_2115));
AND2X1 g65321(.A (n_3025), .B (n_1549), .Y (n_2457));
OR2X1 g65323(.A (n_1559), .B (n_10499), .Y (n_1548));
NAND2X1 g65327(.A (g3821), .B (n_4314), .Y (n_1547));
AOI21X1 g65345(.A0 (n_442), .A1 (n_241), .B0 (n_9371), .Y (n_2677));
NAND3X1 g65358(.A (n_1313), .B (g4076), .C (n_245), .Y (n_1546));
NAND2X1 g65366(.A (g5821), .B (n_4327), .Y (n_1545));
NOR2X1 g65373(.A (n_956), .B (n_2111), .Y (n_1544));
AND2X1 g65375(.A (n_1536), .B (n_1543), .Y (n_6394));
NAND3X1 g65379(.A (n_1559), .B (n_1541), .C (n_1540), .Y (n_1542));
NAND2X1 g65380(.A (g3119), .B (n_4316), .Y (n_1539));
NOR2X1 g65381(.A (n_965), .B (n_1263), .Y (n_2113));
NAND3X1 g65383(.A (n_10499), .B (n_1538), .C (n_11221), .Y (n_2451));
NAND2X1 g65391(.A (n_1536), .B (n_6399), .Y (n_1537));
NAND2X1 g65402(.A (g5475), .B (n_4329), .Y (n_1535));
AOI22X1 g65406(.A0 (n_608), .A1 (n_1533), .B0 (n_1532), .B1 (n_1531),.Y (n_1534));
AOI22X1 g65407(.A0 (n_620), .A1 (n_1529), .B0 (n_1528), .B1 (n_1527),.Y (n_1530));
NAND3X1 g65412(.A (n_1488), .B (g5272), .C (g25114), .Y (n_11195));
AOI22X1 g65416(.A0 (n_675), .A1 (n_368), .B0 (n_450), .B1 (n_1524),.Y (n_1525));
AOI22X1 g65431(.A0 (n_611), .A1 (n_362), .B0 (n_380), .B1 (n_1522),.Y (n_1523));
AOI22X1 g65451(.A0 (n_1520), .A1 (n_1519), .B0 (n_1518), .B1(n_1517), .Y (n_1521));
AOI22X1 g65458(.A0 (n_1515), .A1 (n_278), .B0 (n_1514), .B1(n_10996), .Y (n_1516));
AOI22X1 g65489(.A0 (n_1510), .A1 (g25167), .B0 (n_1509), .B1(n_10616), .Y (n_1511));
AOI22X1 g65490(.A0 (n_1506), .A1 (n_213), .B0 (n_1505), .B1(n_10789), .Y (n_1507));
XOR2X1 g65505(.A (g1579), .B (n_1502), .Y (n_1503));
INVX2 g65507(.A (n_1845), .Y (n_2127));
INVX1 g65509(.A (n_1500), .Y (n_2119));
INVX1 g65513(.A (n_1848), .Y (n_2131));
INVX2 g65514(.A (n_1854), .Y (n_2143));
INVX1 g65517(.A (n_6806), .Y (n_2447));
INVX2 g65518(.A (n_8548), .Y (n_1499));
INVX2 g65526(.A (n_1494), .Y (n_2133));
INVX1 g65614(.A (n_1493), .Y (n_1662));
OR2X1 g65630(.A (n_581), .B (n_3849), .Y (n_2062));
NAND2X1 g65635(.A (n_745), .B (g7916), .Y (n_1491));
AND2X1 g65695(.A (n_1488), .B (g25114), .Y (n_2077));
NOR2X1 g65702(.A (n_807), .B (n_1486), .Y (n_1487));
NOR2X1 g65712(.A (n_744), .B (n_1482), .Y (n_1483));
NAND2X1 g65718(.A (n_1480), .B (n_1177), .Y (n_1481));
NOR2X1 g65720(.A (n_786), .B (g4049), .Y (n_1479));
NAND2X1 g65724(.A (n_1147), .B (n_1584), .Y (n_1478));
NAND2X1 g65726(.A (n_1476), .B (n_1222), .Y (n_1477));
NOR2X1 g65729(.A (n_814), .B (n_1482), .Y (n_1475));
NOR2X1 g65732(.A (n_11124), .B (g3698), .Y (n_1474));
NOR2X1 g65734(.A (n_794), .B (g3347), .Y (n_1473));
NAND2X1 g65735(.A (n_1158), .B (n_1471), .Y (n_1472));
NAND2X1 g65738(.A (n_1149), .B (n_1471), .Y (n_1470));
NOR2X1 g65740(.A (n_810), .B (n_1468), .Y (n_1469));
NOR2X1 g65741(.A (n_1468), .B (n_411), .Y (n_1467));
NAND2X1 g65744(.A (n_1412), .B (n_1476), .Y (n_1466));
NOR2X1 g65746(.A (n_718), .B (n_1464), .Y (n_1465));
NAND2X1 g65748(.A (n_1480), .B (n_1227), .Y (n_1463));
NAND2X1 g65752(.A (n_1734), .B (n_1267), .Y (n_1462));
AND2X1 g65757(.A (n_2432), .B (n_1461), .Y (n_2039));
NOR2X1 g65759(.A (n_739), .B (n_1459), .Y (n_1460));
NAND2X1 g65768(.A (n_1194), .B (n_1455), .Y (n_1456));
NAND2X1 g65771(.A (n_6399), .B (n_6398), .Y (n_1454));
NAND2X1 g65772(.A (n_1403), .B (n_1480), .Y (n_1453));
NAND2X1 g65774(.A (n_1455), .B (n_1145), .Y (n_1452));
NAND2X1 g65776(.A (n_1450), .B (n_1210), .Y (n_1451));
NAND2X1 g65780(.A (n_1207), .B (n_1450), .Y (n_1449));
NAND2X1 g65785(.A (n_1201), .B (n_1450), .Y (n_1448));
NAND2X1 g65790(.A (n_1450), .B (n_1199), .Y (n_1447));
NAND2X1 g65795(.A (n_1445), .B (n_1216), .Y (n_1446));
NAND2X1 g65801(.A (n_1442), .B (g1536), .Y (n_1444));
NOR2X1 g65802(.A (n_1442), .B (n_3849), .Y (n_1443));
NAND2X1 g65814(.A (n_1440), .B (n_1191), .Y (n_1441));
NAND2X1 g65820(.A (n_1185), .B (n_1440), .Y (n_1439));
NAND2X1 g65821(.A (n_1399), .B (n_1480), .Y (n_1438));
NAND2X1 g65826(.A (n_1455), .B (n_1169), .Y (n_1437));
NAND2X1 g65828(.A (n_1181), .B (n_1440), .Y (n_1436));
NAND2X1 g65831(.A (n_1440), .B (n_1175), .Y (n_1435));
INVX1 g65836(.A (n_1434), .Y (n_2067));
NAND2X1 g65842(.A (n_1471), .B (n_1143), .Y (n_1433));
NAND2X1 g65844(.A (n_1395), .B (n_1445), .Y (n_1432));
NAND2X1 g65852(.A (n_1246), .B (n_1455), .Y (n_1431));
NOR2X1 g65860(.A (n_748), .B (g4616), .Y (n_1429));
NOR2X1 g65863(.A (n_893), .B (n_1486), .Y (n_1428));
NAND2X1 g65869(.A (n_1584), .B (n_1135), .Y (n_1427));
NAND2X1 g65872(.A (n_772), .B (n_1173), .Y (n_1655));
AND2X1 g65873(.A (n_6406), .B (n_6398), .Y (n_6404));
NOR2X1 g65882(.A (g4737), .B (n_8776), .Y (n_1426));
NAND2X1 g62021(.A (g_18902), .B (n_4754), .Y (n_2345));
NAND2X1 g65894(.A (n_1476), .B (n_1234), .Y (n_1425));
NAND2X1 g65898(.A (n_1407), .B (n_1476), .Y (n_1424));
NOR2X1 g65905(.A (n_791), .B (n_1325), .Y (n_1423));
INVX1 g65910(.A (n_1422), .Y (n_4637));
NAND3X1 g65918(.A (n_11113), .B (n_719), .C (g_20951), .Y (n_1652));
NAND2X1 g65932(.A (n_1471), .B (n_1214), .Y (n_1419));
NAND2X1 g65933(.A (n_1584), .B (n_896), .Y (n_1418));
NOR2X1 g65937(.A (n_789), .B (n_659), .Y (n_1417));
NAND2X1 g65938(.A (n_1394), .B (n_1445), .Y (n_1416));
NAND2X1 g65940(.A (n_1445), .B (n_585), .Y (n_1415));
NAND2X1 g65942(.A (n_3812), .B (n_6406), .Y (n_1414));
NAND2X1 g65947(.A (n_1412), .B (n_1411), .Y (n_1413));
NAND2X1 g65950(.A (n_877), .B (n_6923), .Y (n_1409));
NAND2X1 g65952(.A (n_1407), .B (n_1411), .Y (n_1408));
NAND2X1 g65965(.A (n_1403), .B (n_1402), .Y (n_1404));
NAND2X1 g65967(.A (n_1403), .B (n_1762), .Y (n_1401));
NAND2X1 g65975(.A (n_1399), .B (n_1402), .Y (n_1400));
NAND2X1 g65978(.A (n_1399), .B (n_1762), .Y (n_1398));
NAND2X1 g65983(.A (n_1407), .B (n_1777), .Y (n_1397));
NAND2X1 g62041(.A (n_4757), .B (n_1599), .Y (n_1646));
OR2X1 g65991(.A (n_1395), .B (n_1394), .Y (n_1396));
NAND2X1 g65995(.A (n_1394), .B (n_1718), .Y (n_1393));
NAND2X1 g65996(.A (n_1394), .B (n_1391), .Y (n_1392));
AOI21X1 g66003(.A0 (g5188), .A1 (n_388), .B0 (n_1402), .Y (n_1390));
AOI21X1 g66009(.A0 (g5535), .A1 (n_383), .B0 (n_1411), .Y (n_1388));
AOI21X1 g66017(.A0 (g5881), .A1 (n_215), .B0 (n_1382), .Y (n_1384));
OAI21X1 g66018(.A0 (g17646), .A1 (g13068), .B0 (n_779), .Y (n_1381));
AOI21X1 g66021(.A0 (g6227), .A1 (n_330), .B0 (n_1377), .Y (n_1380));
AOI22X1 g66027(.A0 (n_10107), .A1 (n_723), .B0 (n_10108), .B1(n_552), .Y (n_10551));
AOI21X1 g66028(.A0 (g6573), .A1 (n_261), .B0 (n_1391), .Y (n_1375));
AOI21X1 g66030(.A0 (g3179), .A1 (n_370), .B0 (n_1370), .Y (n_1373));
AOI21X1 g66036(.A0 (g3530), .A1 (n_365), .B0 (n_1367), .Y (n_1369));
AOI21X1 g66046(.A0 (g3881), .A1 (n_303), .B0 (n_1364), .Y (n_1366));
AOI21X1 g66080(.A0 (n_6527), .A1 (n_3388), .B0 (n_3391), .Y (n_1363));
NAND4X1 g66086(.A (g17711), .B (g17580), .C (g12300), .D (g14694), .Y(n_2881));
NAND4X1 g66090(.A (g17778), .B (g17688), .C (g12470), .D (g14828), .Y(n_2871));
NAND4X1 g66095(.A (n_110), .B (g5046), .C (n_1356), .D (g5052), .Y(n_2044));
OAI21X1 g61479(.A0 (n_556), .A1 (g1333), .B0 (g12923), .Y (n_2060));
DFFSRX1 g3267_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16718), .Q (g16603), .QN ());
NAND2X1 g65420(.A (n_709), .B (n_1353), .Y (n_1354));
DFFSRX1 g3618_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g16744), .Q (g16627), .QN ());
NAND2X1 g66596(.A (g1489), .B (n_9717), .Y (n_1628));
INVX1 g66633(.A (n_10214), .Y (n_1625));
AND2X1 g66661(.A (n_1352), .B (g8719), .Y (n_2001));
NAND3X1 g61513(.A (g19334), .B (n_325), .C (n_496), .Y (n_1351));
NOR2X1 g66878(.A (n_7260), .B (g4349), .Y (n_1349));
NAND2X1 g63875(.A (n_1331), .B (n_10119), .Y (n_2710));
OR2X1 g63876(.A (n_1331), .B (n_10119), .Y (n_1330));
INVX1 g63892(.A (n_1840), .Y (n_1329));
NAND2X1 g63894(.A (n_1328), .B (n_10112), .Y (n_2696));
OR2X1 g63896(.A (n_1328), .B (n_10112), .Y (n_1327));
NOR2X1 g65797(.A (n_1486), .B (n_1325), .Y (n_1326));
NAND2X1 g65962(.A (n_1412), .B (n_1777), .Y (n_1322));
INVX1 g66757(.A (n_1321), .Y (n_2019));
DFFSRX1 g6675_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12470), .Q (g14828), .QN ());
DFFSRX1 g5637_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12300), .Q (g14694), .QN ());
OR2X1 g61538(.A (n_470), .B (n_724), .Y (n_1315));
NAND3X1 g65343(.A (n_1313), .B (n_1312), .C (n_118), .Y (n_1737));
NOR2X1 g62659(.A (n_8585), .B (g3343), .Y (n_1311));
NOR2X1 g62660(.A (n_1272), .B (g3694), .Y (n_1310));
OR2X1 g64604(.A (n_980), .B (n_1307), .Y (n_1308));
NOR2X1 g65703(.A (n_1524), .B (n_433), .Y (n_1304));
AOI21X1 g64704(.A0 (n_1299), .A1 (g34028), .B0 (n_680), .Y (n_1300));
NAND2X1 g65897(.A (n_8796), .B (n_8591), .Y (n_1298));
XOR2X1 g64780(.A (n_1295), .B (n_982), .Y (n_1296));
NAND3X1 g64942(.A (n_663), .B (g1564), .C (g1554), .Y (n_2938));
NAND3X1 g64954(.A (n_971), .B (n_518), .C (n_8799), .Y (n_2945));
NAND3X1 g64966(.A (n_1093), .B (n_2443), .C (g5563), .Y (n_1293));
NAND3X1 g64968(.A (n_1011), .B (n_2432), .C (g6601), .Y (n_1292));
NOR2X1 g65279(.A (n_1290), .B (g_22379), .Y (n_1291));
DFFSRX1 g3983_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g11418), .Q (g13966), .QN ());
NAND2X1 g66779(.A (n_1285), .B (n_11055), .Y (n_1286));
AOI21X1 g65228(.A0 (n_374), .A1 (n_4982), .B0 (g4749), .Y (n_1283));
AOI21X1 g65230(.A0 (n_339), .A1 (n_4978), .B0 (g4771), .Y (n_1282));
NAND2X1 g65320(.A (n_471), .B (n_1285), .Y (n_1279));
NAND2X1 g65352(.A (n_1820), .B (g8839), .Y (n_1278));
NOR2X1 g65370(.A (n_1276), .B (n_1275), .Y (n_1277));
NOR2X1 g65397(.A (g4878), .B (n_1274), .Y (n_1826));
INVX1 g66421(.A (n_1272), .Y (n_1273));
AOI21X1 g65445(.A0 (g34026), .A1 (g21245), .B0 (n_676), .Y (n_1271));
NAND2X1 g66414(.A (n_596), .B (n_10013), .Y (n_5378));
XOR2X1 g66025(.A (g6159), .B (n_3589), .Y (n_1269));
DFFSRX1 g6023_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17819), .Q (g14673), .QN ());
DFFSRX1 g6715_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17871), .Q (g14749), .QN ());
DFFSRX1 g4477_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g4474), .Q (g4477), .QN ());
NAND2X1 g65615(.A (n_771), .B (g5029), .Y (n_1493));
NAND2X1 g65616(.A (n_1267), .B (n_3624), .Y (n_1268));
NOR2X1 g65617(.A (n_578), .B (g5511), .Y (n_1772));
INVX1 g65618(.A (n_1554), .Y (n_1266));
NAND2X1 g65625(.A (n_1264), .B (n_1214), .Y (n_4324));
NOR2X1 g65626(.A (n_566), .B (g6203), .Y (n_1770));
INVX1 g65633(.A (n_1263), .Y (n_2153));
INVX1 g65636(.A (n_3025), .Y (n_1262));
NOR2X1 g65639(.A (n_580), .B (g3506), .Y (n_1752));
NAND2X1 g65640(.A (g1950), .B (n_579), .Y (n_1261));
NAND2X1 g65642(.A (g1816), .B (n_557), .Y (n_1260));
NAND2X1 g65647(.A (g2084), .B (n_558), .Y (n_1257));
NAND2X1 g65649(.A (n_10724), .B (g7916), .Y (n_1255));
NOR2X1 g65651(.A (n_575), .B (g3857), .Y (n_1744));
INVX1 g65655(.A (n_1812), .Y (g26801));
INVX1 g65666(.A (n_1252), .Y (n_4628));
NOR2X1 g65669(.A (n_587), .B (g6549), .Y (n_1765));
NAND2X1 g65670(.A (n_594), .B (n_662), .Y (n_1251));
NOR2X1 g65674(.A (n_479), .B (g5164), .Y (n_1763));
INVX1 g65675(.A (n_1550), .Y (n_1250));
NOR2X1 g65681(.A (n_565), .B (g3155), .Y (n_1767));
NAND2X1 g65694(.A (n_653), .B (n_8677), .Y (n_1576));
NOR2X1 g65696(.A (n_1531), .B (n_187), .Y (n_1248));
AND2X1 g65697(.A (n_1246), .B (n_1245), .Y (n_1247));
AND2X1 g65709(.A (n_1243), .B (n_1242), .Y (n_1244));
NAND3X1 g65714(.A (g2130), .B (n_1240), .C (g2145), .Y (n_1241));
NOR2X1 g65719(.A (n_673), .B (n_1154), .Y (n_1239));
INVX1 g65722(.A (n_4617), .Y (n_1238));
NAND2X1 g65730(.A (n_1236), .B (n_827), .Y (n_1237));
NAND2X1 g65731(.A (n_1411), .B (n_1234), .Y (n_1235));
NOR2X1 g65742(.A (n_1464), .B (n_1224), .Y (n_1232));
NAND2X1 g65743(.A (n_1230), .B (n_836), .Y (n_1231));
AND2X1 g65751(.A (n_1762), .B (n_1227), .Y (n_1228));
NAND3X1 g65753(.A (n_269), .B (n_812), .C (g2453), .Y (n_1226));
NOR2X1 g65754(.A (n_822), .B (n_1224), .Y (n_1225));
AND2X1 g65756(.A (n_1411), .B (n_1222), .Y (n_1223));
NOR2X1 g65758(.A (n_3391), .B (n_3388), .Y (n_1221));
INVX1 g65761(.A (n_1219), .Y (n_1220));
NAND2X1 g65767(.A (n_1718), .B (n_1216), .Y (n_1217));
NAND2X1 g65770(.A (n_1723), .B (n_1214), .Y (n_1215));
NOR2X1 g65777(.A (n_1212), .B (n_3812), .Y (n_1213));
NAND2X1 g65778(.A (n_1751), .B (n_1210), .Y (n_1211));
NAND2X1 g65779(.A (n_1367), .B (n_1210), .Y (n_1209));
AND2X1 g65782(.A (n_1207), .B (n_1206), .Y (n_1208));
NOR2X1 g65783(.A (n_817), .B (n_1224), .Y (n_1205));
AND2X1 g65788(.A (n_1201), .B (n_1206), .Y (n_1202));
AND2X1 g65791(.A (n_1751), .B (n_1199), .Y (n_1200));
AND2X1 g65792(.A (n_1367), .B (n_1199), .Y (n_1198));
AND2X1 g65808(.A (n_1194), .B (n_1245), .Y (n_1195));
NAND3X1 g65812(.A (n_291), .B (n_806), .C (g1894), .Y (n_1193));
NAND2X1 g65816(.A (n_1743), .B (n_1191), .Y (n_1192));
NAND2X1 g65818(.A (n_1364), .B (n_1191), .Y (n_1189));
AND2X1 g65819(.A (n_8832), .B (g7916), .Y (n_1188));
AND2X1 g65824(.A (n_1777), .B (n_1222), .Y (n_1187));
AND2X1 g65825(.A (n_1185), .B (n_1184), .Y (n_1186));
NAND2X1 g65827(.A (n_1024), .B (n_10563), .Y (n_1183));
AND2X1 g65829(.A (n_1181), .B (n_1184), .Y (n_1182));
NAND2X1 g65830(.A (n_1179), .B (n_1165), .Y (n_1180));
NAND2X1 g65833(.A (n_1402), .B (n_1177), .Y (n_1178));
AND2X1 g65834(.A (n_1743), .B (n_1175), .Y (n_1176));
NAND2X1 g65837(.A (n_644), .B (n_11209), .Y (n_1434));
AND2X1 g65839(.A (n_1364), .B (n_1175), .Y (n_1174));
OR2X1 g65840(.A (n_1173), .B (g5029), .Y (n_7010));
NAND2X1 g65856(.A (n_1725), .B (n_1169), .Y (n_1170));
NOR2X1 g65858(.A (n_1527), .B (n_382), .Y (n_1168));
NAND2X1 g65859(.A (n_1391), .B (n_1216), .Y (n_1167));
NAND2X1 g65864(.A (n_978), .B (n_1165), .Y (n_1166));
NAND2X1 g65870(.A (n_1762), .B (n_1177), .Y (n_1164));
NAND2X1 g65875(.A (g_7220), .B (g8291), .Y (n_1731));
NAND3X1 g65880(.A (n_444), .B (n_804), .C (g1760), .Y (n_1163));
NAND3X1 g65881(.A (n_377), .B (n_730), .C (g2319), .Y (n_1162));
NAND2X1 g65885(.A (n_1160), .B (n_831), .Y (n_1161));
AND2X1 g65886(.A (n_1158), .B (n_1264), .Y (n_1159));
NOR2X1 g65892(.A (n_795), .B (n_1154), .Y (n_1155));
NAND2X1 g65893(.A (n_1377), .B (n_1214), .Y (n_1153));
AND2X1 g65902(.A (n_1395), .B (n_590), .Y (n_1152));
AND2X1 g65903(.A (n_1149), .B (n_1264), .Y (n_1150));
AND2X1 g65904(.A (n_1147), .B (n_1242), .Y (n_1148));
AND2X1 g65906(.A (n_1382), .B (n_1145), .Y (n_1146));
AND2X1 g65907(.A (n_1377), .B (n_1143), .Y (n_1144));
NAND2X1 g65911(.A (n_1179), .B (g13272), .Y (n_1422));
NAND2X1 g65925(.A (n_1138), .B (n_839), .Y (n_1139));
NAND2X1 g65926(.A (g5913), .B (n_10508), .Y (n_1137));
INVX1 g65929(.A (n_1536), .Y (n_6402));
NAND2X1 g65931(.A (n_1370), .B (n_1135), .Y (n_1136));
NAND3X1 g65945(.A (g2130), .B (g2138), .C (g2145), .Y (n_1133));
NAND2X1 g65946(.A (n_1777), .B (n_1234), .Y (n_1131));
NAND2X1 g65949(.A (n_1181), .B (n_1743), .Y (n_1130));
NAND2X1 g65955(.A (n_1158), .B (n_1723), .Y (n_1128));
NAND2X1 g65956(.A (n_1149), .B (n_1723), .Y (n_1127));
INVX1 g65958(.A (n_1124), .Y (n_1405));
NAND2X1 g65960(.A (n_1147), .B (n_1370), .Y (n_1123));
NAND2X1 g65963(.A (n_1395), .B (n_1718), .Y (n_1122));
NAND2X1 g65966(.A (n_1147), .B (n_1758), .Y (n_1121));
NAND2X1 g65968(.A (n_1246), .B (n_1725), .Y (n_1120));
NAND2X1 g65971(.A (n_1207), .B (n_1751), .Y (n_1119));
NAND2X1 g65972(.A (n_1207), .B (n_1367), .Y (n_1118));
NAND2X1 g65973(.A (n_1201), .B (n_1751), .Y (n_1117));
NAND2X1 g65974(.A (n_1201), .B (n_1367), .Y (n_1116));
OR2X1 g65976(.A (n_1207), .B (n_1201), .Y (n_1115));
NAND2X1 g65977(.A (n_1194), .B (n_1382), .Y (n_1114));
OR2X1 g65979(.A (n_1185), .B (n_1181), .Y (n_1113));
NAND2X1 g65980(.A (n_1185), .B (n_1743), .Y (n_1112));
NAND2X1 g65981(.A (n_1185), .B (n_1364), .Y (n_1111));
NAND2X1 g65982(.A (n_1181), .B (n_1364), .Y (n_1110));
OR2X1 g65985(.A (n_1243), .B (n_1147), .Y (n_1109));
NAND2X1 g65988(.A (n_1194), .B (n_1725), .Y (n_1108));
NAND2X1 g65989(.A (n_1158), .B (n_1377), .Y (n_1107));
NAND2X1 g65990(.A (n_1149), .B (n_1377), .Y (n_1106));
NAND2X1 g65993(.A (n_1243), .B (n_1370), .Y (n_1105));
NAND2X1 g65997(.A (n_1246), .B (n_1382), .Y (n_1104));
NAND2X1 g65998(.A (n_1395), .B (n_1391), .Y (n_1103));
NAND2X1 g65999(.A (n_1243), .B (n_1758), .Y (n_1102));
XOR2X1 g66000(.A (g5120), .B (n_3618), .Y (n_1101));
OAI21X1 g66014(.A0 (n_423), .A1 (n_11050), .B0 (n_1100), .Y (n_1845));
XOR2X1 g66031(.A (g6505), .B (n_3604), .Y (n_1099));
XOR2X1 g66032(.A (g5813), .B (n_3611), .Y (n_1098));
OAI21X1 g66037(.A0 (n_11160), .A1 (g_6165), .B0 (n_818), .Y (n_1848));
XOR2X1 g66052(.A (g5467), .B (n_3616), .Y (n_1097));
OAI21X1 g66058(.A0 (n_10369), .A1 (g_4409), .B0 (n_823), .Y (n_1854));
AOI21X1 g66060(.A0 (n_512), .A1 (g4601), .B0 (n_820), .Y (n_1096));
XOR2X1 g66069(.A (n_364), .B (g_22552), .Y (n_1095));
NAND2X1 g66732(.A (g17577), .B (g17519), .Y (n_1094));
AOI21X1 g66075(.A0 (n_776), .A1 (n_409), .B0 (n_1093), .Y (n_1494));
NAND4X1 g66085(.A (g17674), .B (g17519), .C (g12238), .D (g14662), .Y(n_3171));
NAND4X1 g66087(.A (g_15380), .B (g_15381), .C (n_413), .D (g_16792),.Y (n_1090));
NAND4X1 g66093(.A (g17760), .B (g17649), .C (g12422), .D (g14779), .Y(n_2729));
NAND4X1 g66094(.A (g17739), .B (g17607), .C (g12350), .D (g14738), .Y(n_2732));
NOR2X1 g65622(.A (n_589), .B (g5857), .Y (n_1727));
MX2X1 g66151(.A (n_527), .B (g14662), .S0 (g17674), .Y (n_1085));
MX2X1 g66152(.A (n_669), .B (g14694), .S0 (g17711), .Y (n_1084));
MX2X1 g66153(.A (n_549), .B (g14779), .S0 (g17760), .Y (n_1083));
MX2X1 g66155(.A (n_538), .B (g14828), .S0 (g17778), .Y (n_1082));
MX2X1 g66157(.A (g_22552), .B (n_364), .S0 (g_16404), .Y (n_1081));
XOR2X1 g66160(.A (g5527), .B (n_1234), .Y (n_1079));
XOR2X1 g66161(.A (g5180), .B (n_1177), .Y (n_1077));
XOR2X1 g66168(.A (g3171), .B (n_1135), .Y (n_1075));
XOR2X1 g66169(.A (g3522), .B (n_1210), .Y (n_1074));
XOR2X1 g66172(.A (g6219), .B (n_1214), .Y (n_1072));
XOR2X1 g66181(.A (g6565), .B (n_1216), .Y (n_1071));
XOR2X1 g66188(.A (g5873), .B (n_1169), .Y (n_1069));
DFFSRX1 g5331_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17787), .Q (g14597), .QN ());
DFFSRX1 g4012_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13966), .Q (g16775), .QN ());
INVX1 g66355(.A (n_1064), .Y (n_1065));
INVX1 g66390(.A (n_1062), .Y (n_1063));
INVX1 g66559(.A (n_1059), .Y (n_1060));
INVX1 g66566(.A (n_2339), .Y (n_1058));
INVX1 g66607(.A (n_1055), .Y (n_4878));
NAND2X1 g66642(.A (g17604), .B (g17580), .Y (n_1054));
NOR2X1 g66693(.A (n_5917), .B (g2351), .Y (n_1053));
NOR2X1 g66743(.A (n_5921), .B (g2485), .Y (n_1052));
NAND2X1 g66758(.A (g3466), .B (n_10950), .Y (n_1321));
DFFSRX1 g6369_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17845), .Q (g14705), .QN ());
NAND2X1 g66799(.A (g17685), .B (g17649), .Y (n_1046));
NOR2X1 g66843(.A (n_5925), .B (g1926), .Y (n_1044));
INVX1 g66846(.A (n_3459), .Y (n_1043));
NOR2X1 g66904(.A (n_5996), .B (g1792), .Y (n_1040));
DFFSRX1 g5677_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17813), .Q (g14635), .QN ());
INVX2 g67909(.A (n_5402), .Y (n_3894));
INVX1 g62237(.A (n_4754), .Y (n_2878));
AND2X1 g62259(.A (n_8591), .B (g13259), .Y (n_4764));
AND2X1 g62262(.A (n_8832), .B (g13259), .Y (n_4761));
OR2X1 g65994(.A (n_10567), .B (n_1024), .Y (n_10550));
NAND2X1 g66590(.A (g17722), .B (g17688), .Y (n_1021));
OR2X1 g65992(.A (n_1158), .B (n_1149), .Y (n_1017));
AND2X1 g65396(.A (g4878), .B (n_1274), .Y (n_1016));
NOR2X1 g61630(.A (g4434), .B (n_596), .Y (n_1015));
AND2X1 g63893(.A (n_1307), .B (g4659), .Y (n_1840));
NOR2X1 g65733(.A (n_1522), .B (n_418), .Y (n_1014));
OR2X1 g65389(.A (n_989), .B (n_10499), .Y (n_1013));
AOI21X1 g66081(.A0 (n_11185), .A1 (n_322), .B0 (n_1011), .Y (n_1500));
DFFSRX1 g5630_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17580), .Q (g17604), .QN ());
DFFSRX1 g5290_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12238), .Q (g14662), .QN ());
DFFSRX1 g4864_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g34034), .Q (g34035), .QN ());
DFFSRX1 g6329_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12422), .Q (g14779), .QN ());
DFFSRX1 g6668_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17688), .Q (g17722), .QN ());
DFFSRX1 g5983_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12350), .Q (g14738), .QN ());
DFFSRX1 g3632_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g11388), .Q (g13926), .QN ());
DFFSRX1 g3281_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g11349), .Q (g13895), .QN ());
DFFSRX1 g6322_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17649), .Q (g17685), .QN ());
OR2X1 g65954(.A (n_1194), .B (n_1246), .Y (n_1002));
DFFSRX1 g5283_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17519), .Q (g17577), .QN ());
NAND2X1 g65765(.A (n_1382), .B (n_1169), .Y (n_999));
XOR2X1 g66174(.A (g3873), .B (n_1191), .Y (n_998));
NOR2X1 g65736(.A (n_983), .B (n_1154), .Y (n_995));
NOR2X1 g65372(.A (n_151), .B (g4878), .Y (n_994));
NAND2X1 g65745(.A (n_1758), .B (n_1135), .Y (n_993));
OR2X1 g65721(.A (g_9174), .B (g2980), .Y (n_992));
NOR2X1 g65329(.A (n_6707), .B (n_989), .Y (n_991));
NAND4X1 g64601(.A (n_988), .B (n_987), .C (n_986), .D (g4688), .Y(n_4839));
INVX2 g68008(.A (g25219), .Y (n_1695));
INVX1 g66416(.A (n_983), .Y (n_1412));
NOR2X1 g64840(.A (n_474), .B (n_307), .Y (n_1331));
NOR2X1 g64849(.A (n_982), .B (n_1295), .Y (n_1328));
NOR3X1 g64899(.A (g_16404), .B (g_22552), .C (n_364), .Y (n_5582));
XOR2X1 g66061(.A (n_2485), .B (g1472), .Y (n_981));
NOR2X1 g64914(.A (n_69), .B (g4653), .Y (n_980));
INVX1 g66447(.A (n_978), .Y (n_1442));
NOR2X1 g66793(.A (g3171), .B (g3179), .Y (n_1584));
OAI21X1 g65677(.A0 (g3480), .A1 (g3494), .B0 (n_10949), .Y (n_1550));
XOR2X1 g66034(.A (n_1799), .B (n_2699), .Y (n_977));
OAI21X1 g65683(.A0 (g5485), .A1 (g5499), .B0 (n_8921), .Y (n_1631));
XOR2X1 g66033(.A (n_975), .B (n_6025), .Y (n_976));
OR2X1 g65679(.A (n_948), .B (g4628), .Y (n_974));
DFFSRX1 g4674_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g34026), .Q (g34027), .QN ());
DFFSRX1 g4681_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g34027), .Q (g34028), .QN ());
NAND2X1 g65667(.A (n_908), .B (g13272), .Y (n_1252));
NAND2X1 g65653(.A (n_973), .B (n_1234), .Y (n_4329));
NAND2X1 g65657(.A (n_970), .B (n_1177), .Y (n_1812));
XOR2X1 g66026(.A (g1300), .B (n_3383), .Y (n_969));
NAND3X1 g65861(.A (n_196), .B (n_6967), .C (g5057), .Y (n_2045));
NAND2X1 g65621(.A (n_1245), .B (n_1169), .Y (n_4327));
OR2X1 g65623(.A (g2509), .B (n_8632), .Y (n_967));
INVX1 g65627(.A (n_1630), .Y (n_965));
OR2X1 g65631(.A (g2375), .B (n_8627), .Y (n_963));
NOR2X1 g65634(.A (n_343), .B (n_9297), .Y (n_1263));
NAND2X1 g65638(.A (n_1206), .B (n_1210), .Y (n_4320));
OR2X1 g65646(.A (n_309), .B (g17423), .Y (n_961));
NOR2X1 g65654(.A (n_429), .B (g2357), .Y (n_958));
OR2X1 g65660(.A (n_295), .B (g17400), .Y (n_957));
NAND2X1 g65661(.A (n_1312), .B (n_955), .Y (n_956));
NAND2X1 g65662(.A (n_1242), .B (n_1135), .Y (n_4316));
OR2X1 g65663(.A (n_220), .B (n_10871), .Y (n_954));
OAI21X1 g65664(.A0 (g3129), .A1 (g3143), .B0 (g35), .Y (n_3030));
OR2X1 g65668(.A (g2241), .B (n_8534), .Y (n_952));
AND2X1 g65671(.A (n_188), .B (n_955), .Y (n_1313));
NAND2X1 g65672(.A (n_590), .B (n_1216), .Y (n_4322));
OAI21X1 g65673(.A0 (g3831), .A1 (g3845), .B0 (n_10949), .Y (n_1549));
NOR2X1 g65678(.A (n_302), .B (g2112), .Y (n_950));
NAND2X1 g65680(.A (n_948), .B (g4628), .Y (n_2980));
NOR2X1 g65682(.A (n_436), .B (g2671), .Y (n_947));
INVX1 g68403(.A (n_946), .Y (n_3707));
NOR2X1 g65684(.A (n_298), .B (g1798), .Y (n_943));
OR2X1 g65685(.A (g2643), .B (n_10720), .Y (n_942));
OR2X1 g65686(.A (g1682), .B (n_10271), .Y (n_940));
AND2X1 g65723(.A (n_899), .B (g13272), .Y (n_4617));
NAND2X1 g65725(.A (n_323), .B (n_2550), .Y (n_938));
XOR2X1 g66038(.A (g3111), .B (n_3609), .Y (n_937));
NAND2X1 g65775(.A (n_336), .B (n_933), .Y (n_934));
NAND2X1 g65789(.A (n_441), .B (n_2306), .Y (n_932));
AND2X1 g65793(.A (n_1199), .B (n_1206), .Y (n_931));
NAND3X1 g65805(.A (n_928), .B (g1624), .C (n_677), .Y (n_929));
NAND2X1 g65807(.A (n_240), .B (n_926), .Y (n_927));
NAND3X1 g65809(.A (n_399), .B (n_674), .C (g2028), .Y (n_925));
NOR3X1 g65822(.A (g_21778), .B (n_273), .C (g_19113), .Y (n_924));
OR4X1 g65832(.A (n_10113), .B (g1564), .C (g1554), .D (g1548), .Y(n_2108));
OR2X1 g66729(.A (g8416), .B (g7916), .Y (n_923));
AND2X1 g65841(.A (n_1175), .B (n_1184), .Y (n_921));
NOR2X1 g65850(.A (n_218), .B (n_143), .Y (n_10905));
NAND3X1 g65854(.A (n_919), .B (n_619), .C (g2185), .Y (n_920));
OR4X1 g65855(.A (g2657), .B (g2523), .C (g2255), .D (g2389), .Y(n_918));
AND2X1 g65857(.A (n_916), .B (n_8534), .Y (n_917));
NAND2X1 g65862(.A (n_376), .B (n_2293), .Y (n_915));
NAND2X1 g65877(.A (g1950), .B (n_6790), .Y (n_914));
AND2X1 g65883(.A (n_911), .B (n_8627), .Y (n_912));
AND2X1 g65884(.A (n_6399), .B (n_3641), .Y (n_1543));
AND2X1 g65888(.A (n_1145), .B (n_1245), .Y (n_910));
NAND2X1 g65899(.A (n_908), .B (n_1165), .Y (n_909));
NAND2X1 g65912(.A (n_408), .B (n_2780), .Y (n_906));
AND2X1 g65924(.A (n_904), .B (n_8632), .Y (n_905));
AND2X1 g65927(.A (n_902), .B (n_10720), .Y (n_903));
NOR2X1 g65930(.A (n_901), .B (n_3812), .Y (n_1536));
NAND2X1 g65935(.A (n_1165), .B (n_899), .Y (n_900));
NAND3X1 g65939(.A (g2130), .B (g2138), .C (n_308), .Y (n_898));
AND2X1 g65941(.A (n_896), .B (n_1242), .Y (n_897));
NAND3X1 g65943(.A (n_351), .B (n_610), .C (g2587), .Y (n_895));
NAND2X1 g65944(.A (n_338), .B (n_2521), .Y (n_894));
INVX1 g66380(.A (n_1718), .Y (n_893));
AOI21X1 g65987(.A0 (g_20073), .A1 (g_12433), .B0 (n_891), .Y(n_10552));
XOR2X1 g66002(.A (n_1813), .B (n_2718), .Y (n_890));
XOR2X1 g66006(.A (n_1794), .B (n_3007), .Y (n_888));
XOR2X1 g66008(.A (n_1810), .B (n_3011), .Y (n_887));
XOR2X1 g66011(.A (n_885), .B (n_5975), .Y (n_886));
XOR2X1 g66012(.A (n_883), .B (n_5978), .Y (n_884));
XOR2X1 g66016(.A (n_1807), .B (n_2684), .Y (n_882));
XOR2X1 g66020(.A (n_2084), .B (n_2704), .Y (n_881));
XOR2X1 g66022(.A (n_1805), .B (n_2686), .Y (n_880));
INVX1 g66451(.A (n_876), .Y (n_877));
AND2X1 g66737(.A (n_11177), .B (g17722), .Y (n_1461));
XOR2X1 g66035(.A (n_871), .B (n_4946), .Y (n_872));
OAI21X1 g65637(.A0 (g5138), .A1 (g5152), .B0 (n_10949), .Y (n_3025));
XOR2X1 g66043(.A (g3813), .B (n_3596), .Y (n_868));
XOR2X1 g66045(.A (n_866), .B (n_5972), .Y (n_867));
XOR2X1 g66047(.A (n_864), .B (n_5961), .Y (n_8755));
XOR2X1 g66048(.A (n_862), .B (n_5953), .Y (n_863));
XOR2X1 g66049(.A (n_860), .B (n_6017), .Y (n_861));
XOR2X1 g66050(.A (n_858), .B (n_5969), .Y (n_859));
XOR2X1 g66051(.A (n_856), .B (n_5964), .Y (n_857));
XOR2X1 g66054(.A (n_854), .B (n_4948), .Y (n_855));
XOR2X1 g66055(.A (n_852), .B (n_6020), .Y (n_10554));
XOR2X1 g66059(.A (n_2556), .B (g_16456), .Y (n_851));
XOR2X1 g66062(.A (n_2535), .B (g1478), .Y (n_849));
XOR2X1 g66070(.A (n_2529), .B (g_11413), .Y (n_848));
XOR2X1 g66072(.A (n_846), .B (n_4942), .Y (n_847));
XOR2X1 g66082(.A (g3462), .B (n_3601), .Y (n_845));
OAI21X1 g65620(.A0 (g5831), .A1 (g5845), .B0 (n_8921), .Y (n_1554));
NAND4X1 g66091(.A (g4489), .B (g4483), .C (g4492), .D (g4486), .Y(n_1562));
AOI22X1 g66092(.A0 (g3333), .A1 (g34035), .B0 (n_843), .B1 (g34034),.Y (n_844));
MX2X1 g66156(.A (n_371), .B (g14738), .S0 (g17739), .Y (n_842));
XOR2X1 g66158(.A (g1691), .B (n_4527), .Y (n_841));
XOR2X1 g66159(.A (n_4531), .B (n_839), .Y (n_840));
XOR2X1 g66163(.A (n_1796), .B (n_2692), .Y (n_838));
XOR2X1 g66166(.A (n_4187), .B (n_836), .Y (n_837));
XOR2X1 g66170(.A (g1448), .B (n_2538), .Y (n_835));
XOR2X1 g66171(.A (g2093), .B (n_4183), .Y (n_834));
XOR2X1 g66177(.A (g2250), .B (n_4906), .Y (n_833));
XOR2X1 g66178(.A (n_4529), .B (n_831), .Y (n_832));
XOR2X1 g66180(.A (g_18869), .B (n_2244), .Y (n_830));
XOR2X1 g66183(.A (g2652), .B (n_4726), .Y (n_829));
XOR2X1 g66184(.A (n_4190), .B (n_827), .Y (n_828));
CLKBUFX1 g66185(.A (n_6707), .Y (n_1559));
INVX1 g66208(.A (g_7220), .Y (n_826));
DFFSRX1 g3310_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13895), .Q (g16718), .QN ());
INVX1 g66284(.A (n_823), .Y (n_824));
INVX1 g66300(.A (n_822), .Y (n_1403));
INVX1 g66303(.A (n_820), .Y (n_821));
INVX1 g66312(.A (n_818), .Y (n_819));
INVX1 g66332(.A (n_817), .Y (n_1399));
INVX1 g66703(.A (n_6552), .Y (n_816));
INVX1 g66342(.A (n_1758), .Y (n_814));
NOR2X1 g66356(.A (n_812), .B (g2485), .Y (n_1064));
INVX1 g66370(.A (n_1723), .Y (n_810));
INVX1 g66377(.A (n_1138), .Y (n_808));
INVX1 g66386(.A (n_1391), .Y (n_807));
NOR2X1 g66391(.A (n_806), .B (g1926), .Y (n_1062));
AND2X1 g66392(.A (n_804), .B (g1792), .Y (n_805));
INVX1 g66422(.A (n_4682), .Y (n_1272));
INVX1 g66434(.A (n_802), .Y (n_803));
INVX1 g66454(.A (n_800), .Y (n_801));
NOR2X1 g66483(.A (n_804), .B (g1792), .Y (n_1667));
INVX1 g66485(.A (n_799), .Y (n_1599));
INVX1 g66489(.A (n_1236), .Y (n_798));
NOR2X1 g66492(.A (n_448), .B (n_662), .Y (n_797));
INVX1 g66505(.A (n_795), .Y (n_1407));
INVX1 g66516(.A (n_8572), .Y (n_794));
INVX1 g66520(.A (n_1160), .Y (n_793));
INVX1 g66535(.A (n_791), .Y (n_1394));
AND2X1 g66548(.A (n_812), .B (g2485), .Y (n_790));
INVX1 g66550(.A (n_3391), .Y (n_789));
INVX1 g66578(.A (n_6808), .Y (n_786));
NOR2X1 g66598(.A (g6565), .B (g6573), .Y (n_1445));
NOR2X1 g66599(.A (g4349), .B (n_1627), .Y (n_1734));
NAND2X1 g66608(.A (g3817), .B (n_10949), .Y (n_1055));
INVX1 g66613(.A (n_590), .Y (n_1325));
NAND2X1 g66618(.A (g4401), .B (g4392), .Y (n_784));
NOR2X1 g66619(.A (g1636), .B (n_4120), .Y (n_783));
NOR2X1 g66622(.A (g3522), .B (g3530), .Y (n_1450));
NOR2X1 g66625(.A (n_5928), .B (g2619), .Y (n_782));
OR2X1 g66639(.A (n_6967), .B (n_1356), .Y (n_2679));
AND2X1 g66649(.A (n_424), .B (g17646), .Y (n_1458));
NAND2X1 g66654(.A (g5817), .B (n_10950), .Y (n_6398));
NOR2X1 g66659(.A (g3873), .B (g3881), .Y (n_1440));
NOR2X1 g66663(.A (g6219), .B (g6227), .Y (n_1471));
NAND2X1 g66674(.A (n_3439), .B (n_659), .Y (n_780));
NAND2X1 g66682(.A (g17646), .B (g17607), .Y (n_779));
INVX1 g66353(.A (n_1230), .Y (n_778));
INVX1 g66711(.A (n_1538), .Y (n_777));
AND2X1 g66736(.A (n_776), .B (g17604), .Y (n_1484));
NOR2X1 g66759(.A (n_5941), .B (g2217), .Y (n_775));
INVX1 g66774(.A (n_771), .Y (n_772));
NOR2X1 g66784(.A (g1657), .B (n_5936), .Y (n_769));
INVX1 g66458(.A (n_10578), .Y (n_11217));
DFFSRX1 g4688_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g34028), .Q (), .QN (g4688));
NOR2X1 g66851(.A (n_10213), .B (n_11129), .Y (n_10206));
NOR2X1 g66867(.A (n_5932), .B (g2060), .Y (n_765));
AND2X1 g66870(.A (g25219), .B (g17577), .Y (n_1488));
NAND2X1 g66891(.A (g6163), .B (n_10949), .Y (n_6406));
NOR2X1 g66720(.A (g5873), .B (g5881), .Y (n_1455));
AND2X1 g66660(.A (n_11157), .B (g17685), .Y (n_1457));
INVX1 g66315(.A (n_747), .Y (n_748));
AND2X1 g62238(.A (n_746), .B (g13259), .Y (n_4754));
AND2X1 g62244(.A (n_745), .B (g13259), .Y (n_4757));
INVX1 g66292(.A (n_1370), .Y (n_744));
INVX1 g68093(.A (n_740), .Y (n_741));
INVX1 g66479(.A (n_1725), .Y (n_739));
NOR2X1 g66560(.A (n_730), .B (g2351), .Y (n_1059));
INVX2 g67032(.A (n_2421), .Y (n_2376));
DFFSRX1 g3661_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13926), .Q (g16744), .QN ());
OAI21X1 g61595(.A0 (g4401), .A1 (g4434), .B0 (n_243), .Y (n_724));
INVX1 g66918(.A (n_723), .Y (n_3042));
XOR2X1 g66077(.A (n_2280), .B (g_20563), .Y (n_722));
DFFSRX1 g5976_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17607), .Q (g17646), .QN ());
AOI21X1 g65984(.A0 (n_563), .A1 (g4311), .B0 (n_404), .Y (n_720));
INVX1 g68169(.A (n_719), .Y (n_1352));
INVX1 g66529(.A (n_1402), .Y (n_718));
XOR2X1 g66083(.A (n_716), .B (n_5958), .Y (n_717));
XOR2X1 g66079(.A (n_714), .B (n_5229), .Y (n_715));
INVX1 g66186(.A (n_10678), .Y (n_11221));
NOR2X1 g66508(.A (n_10213), .B (n_11187), .Y (n_10185));
OAI21X1 g65964(.A0 (n_2861), .A1 (n_3181), .B0 (g4473), .Y (n_709));
NOR2X1 g66863(.A (g5180), .B (g5188), .Y (n_1480));
OAI21X1 g65959(.A0 (g_10715), .A1 (n_708), .B0 (g_12791), .Y(n_1124));
NOR2X1 g66860(.A (g5527), .B (g5535), .Y (n_1476));
NOR2X1 g66746(.A (n_490), .B (n_11203), .Y (n_10809));
AND2X1 g66497(.A (n_730), .B (g2351), .Y (n_707));
NAND2X1 g65659(.A (n_1184), .B (n_1191), .Y (n_4314));
NOR2X1 g65762(.A (n_204), .B (n_7247), .Y (n_1219));
OR2X1 g62605(.A (g19334), .B (g7916), .Y (n_705));
INVX1 g66819(.A (n_1541), .Y (n_3323));
NAND2X1 g65728(.A (n_234), .B (n_2258), .Y (n_704));
INVX2 g68056(.A (n_2208), .Y (n_1023));
NAND2X1 g65717(.A (g2084), .B (n_7101), .Y (n_702));
NAND2X1 g65713(.A (n_745), .B (n_8796), .Y (n_698));
AND2X1 g66473(.A (n_806), .B (g1926), .Y (n_697));
XOR2X1 g65515(.A (g5084), .B (g5092), .Y (n_696));
AND2X1 g65515_and(.A (g5084), .B (g5092), .Y (n_1580));
XOR2X1 g65521(.A (g4258), .B (g4264), .Y (n_695));
AND2X1 g65521_and(.A (g4258), .B (g4264), .Y (n_1582));
XOR2X1 g65506(.A (n_11163), .B (g_20268), .Y (n_694));
AND2X1 g65506_and(.A (n_11163), .B (g_20268), .Y (n_693));
NOR2X1 g66394(.A (n_482), .B (g5188), .Y (n_1762));
NAND2X1 g66461(.A (g_21778), .B (n_691), .Y (n_692));
NAND2X1 g66435(.A (n_690), .B (g_3974), .Y (n_802));
INVX1 g68404(.A (n_10224), .Y (n_946));
XOR2X1 g66044(.A (g3827), .B (g3821), .Y (n_688));
DFFSRX1 g358_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8719), .Q (n_11116), .QN ());
OR2X1 g66493(.A (n_3789), .B (g1728), .Y (n_3948));
DFFSRX1 g4210_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8788), .Q (g8789), .QN ());
OR2X1 g66490(.A (n_804), .B (g1760), .Y (n_1236));
AND2X1 g66456(.A (n_11110), .B (g_21318), .Y (n_1024));
NAND2X1 g66417(.A (g5511), .B (n_686), .Y (n_983));
NOR2X1 g66811(.A (g4991), .B (n_684), .Y (n_685));
NOR2X1 g64908(.A (n_19), .B (g4688), .Y (n_680));
NOR2X1 g64915(.A (g4688), .B (n_294), .Y (n_1307));
NOR2X1 g66452(.A (n_6922), .B (g_20208), .Y (n_876));
NOR2X1 g66450(.A (g3857), .B (n_678), .Y (n_1181));
NOR2X1 g66437(.A (g1657), .B (n_677), .Y (g25167));
NOR2X1 g65879(.A (n_20), .B (n_988), .Y (n_676));
AND2X1 g66442(.A (n_674), .B (g2060), .Y (n_675));
AND2X1 g66387(.A (n_661), .B (g6573), .Y (n_1391));
DFFSRX1 g4405_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7243), .Q (g4405), .QN ());
INVX1 g66781(.A (n_673), .Y (n_1222));
DFFSRX1 g5623_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17711), .Q (g17580), .QN ());
DFFSRX1 g1333_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8475), .Q (g1333), .QN ());
DFFSRX1 g1459_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g19357), .Q (g13272), .QN ());
NAND2X1 g66418(.A (n_3943), .B (g1996), .Y (n_670));
DFFSRX1 g1236_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g10500), .Q (g1236), .QN ());
NAND2X1 g66427(.A (n_3943), .B (g2070), .Y (n_667));
AND2X1 g66347(.A (n_626), .B (g3881), .Y (n_1364));
OR2X1 g66425(.A (n_3943), .B (g1996), .Y (n_4318));
NOR2X1 g66423(.A (n_128), .B (n_6979), .Y (n_4682));
NAND2X1 g66313(.A (n_11160), .B (g_6165), .Y (n_818));
NOR2X1 g66448(.A (n_10197), .B (n_224), .Y (n_978));
NOR2X1 g66433(.A (g3506), .B (n_664), .Y (n_1201));
MX2X1 g66131(.A (g_21806), .B (g_19241), .S0 (g_20268), .Y (n_1290));
INVX1 g65516(.A (n_982), .Y (n_663));
DFFSRX1 g979_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13259), .Q (n_10125), .QN ());
NOR2X1 g66381(.A (n_661), .B (g6573), .Y (n_1718));
OAI21X1 g65629(.A0 (g6523), .A1 (g6537), .B0 (g35), .Y (n_1630));
DFFSRX1 g4308_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9251), .Q (g4308), .QN ());
DFFSRX1 g4474_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g4467), .Q (g4474), .QN ());
XOR2X1 g66165(.A (g4308), .B (g9251), .Y (n_1570));
XOR2X1 g66179(.A (g1548), .B (g1430), .Y (n_652));
NAND3X1 g65815(.A (n_50), .B (g1178), .C (g_20614), .Y (n_1636));
XOR2X1 g66175(.A (g_22600), .B (g_22371), .Y (n_650));
NAND3X1 g65845(.A (g1367), .B (g1379), .C (g1345), .Y (n_1276));
MX2X1 g61436(.A (g10527), .B (g12923), .S0 (g17423), .Y (n_649));
INVX1 g66800(.A (n_647), .Y (n_648));
INVX1 g66740(.A (n_10622), .Y (n_10180));
XOR2X1 g66053(.A (g8786), .B (n_10867), .Y (n_643));
DFFSRX1 g55_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_628), .Q (g55), .QN ());
INVX1 g66733(.A (n_4760), .Y (n_4791));
XOR2X1 g66074(.A (g5827), .B (g5821), .Y (n_639));
DFFSRX1 g6000_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17646), .Q (g13068), .QN ());
XOR2X1 g66076(.A (g3476), .B (g3470), .Y (n_638));
AOI22X1 g66088(.A0 (g2936), .A1 (g2941), .B0 (g2950), .B1 (g2955), .Y(n_637));
AOI22X1 g66089(.A0 (g_14342), .A1 (g_19414), .B0 (g_10715), .B1(g_12791), .Y (n_636));
OR2X1 g66378(.A (n_812), .B (g2453), .Y (n_1138));
OAI21X1 g61476(.A0 (g1395), .A1 (g1404), .B0 (g12923), .Y (n_635));
NAND2X1 g66455(.A (n_8587), .B (g_4050), .Y (n_800));
DFFSRX1 g990_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8416), .Q (g_15287), .QN ());
XOR2X1 g66164(.A (g4281), .B (g8839), .Y (n_1820));
XOR2X1 g66176(.A (g_14535), .B (g8358), .Y (n_1732));
NOR2X1 g66375(.A (g1636), .B (n_629), .Y (g25259));
DFFSRX1 g34_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(n_628), .Q (g_9174), .QN ());
DFFSRX1 g6711_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13099), .Q (g17871), .QN ());
DFFSRX1 g5112_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9553), .Q (), .QN (g5112));
DFFSRX1 g218_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8291), .Q (g_7220), .QN ());
DFFSRX1 g6019_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13068), .Q (g17819), .QN ());
DFFSRX1 g5327_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13039), .Q (g17787), .QN ());
DFFSRX1 g6365_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13085), .Q (g17845), .QN ());
AND2X1 g66373(.A (g5857), .B (n_627), .Y (n_1194));
DFFSRX1 g1579_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g10527), .Q (), .QN (g1579));
NOR2X1 g66712(.A (n_416), .B (n_251), .Y (n_1538));
AND2X1 g66371(.A (g6219), .B (n_617), .Y (n_1723));
NOR2X1 g66277(.A (n_626), .B (g3881), .Y (n_1743));
NOR2X1 g66278(.A (n_609), .B (g6395), .Y (n_3277));
NOR2X1 g66283(.A (n_674), .B (g2060), .Y (n_1515));
NAND2X1 g66285(.A (n_10369), .B (g_4409), .Y (n_823));
NOR2X1 g66293(.A (g3171), .B (n_553), .Y (n_1370));
NAND2X1 g66294(.A (n_6742), .B (g2629), .Y (n_624));
NOR2X1 g66307(.A (g3155), .B (n_623), .Y (n_1147));
NAND2X1 g66316(.A (g4608), .B (n_3624), .Y (n_747));
DFFSRX1 g6315_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17760), .Q (g17649), .QN ());
AND2X1 g66320(.A (g3506), .B (n_664), .Y (n_1207));
NAND2X1 g66333(.A (g5164), .B (n_621), .Y (n_817));
NOR2X1 g66336(.A (g5857), .B (n_627), .Y (n_1246));
AND2X1 g66345(.A (n_619), .B (g2217), .Y (n_620));
NAND2X1 g66346(.A (n_6742), .B (g2555), .Y (n_618));
OR2X1 g66354(.A (n_806), .B (g1894), .Y (n_1230));
NOR2X1 g66366(.A (n_11071), .B (n_134), .Y (n_2600));
NOR2X1 g66367(.A (g6219), .B (n_617), .Y (n_1377));
NOR2X1 g66368(.A (n_619), .B (g2217), .Y (n_1520));
AND2X1 g66382(.A (n_11165), .B (g_8864), .Y (n_1011));
AND2X1 g66384(.A (g3155), .B (n_623), .Y (n_1243));
AND2X1 g66385(.A (n_11071), .B (n_134), .Y (n_3275));
NOR2X1 g66389(.A (n_616), .B (g3530), .Y (n_1751));
AND2X1 g66407(.A (n_616), .B (g3530), .Y (n_1367));
XOR2X1 g66073(.A (g3125), .B (g3119), .Y (n_615));
AND2X1 g66424(.A (g6203), .B (n_612), .Y (n_1158));
AND2X1 g66428(.A (n_610), .B (g2619), .Y (n_611));
AND2X1 g66460(.A (n_609), .B (g6395), .Y (n_2325));
OR2X1 g66465(.A (n_4301), .B (g2153), .Y (n_4109));
AND2X1 g66469(.A (g1657), .B (n_677), .Y (n_608));
OR2X1 g66487(.A (n_3939), .B (g2421), .Y (n_4122));
NOR2X1 g66494(.A (n_8637), .B (n_10818), .Y (n_607));
AND2X1 g66507(.A (n_10197), .B (n_224), .Y (n_1179));
OR2X1 g66513(.A (g4608), .B (n_3624), .Y (n_1831));
NOR2X1 g66519(.A (n_610), .B (g2619), .Y (n_1506));
AND2X1 g66523(.A (g3857), .B (n_678), .Y (n_1185));
NOR2X1 g66531(.A (n_610), .B (g2587), .Y (n_1522));
OR2X1 g66532(.A (n_3782), .B (g1862), .Y (n_3945));
OR2X1 g66536(.A (g6549), .B (n_603), .Y (n_791));
NOR2X1 g66538(.A (g6203), .B (n_612), .Y (n_1149));
NOR2X1 g66551(.A (n_95), .B (g_17426), .Y (n_3391));
AND2X1 g66553(.A (n_455), .B (n_11198), .Y (n_11101));
XOR2X1 g66010(.A (g6519), .B (g6513), .Y (n_600));
OR2X1 g66357(.A (g1592), .B (n_347), .Y (n_3938));
NOR2X1 g66570(.A (n_598), .B (g4966), .Y (n_599));
AND2X1 g66571(.A (n_191), .B (n_10657), .Y (n_2597));
NAND2X1 g66572(.A (g4388), .B (n_596), .Y (n_597));
NAND2X1 g66573(.A (g4430), .B (n_596), .Y (n_595));
NAND2X1 g66575(.A (n_10139), .B (n_6967), .Y (n_1173));
AND2X1 g66577(.A (n_6979), .B (n_128), .Y (n_11128));
AND2X1 g66582(.A (n_401), .B (g_3381), .Y (n_1093));
INVX1 g66586(.A (n_1267), .Y (n_594));
INVX1 g66603(.A (n_1468), .Y (n_1143));
INVX1 g66605(.A (n_591), .Y (n_592));
NAND2X1 g66617(.A (n_627), .B (n_215), .Y (n_589));
NOR2X1 g66624(.A (n_413), .B (n_456), .Y (n_588));
NAND2X1 g66635(.A (n_603), .B (n_261), .Y (n_587));
INVX1 g66646(.A (n_1486), .Y (n_585));
NOR2X1 g66653(.A (n_10630), .B (n_10634), .Y (n_584));
INVX1 g66666(.A (n_908), .Y (n_581));
NAND2X1 g66675(.A (n_664), .B (n_365), .Y (n_580));
INVX1 g66708(.A (n_6790), .Y (n_579));
NAND2X1 g66717(.A (n_686), .B (n_383), .Y (n_578));
INVX1 g66722(.A (n_970), .Y (n_1224));
NOR2X1 g66350(.A (n_619), .B (g2185), .Y (n_1527));
NAND2X1 g66764(.A (n_678), .B (n_303), .Y (n_575));
NOR2X1 g66768(.A (n_10228), .B (n_10225), .Y (n_8778));
INVX1 g66770(.A (n_411), .Y (n_1264));
NOR2X1 g66775(.A (n_10139), .B (n_379), .Y (n_771));
NAND2X1 g66791(.A (n_572), .B (n_571), .Y (n_2111));
INVX1 g66794(.A (n_1145), .Y (n_1459));
INVX1 g66802(.A (n_1464), .Y (n_1227));
OR2X1 g66806(.A (g8475), .B (g7946), .Y (n_568));
NAND2X1 g66825(.A (n_612), .B (n_330), .Y (n_566));
NAND2X1 g66827(.A (n_623), .B (n_370), .Y (n_565));
NAND2X1 g66830(.A (n_563), .B (n_327), .Y (n_564));
INVX1 g66841(.A (n_561), .Y (n_562));
INVX1 g66854(.A (n_7101), .Y (n_558));
DFFSRX1 g1116_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g19334), .Q (g13259), .QN ());
INVX1 g66868(.A (n_7024), .Y (n_557));
OR2X1 g66874(.A (g19357), .B (g7946), .Y (n_556));
NOR2X1 g66889(.A (n_297), .B (n_406), .Y (n_3365));
AND2X1 g66343(.A (g3171), .B (n_553), .Y (n_1758));
INVX1 g66919(.A (n_552), .Y (n_723));
DFFSRX1 g1087_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17400), .Q (g_18330), .QN ());
DFFSRX1 g4878_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g34036), .Q (), .QN (g4878));
XOR2X1 g66001(.A (g5128), .B (g5134), .Y (n_540));
INVX1 g66664(.A (n_973), .Y (n_1154));
NOR2X1 g66311(.A (n_522), .B (g5535), .Y (n_1777));
DFFSRX1 g5654_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17604), .Q (g13049), .QN ());
NOR2X1 g66337(.A (g1389), .B (n_6782), .Y (n_3364));
DFFSRX1 g6012_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14738), .Q (g17739), .QN ());
DFFSRX1 g4871_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g34035), .Q (g34036), .QN ());
INVX1 g66669(.A (n_901), .Y (n_1212));
DFFSRX1 g5666_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14694), .Q (g17711), .QN ());
DFFSRX1 g1426_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17404), .Q (g17423), .QN ());
DFFSRX1 g5969_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17739), .Q (g17607), .QN ());
DFFSRX1 g6661_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17778), .Q (g17688), .QN ());
DFFSRX1 g5308_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17577), .Q (g13039), .QN ());
NAND2X1 g66329(.A (n_103), .B (n_11050), .Y (n_1100));
AND2X1 g66658(.A (n_523), .B (g6736), .Y (n_524));
AND2X1 g66325(.A (n_522), .B (g5535), .Y (n_1411));
NOR2X1 g66655(.A (n_8913), .B (n_10818), .Y (n_521));
INVX1 g68267(.A (n_10314), .Y (n_519));
MX2X1 g61555(.A (g10500), .B (g12919), .S0 (g17400), .Y (n_515));
DFFSRX1 g4411_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7257), .Q (g4411), .QN ());
DFFSRX1 g4452_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7245), .Q (g4452), .QN ());
INVX1 g67211(.A (g4584), .Y (n_3624));
NOR2X1 g66304(.A (n_512), .B (g4601), .Y (n_820));
DFFSRX1 g1242_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12919), .Q (), .QN (g1242));
OR2X1 g66301(.A (g5164), .B (n_621), .Y (n_822));
OR2X1 g66379(.A (g2984), .B (n_628), .Y (n_511));
NAND3X1 g65813(.A (g_22306), .B (g_12465), .C (g_19911), .Y (n_989));
OR2X1 g66290(.A (n_6742), .B (g2555), .Y (n_4118));
DFFSRX1 g1083_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17316), .Q (g17400), .QN ());
INVX1 g68012(.A (n_503), .Y (n_504));
INVX2 g68057(.A (n_776), .Y (n_2208));
DFFSRX1 g5673_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13049), .Q (g17813), .QN ());
INVX1 g68119(.A (n_10245), .Y (n_2177));
OAI21X1 g61586(.A0 (g_18488), .A1 (n_8508), .B0 (g12919), .Y (n_496));
INVX4 g67034(.A (n_546), .Y (n_2421));
CLKBUFX1 g68332(.A (n_490), .Y (n_4980));
AND2X1 g66569(.A (n_11038), .B (n_8807), .Y (n_2339));
INVX1 g66906(.A (n_896), .Y (n_1482));
NAND2X1 g66486(.A (n_453), .B (g_19172), .Y (n_799));
INVX1 g68244(.A (n_488), .Y (n_2017));
DFFSRX1 g4297_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g10122), .Q (g4297), .QN ());
DFFSRX1 g1422_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17320), .Q (g17404), .QN ());
OR2X1 g66506(.A (g5511), .B (n_686), .Y (n_795));
INVX1 g66872(.A (n_486), .Y (n_487));
INVX1 g68170(.A (g_20952), .Y (n_719));
AND2X1 g66530(.A (n_482), .B (g5188), .Y (n_1402));
DFFSRX1 g6346_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17685), .Q (g13085), .QN ());
AND2X1 g66526(.A (g6549), .B (n_603), .Y (n_1395));
OR2X1 g66521(.A (n_730), .B (g2319), .Y (n_1160));
NAND2X1 g66883(.A (n_621), .B (n_388), .Y (n_479));
DFFSRX1 g4291_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g9019), .Q (g4291), .QN ());
OR2X1 g66511(.A (n_4038), .B (g2287), .Y (n_4124));
INVX1 g66864(.A (n_4631), .Y (n_4679));
INVX1 g65512(.A (n_474), .Y (n_971));
DFFSRX1 g5276_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17674), .Q (g17519), .QN ());
DFFSRX1 g5320_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14662), .Q (g17674), .QN ());
DFFSRX1 g1322_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g13272), .Q (g1322), .QN ());
DFFSRX1 g4188_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g11447), .Q (g8783), .QN ());
DFFSRX1 g1430_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17423), .Q (g1430), .QN ());
DFFSRX1 g4194_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8783), .Q (g8784), .QN ());
DFFSRX1 g4200_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8785), .Q (g8786), .QN ());
DFFSRX1 g191_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8358), .Q (g_14535), .QN ());
DFFSRX1 g6358_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14779), .Q (g17760), .QN ());
DFFSRX1 g1585_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g12923), .Q (), .QN (g1585));
NAND3X1 g65763(.A (g_10715), .B (g_15740), .C (g_12791), .Y (n_471));
XOR2X1 g66064(.A (g4388), .B (g4430), .Y (n_470));
XOR2X1 g66167(.A (n_10128), .B (g_18330), .Y (n_469));
INVX2 g66848(.A (n_10426), .Y (n_3459));
DFFSRX1 g1079_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17291), .Q (g17316), .QN ());
DFFSRX1 g4443_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g7260), .Q (g4443), .QN ());
NOR2X1 g66491(.A (n_674), .B (g2028), .Y (n_1524));
DFFSRX1 g6692_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g17722), .Q (g13099), .QN ());
INVX1 g68094(.A (n_10213), .Y (n_740));
DFFSRX1 g4281_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8839), .Q (g4281), .QN ());
INVX1 g67943(.A (n_464), .Y (g11349));
NOR2X1 g66488(.A (g1624), .B (n_677), .Y (n_1531));
INVX1 g66600(.A (n_1199), .Y (n_463));
XOR2X1 g66162(.A (g4291), .B (g9019), .Y (n_1556));
AND2X1 g66580(.A (n_459), .B (g5881), .Y (n_1382));
NAND2X1 g61309(.A (g1521), .B (n_460), .Y (n_461));
NOR2X1 g66480(.A (n_459), .B (g5881), .Y (n_1725));
INVX1 g66815(.A (n_1175), .Y (n_458));
DFFSRX1 g4197_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8784), .Q (g8785), .QN ());
DFFSRX1 g4204_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8786), .Q (g8787), .QN ());
CLKBUFX1 g66820(.A (n_6762), .Y (n_1541));
DFFSRX1 g4180_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8789), .Q (n_10871), .QN ());
NAND2X1 g66475(.A (g1442), .B (n_412), .Y (n_1729));
DFFSRX1 g4207_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g8787), .Q (g8788), .QN ());
INVX1 g68017(.A (n_1285), .Y (n_456));
INVX1 g67958(.A (n_2150), .Y (n_1540));
DFFSRX1 g6704_reg(.RN (n_6421), .SN (1'b1), .CK (blif_clk_net), .D(g14828), .Q (g17778), .QN ());
NOR2X1 g66552(.A (n_455), .B (n_11198), .Y (n_10508));
INVX1 g68333(.A (n_455), .Y (n_490));
NOR2X1 g66641(.A (g6336), .B (g6395), .Y (n_2413));
NOR2X1 g66809(.A (g2098), .B (g1964), .Y (n_442));
INVX1 g68245(.A (g_20951), .Y (n_488));
NOR2X1 g66805(.A (g1894), .B (g1926), .Y (n_441));
NAND2X1 g66804(.A (g_18330), .B (n_10128), .Y (n_474));
NAND2X1 g66801(.A (g1894), .B (g1926), .Y (n_647));
OR2X1 g66786(.A (g2537), .B (g2417), .Y (n_436));
AND2X1 g66816(.A (g3857), .B (g3863), .Y (n_1175));
INVX1 g67902(.A (g34034), .Y (n_477));
NAND2X1 g66760(.A (g1548), .B (g1430), .Y (n_982));
OR2X1 g66778(.A (g2338), .B (g2491), .Y (n_429));
NOR2X1 g66730(.A (g1844), .B (g1710), .Y (n_428));
INVX1 g68229(.A (n_6782), .Y (n_1275));
NOR2X1 g66885(.A (n_11071), .B (g6741), .Y (n_2435));
NOR2X1 g66792(.A (g2126), .B (g1992), .Y (n_425));
INVX1 g61358(.A (n_460), .Y (n_2474));
INVX1 g67026(.A (n_423), .Y (n_424));
INVX1 g67975(.A (n_417), .Y (n_659));
AND2X1 g66795(.A (g5857), .B (g5863), .Y (n_1145));
OR2X1 g61462(.A (g1404), .B (g12923), .Y (n_415));
NAND2X1 g66771(.A (g6219), .B (g6227), .Y (n_411));
INVX2 g67915(.A (n_690), .Y (n_5402));
INVX1 g67886(.A (g12238), .Y (n_465));
INVX1 g67798(.A (n_409), .Y (g12300));
NOR2X1 g66696(.A (g2453), .B (g2485), .Y (n_408));
INVX1 g67783(.A (n_6922), .Y (n_5663));
AND2X1 g66796(.A (g3873), .B (g3881), .Y (n_1184));
INVX1 g68058(.A (n_401), .Y (n_776));
NOR2X1 g65890(.A (g34035), .B (g34036), .Y (n_1578));
AND2X1 g66731(.A (g6336), .B (g6395), .Y (n_2352));
NOR2X1 g66728(.A (g2319), .B (g2351), .Y (n_376));
INVX1 g67169(.A (g17688), .Y (n_538));
NAND2X1 g66716(.A (g5124), .B (g35), .Y (n_3641));
AND2X1 g66718(.A (n_10660), .B (g5698), .Y (n_374));
INVX1 g67984(.A (n_367), .Y (n_2252));
INVX1 g68445(.A (g12422), .Y (n_660));
INVX1 g67009(.A (g17580), .Y (n_669));
NOR2X1 g66721(.A (g1664), .B (g1644), .Y (n_353));
AND2X1 g66723(.A (g5180), .B (g5188), .Y (n_970));
NAND2X1 g66724(.A (g4467), .B (g4473), .Y (n_1353));
NOR2X1 g66584(.A (g4141), .B (g4082), .Y (n_1312));
NOR2X1 g66587(.A (g4311), .B (n_662), .Y (n_1267));
NOR2X1 g66597(.A (g8787), .B (g8786), .Y (n_344));
AND2X1 g66907(.A (g3155), .B (g3161), .Y (n_896));
NOR2X1 g66620(.A (g6177), .B (g6191), .Y (n_343));
NAND2X1 g66627(.A (g2629), .B (g2555), .Y (n_342));
AND2X1 g66629(.A (n_10657), .B (g5644), .Y (n_2443));
AND2X1 g66902(.A (n_7247), .B (g4621), .Y (n_948));
NOR2X1 g66657(.A (g2685), .B (g2551), .Y (n_340));
AND2X1 g66673(.A (g2185), .B (g2217), .Y (n_1517));
AND2X1 g66686(.A (g6395), .B (g6390), .Y (n_339));
AND2X1 g66692(.A (g6509), .B (g35), .Y (n_3812));
NOR2X1 g66739(.A (g1624), .B (g1657), .Y (n_338));
NOR2X1 g66754(.A (g2587), .B (g2619), .Y (n_336));
NAND2X1 g66803(.A (g5164), .B (g5170), .Y (n_1464));
AND2X1 g66813(.A (n_11071), .B (g6741), .Y (n_2432));
NOR2X1 g66834(.A (g2066), .B (g2047), .Y (n_335));
OR2X1 g66838(.A (g7260), .B (g7245), .Y (n_334));
NAND2X1 g66842(.A (g1760), .B (g1792), .Y (n_561));
INVX1 g68439(.A (g11418), .Y (n_491));
AND2X1 g66873(.A (g2453), .B (g2485), .Y (n_486));
NOR2X1 g66886(.A (g1183), .B (n_8769), .Y (n_746));
AND2X1 g66699(.A (g3171), .B (g3179), .Y (n_1242));
INVX2 g67035(.A (n_423), .Y (n_546));
AND2X1 g66742(.A (g5873), .B (g5881), .Y (n_1245));
NOR2X1 g66725(.A (n_10657), .B (g5644), .Y (n_2439));
AND2X1 g66665(.A (g5527), .B (g5535), .Y (n_973));
OR2X1 g61584(.A (n_8508), .B (g12919), .Y (n_325));
AND2X1 g66670(.A (g3115), .B (g35), .Y (n_901));
NOR2X1 g66702(.A (g1760), .B (g1792), .Y (n_323));
INVX1 g68290(.A (n_322), .Y (g12470));
OR2X1 g66824(.A (g7257), .B (g7243), .Y (n_316));
NOR2X1 g66808(.A (g4153), .B (g4172), .Y (n_311));
OR2X1 g66652(.A (g17404), .B (g17320), .Y (n_309));
INVX1 g68232(.A (n_307), .Y (n_518));
NAND2X1 g66647(.A (g6549), .B (g6555), .Y (n_1486));
NOR2X1 g66871(.A (g4054), .B (g3990), .Y (n_4988));
OR2X1 g66861(.A (g1978), .B (g1858), .Y (n_302));
OR2X1 g66630(.A (g1779), .B (g1932), .Y (n_298));
OR2X1 g66831(.A (g17316), .B (g17291), .Y (n_295));
NAND2X1 g66881(.A (g2070), .B (g1996), .Y (n_290));
AND2X1 g66615(.A (g6565), .B (g6573), .Y (n_590));
NAND2X1 g66604(.A (g6203), .B (g6209), .Y (n_1468));
AND2X1 g66601(.A (g3506), .B (g3512), .Y (n_1199));
NAND2X1 g66782(.A (g5511), .B (g5517), .Y (n_673));
NAND2X1 g66691(.A (g5037), .B (g5033), .Y (n_281));
INVX1 g68274(.A (n_598), .Y (n_653));
INVX4 g68390(.A (g7946), .Y (n_3849));
AND2X1 g66772(.A (n_11201), .B (g6044), .Y (n_268));
INVX1 g66986(.A (g17649), .Y (n_549));
INVX1 g66943(.A (n_684), .Y (n_551));
INVX1 g68184(.A (n_276), .Y (n_3181));
NOR2X1 g66908(.A (g2403), .B (g2269), .Y (n_248));
INVX2 g66920(.A (n_10634), .Y (n_552));
NAND2X1 g61629(.A (g4401), .B (g4434), .Y (n_243));
NOR2X1 g66901(.A (g1830), .B (g1696), .Y (n_241));
NOR2X1 g66895(.A (g2028), .B (g2060), .Y (n_240));
NOR2X1 g66896(.A (g_20073), .B (g_12433), .Y (n_891));
INVX1 g68324(.A (g13966), .Y (n_493));
AND2X1 g66690(.A (g3522), .B (g3530), .Y (n_1206));
NOR2X1 g66890(.A (g2625), .B (g2606), .Y (n_235));
NAND2X1 g66880(.A (g5471), .B (g35), .Y (n_6399));
NOR2X1 g66887(.A (g2185), .B (g2217), .Y (n_234));
AND2X1 g66748(.A (g1183), .B (n_8769), .Y (n_745));
INVX1 g67875(.A (g17519), .Y (n_527));
INVX1 g68277(.A (n_1627), .Y (n_227));
INVX1 g68158(.A (n_691), .Y (n_3550));
INVX1 g68147(.A (n_224), .Y (n_2773));
INVX1 g68142(.A (n_223), .Y (n_3439));
NOR2X1 g66875(.A (n_10197), .B (g1526), .Y (n_899));
NOR2X1 g66866(.A (g1442), .B (g1489), .Y (n_4631));
AND2X1 g66857(.A (n_6979), .B (g3639), .Y (n_6973));
OR2X1 g66839(.A (g11447), .B (g8789), .Y (n_220));
NAND2X1 g66862(.A (g4669), .B (g4653), .Y (n_218));
AND2X1 g66667(.A (n_10197), .B (g1526), .Y (n_908));
AND2X1 g66651(.A (g1322), .B (g1404), .Y (n_1165));
NOR2X1 g66735(.A (g_18902), .B (g_19172), .Y (n_4760));
INVX1 g67944(.A (g_4050), .Y (n_464));
NAND2X1 g66694(.A (g4146), .B (g4157), .Y (n_209));
NOR2X1 g66648(.A (n_6958), .B (g_21651), .Y (n_205));
NAND2X1 g66845(.A (g4621), .B (g4633), .Y (n_204));
NOR2X1 g66783(.A (g5046), .B (g5052), .Y (n_196));
NOR2X1 g66835(.A (g2223), .B (g2204), .Y (n_194));
AND2X1 g66606(.A (g2319), .B (g2351), .Y (n_591));
INVX1 g67208(.A (n_191), .Y (n_4982));
NOR2X1 g66833(.A (g4087), .B (g4098), .Y (n_188));
AND2X1 g66828(.A (n_8509), .B (n_10125), .Y (n_8796));
INVX1 g68344(.A (n_8637), .Y (n_644));
INVX1 g68013(.A (n_10630), .Y (n_503));
CLKBUFX1 g67959(.A (n_8594), .Y (n_2150));
INVX1 g67122(.A (g2667), .Y (n_716));
INVX1 g68456(.A (g_16464), .Y (n_172));
INVX1 g66913(.A (n_3604), .Y (n_247));
INVX1 g67920(.A (g2040), .Y (n_3943));
INVX1 g67195(.A (g2295), .Y (n_1702));
INVX1 g68291(.A (g_8864), .Y (n_322));
INVX1 g68248(.A (g1959), .Y (n_836));
INVX1 g68114(.A (g2250), .Y (n_382));
INVX1 g68367(.A (g2303), .Y (n_1703));
INVX1 g68214(.A (g2704), .Y (n_169));
INVX1 g67742(.A (g5134), .Y (n_168));
INVX1 g68315(.A (g3133), .Y (n_2686));
INVX1 g68117(.A (g3490), .Y (n_1799));
INVX1 g67182(.A (g4653), .Y (n_294));
INVX1 g68211(.A (g4849), .Y (n_165));
INVX1 g67827(.A (g2856), .Y (n_3499));
INVX1 g68217(.A (g2177), .Y (n_919));
INVX1 g68338(.A (n_640), .Y (n_273));
INVX1 g68190(.A (g3147), .Y (n_3253));
INVX1 g67177(.A (g4462), .Y (n_2861));
CLKBUFX1 g68440(.A (g_3974), .Y (g11418));
INVX1 g66950(.A (g_20909), .Y (n_6324));
INVX1 g66955(.A (g2246), .Y (n_4906));
INVX1 g68353(.A (g2988), .Y (n_162));
INVX1 g68354(.A (g1564), .Y (n_1295));
INVX1 g68086(.A (n_3611), .Y (n_202));
INVX1 g67830(.A (g2571), .Y (n_362));
INVX1 g67126(.A (g6519), .Y (n_158));
INVX1 g68357(.A (g5517), .Y (n_686));
INVX1 g67846(.A (g2472), .Y (n_157));
INVX1 g68166(.A (g2527), .Y (n_5229));
INVX1 g68213(.A (g_18112), .Y (n_153));
INVX1 g67039(.A (g2864), .Y (n_271));
INVX1 g67752(.A (g13926), .Y (n_242));
INVX1 g68377(.A (g2898), .Y (n_3501));
INVX1 g67862(.A (g6555), .Y (n_603));
INVX1 g67747(.A (g1834), .Y (n_4948));
INVX1 g68327(.A (g2399), .Y (n_846));
INVX1 g68308(.A (g4035), .Y (n_151));
INVX1 g68254(.A (g4239), .Y (n_150));
INVX1 g67025(.A (g5170), .Y (n_621));
INVX1 g67093(.A (n_1234), .Y (n_383));
INVX1 g66916(.A (g1882), .Y (n_2306));
INVX1 g67012(.A (g2380), .Y (n_4529));
INVX1 g68263(.A (g2315), .Y (n_1677));
INVX1 g67925(.A (g2016), .Y (n_926));
INVX1 g68104(.A (g2384), .Y (n_831));
INVX1 g66997(.A (g5503), .Y (n_2943));
INVX1 g68394(.A (g2122), .Y (n_860));
INVX1 g67989(.A (g2648), .Y (n_4726));
INVX1 g68048(.A (g5406), .Y (n_144));
CLKBUFX1 g67842(.A (g6741), .Y (n_523));
INVX1 g67096(.A (g4659), .Y (n_143));
INVX1 g66970(.A (g2563), .Y (n_380));
INVX1 g68154(.A (g4515), .Y (n_563));
INVX1 g67209(.A (g5644), .Y (n_191));
INVX1 g67203(.A (g2197), .Y (n_4301));
INVX1 g67980(.A (g5849), .Y (n_2940));
INVX1 g67869(.A (g3139), .Y (n_1805));
INVX1 g68298(.A (g4382), .Y (n_5363));
INVX1 g67818(.A (g4593), .Y (n_512));
INVX1 g66962(.A (g2116), .Y (n_6017));
INVX1 g68198(.A (n_2005), .Y (n_412));
INVX1 g67215(.A (g1768), .Y (n_136));
INVX1 g68317(.A (g2643), .Y (n_902));
INVX1 g67099(.A (g1714), .Y (n_6027));
INVX1 g68261(.A (g3841), .Y (n_1796));
INVX1 g66959(.A (n_3589), .Y (n_332));
INVX1 g67864(.A (g1454), .Y (n_2538));
INVX1 g68078(.A (g3684), .Y (n_1818));
INVX1 g67843(.A (g6741), .Y (n_134));
INVX1 g67790(.A (g13895), .Y (n_238));
INVX1 g68365(.A (g2449), .Y (n_1671));
INVX1 g66262(.A (g34027), .Y (n_988));
INVX1 g67966(.A (g2008), .Y (n_1514));
INVX1 g68436(.A (g1848), .Y (n_5978));
INVX1 g67108(.A (g2012), .Y (n_368));
INVX1 g67155(.A (n_5936), .Y (n_677));
INVX1 g68016(.A (g1706), .Y (n_856));
INVX1 g68084(.A (g2361), .Y (n_386));
INVX1 g66980(.A (n_5928), .Y (n_610));
INVX1 g67871(.A (g2279), .Y (n_975));
INVX1 g68124(.A (g2024), .Y (n_278));
INVX1 g67780(.A (g3522), .Y (n_616));
INVX1 g68305(.A (g1982), .Y (n_5975));
INVX1 g68304(.A (g2020), .Y (n_399));
INVX1 g67103(.A (g2407), .Y (n_5972));
INVX1 g67083(.A (g_18488), .Y (n_129));
INVX1 g68260(.A (g1604), .Y (n_1509));
INVX1 g61359(.A (g1339), .Y (n_460));
INVX1 g67991(.A (g2413), .Y (n_866));
INVX1 g68027(.A (g3639), .Y (n_128));
INVX1 g67976(.A (g_16475), .Y (n_417));
INVX1 g67097(.A (g6098), .Y (n_127));
INVX1 g68165(.A (g6565), .Y (n_661));
INVX1 g66914(.A (g5863), .Y (n_627));
INVX1 g68143(.A (g_15016), .Y (n_223));
INVX1 g68296(.A (g20899), .Y (n_2518));
INVX1 g68074(.A (g2917), .Y (n_3463));
INVX1 g67897(.A (n_3616), .Y (n_356));
INVX1 g67930(.A (g_16958), .Y (n_416));
INVX1 g68180(.A (g4601), .Y (n_262));
CLKBUFX1 g68031(.A (g6336), .Y (n_4978));
INVX1 g67753(.A (g_19414), .Y (n_126));
INVX1 g67006(.A (g2681), .Y (n_852));
INVX1 g66991(.A (g6173), .Y (n_125));
INVX1 g67824(.A (g6181), .Y (n_2704));
INVX1 g68415(.A (g6527), .Y (n_3007));
INVX1 g68102(.A (g2145), .Y (n_308));
INVX1 g67934(.A (g2004), .Y (n_450));
INVX1 g68041(.A (g_12791), .Y (n_413));
INVX1 g67148(.A (g_22306), .Y (n_286));
INVX1 g66978(.A (n_1214), .Y (n_330));
INVX1 g67956(.A (g6195), .Y (n_2936));
INVX1 g68209(.A (g1906), .Y (n_3782));
INVX1 g68173(.A (g6209), .Y (n_612));
INVX1 g67014(.A (g2299), .Y (n_1676));
INVX1 g68116(.A (g1437), .Y (n_2535));
INVX1 g66941(.A (n_4339), .Y (n_437));
INVX1 g66938(.A (g2181), .Y (n_1519));
INVX1 g68236(.A (n_5921), .Y (n_812));
INVX1 g67811(.A (g2138), .Y (n_1240));
INVX1 g68408(.A (g1691), .Y (n_187));
INVX1 g67765(.A (g6541), .Y (n_2930));
INVX1 g68225(.A (g3498), .Y (n_2928));
INVX1 g68363(.A (g_21447), .Y (n_3310));
INVX1 g67200(.A (g2771), .Y (n_326));
INVX1 g67806(.A (g1608), .Y (n_1533));
INVX1 g67171(.A (g3161), .Y (n_623));
INVX1 g68196(.A (g1600), .Y (n_1532));
INVX1 g68362(.A (g2533), .Y (n_714));
INVX1 g67756(.A (g3457), .Y (n_3601));
INVX1 g67088(.A (g_20839), .Y (n_2280));
INVX1 g68370(.A (g2583), .Y (n_213));
INVX1 g68201(.A (g4076), .Y (n_118));
INVX1 g67011(.A (g3752), .Y (n_117));
INVX1 g68360(.A (g1379), .Y (n_263));
INVX1 g66935(.A (g2331), .Y (n_4038));
INVX1 g67891(.A (g55), .Y (n_628));
INVX1 g67150(.A (g5873), .Y (n_459));
INVX1 g67949(.A (g1467), .Y (n_2485));
INVX1 g67218(.A (g2429), .Y (n_1713));
INVX1 g68218(.A (g5835), .Y (n_2684));
INVX1 g68334(.A (g5990), .Y (n_455));
INVX1 g68109(.A (n_3618), .Y (n_389));
INVX1 g68282(.A (g1720), .Y (n_878));
INVX1 g66964(.A (g3808), .Y (n_3596));
INVX1 g68233(.A (g1221), .Y (n_307));
INVX1 g68356(.A (g5527), .Y (n_522));
INVX1 g67812(.A (g4843), .Y (n_1274));
INVX1 g68379(.A (n_2458), .Y (n_397));
INVX1 g66925(.A (g_20159), .Y (n_251));
INVX2 g67916(.A (g4040), .Y (n_690));
INVX1 g67884(.A (g5057), .Y (n_110));
INVX1 g67947(.A (g1322), .Y (n_1502));
INVX1 g67939(.A (n_1169), .Y (n_215));
INVX1 g68189(.A (g2227), .Y (n_259));
INVX1 g66956(.A (g9553), .Y (n_107));
INVX1 g67023(.A (g1632), .Y (n_105));
INVX1 g68148(.A (g1526), .Y (n_224));
INVX1 g67037(.A (g6035), .Y (n_103));
INVX1 g66998(.A (g2089), .Y (n_4183));
INVX1 g68130(.A (g2108), .Y (n_862));
INVX1 g68152(.A (g20763), .Y (n_101));
INVX1 g68220(.A (g1616), .Y (n_928));
INVX1 g68286(.A (g4392), .Y (n_596));
INVX1 g66932(.A (g2941), .Y (n_98));
INVX1 g68453(.A (n_662), .Y (n_404));
INVX1 g68458(.A (g1612), .Y (n_2521));
INVX1 g67791(.A (g1484), .Y (n_3383));
INVX1 g68237(.A (g1968), .Y (n_4946));
INVX1 g67844(.A (g_16063), .Y (n_3914));
INVX1 g67165(.A (n_4120), .Y (n_629));
INVX1 g67803(.A (g2437), .Y (n_1714));
INVX1 g67942(.A (g2193), .Y (n_96));
INVX1 g67950(.A (g3484), .Y (n_2699));
INVX1 g68421(.A (g1752), .Y (n_444));
INVX1 g68144(.A (g_10278), .Y (n_95));
INVX1 g67833(.A (g5481), .Y (n_94));
INVX1 g67743(.A (g4483), .Y (n_93));
INVX1 g67941(.A (g1736), .Y (n_1710));
INVX1 g67216(.A (g1236), .Y (n_92));
INVX1 g67836(.A (g2311), .Y (n_377));
INVX1 g66996(.A (g4486), .Y (n_89));
INVX1 g67982(.A (g_16769), .Y (n_2290));
INVX1 g66982(.A (g_9176), .Y (n_6057));
INVX1 g68112(.A (g1554), .Y (n_392));
INVX1 g68125(.A (g2273), .Y (n_6025));
INVX1 g67098(.A (g5752), .Y (n_87));
INVX1 g67080(.A (g_4449), .Y (n_284));
INVX1 g67120(.A (g_15879), .Y (n_86));
INVX1 g66954(.A (g_10715), .Y (n_2583));
INVX1 g67102(.A (g1840), .Y (n_854));
CLKBUFX1 g66944(.A (g4966), .Y (n_684));
INVX1 g66917(.A (g5495), .Y (n_1810));
INVX1 g67758(.A (g3827), .Y (n_85));
INVX1 g68412(.A (g3835), .Y (n_2692));
INVX1 g67145(.A (g_12465), .Y (n_287));
INVX1 g67997(.A (blif_reset_net), .Y (n_6421));
INVX1 g67153(.A (g4057), .Y (n_571));
INVX1 g67776(.A (g2575), .Y (n_933));
INVX1 g67750(.A (g_22464), .Y (n_83));
INVX1 g68417(.A (g2093), .Y (n_433));
INVX1 g67187(.A (g_16571), .Y (n_364));
INVX1 g67084(.A (g2675), .Y (n_6020));
INVX1 g68423(.A (g2433), .Y (n_1670));
INVX1 g67176(.A (g1886), .Y (n_291));
INVX1 g67928(.A (n_2429), .Y (n_453));
INVX1 g68224(.A (g1988), .Y (n_885));
INVX1 g67764(.A (g6187), .Y (n_2084));
INVX1 g68090(.A (g_15381), .Y (n_79));
INVX1 g67094(.A (g_22236), .Y (n_2529));
INVX1 g68322(.A (g1854), .Y (n_883));
INVX1 g66966(.A (g1874), .Y (n_1687));
INVX1 g67183(.A (g2514), .Y (n_4531));
INVX1 g66994(.A (g2465), .Y (n_3939));
INVX1 g67087(.A (g4116), .Y (n_282));
INVX1 g67986(.A (g1536), .Y (n_367));
INVX1 g68043(.A (g2652), .Y (n_418));
INVX1 g67754(.A (g2541), .Y (n_5969));
INVX1 g68132(.A (g1870), .Y (n_1705));
INVX1 g68181(.A (g4093), .Y (n_955));
INVX1 g67823(.A (g5909), .Y (n_75));
INVX1 g68081(.A (g2445), .Y (n_269));
INVX1 g67795(.A (g4417), .Y (n_74));
INVX1 g68099(.A (g1878), .Y (n_1706));
INVX1 g68381(.A (g3873), .Y (n_626));
INVX1 g68091(.A (g3106), .Y (n_3609));
INVX1 g68352(.A (g4311), .Y (n_327));
INVX1 g67788(.A (g2567), .Y (n_1505));
INVX1 g67040(.A (g3512), .Y (n_664));
INVX1 g67808(.A (g_22600), .Y (n_70));
INVX1 g65203(.A (g4688), .Y (n_69));
INVX1 g67142(.A (g1902), .Y (n_67));
INVX1 g68060(.A (g_18220), .Y (n_2556));
INVX1 g67119(.A (g3849), .Y (n_2923));
INVX1 g67900(.A (n_4139), .Y (n_446));
INVX1 g68163(.A (n_5996), .Y (n_804));
INVX1 g68077(.A (g5827), .Y (n_65));
INVX1 g67019(.A (n_5941), .Y (n_619));
INVX1 g68159(.A (g_20268), .Y (n_691));
INVX1 g67077(.A (g3333), .Y (n_64));
INVX1 g68314(.A (g_10556), .Y (n_447));
INVX1 g68372(.A (g2518), .Y (n_839));
INVX1 g68411(.A (g6227), .Y (n_617));
INVX1 g68135(.A (g2375), .Y (n_911));
INVX1 g67963(.A (g1772), .Y (n_3789));
INVX1 g67799(.A (g_3381), .Y (n_409));
INVX1 g68222(.A (g2509), .Y (n_904));
INVX1 g68292(.A (g3476), .Y (n_60));
INVX1 g67895(.A (g3401), .Y (n_59));
INVX1 g67978(.A (g2165), .Y (n_1518));
INVX1 g66947(.A (g_18200), .Y (n_2244));
INVX2 g68275(.A (g4983), .Y (n_598));
INVX1 g66929(.A (n_5917), .Y (n_730));
INVX1 g67196(.A (g2327), .Y (n_57));
INVX1 g68358(.A (g2441), .Y (n_2780));
INVX1 g67021(.A (g2393), .Y (n_4942));
INVX1 g67894(.A (g5180), .Y (n_482));
INVX1 g67860(.A (n_5932), .Y (n_674));
INVX1 g68256(.A (g2036), .Y (n_54));
INVX1 g67111(.A (g3179), .Y (n_553));
INVX1 g68294(.A (g2595), .Y (n_52));
INVX1 g67017(.A (g1936), .Y (n_328));
INVX1 g67774(.A (g1756), .Y (n_1666));
INVX1 g66967(.A (g2173), .Y (n_2258));
INVX1 g67190(.A (g1189), .Y (n_50));
INVX1 g67786(.A (g_16792), .Y (n_10496));
INVX1 g67141(.A (n_5925), .Y (n_806));
INVX1 g67146(.A (g1682), .Y (n_4893));
INVX1 g67979(.A (g1687), .Y (n_4527));
INVX1 g67761(.A (g1636), .Y (n_347));
INVX1 g67105(.A (g4628), .Y (n_46));
INVX1 g67745(.A (g1373), .Y (n_406));
INVX1 g68375(.A (g2265), .Y (n_864));
INVX1 g67160(.A (g_5342), .Y (n_6331));
INVX1 g68383(.A (g2547), .Y (n_858));
INVX1 g67800(.A (g_18590), .Y (n_6252));
INVX1 g68312(.A (g4054), .Y (n_3769));
INVX1 g68320(.A (g4176), .Y (n_43));
INVX1 g67162(.A (g2169), .Y (n_1529));
INVX1 g67188(.A (g3863), .Y (n_678));
INVX1 g68030(.A (g1974), .Y (n_871));
INVX1 g67178(.A (g_6283), .Y (n_40));
INVX1 g66931(.A (g3050), .Y (n_39));
INVX1 g68293(.A (g2848), .Y (n_38));
INVX1 g68264(.A (g_14587), .Y (n_35));
INVX1 g67820(.A (g4119), .Y (n_360));
INVX1 g66953(.A (g2902), .Y (n_3765));
INVX1 g68206(.A (n_1191), .Y (n_303));
INVX1 g67057(.A (g34026), .Y (n_986));
INVX1 g68176(.A (g4112), .Y (n_245));
INVX1 g67970(.A (g5011), .Y (n_843));
INVX1 g67118(.A (n_1177), .Y (n_388));
INVX1 g66990(.A (g2579), .Y (n_351));
INVX1 g67112(.A (g_15801), .Y (n_32));
INVX1 g68194(.A (g_12276), .Y (n_30));
INVX1 g68160(.A (g1724), .Y (n_29));
INVX1 g67822(.A (g1620), .Y (n_1510));
INVX1 g67946(.A (g_22639), .Y (n_28));
INVX1 g67868(.A (g2803), .Y (n_317));
INVX1 g68418(.A (g1821), .Y (n_4190));
INVX1 g67763(.A (g2999), .Y (n_27));
INVX1 g68347(.A (g1744), .Y (n_1711));
INVX1 g67782(.A (g1740), .Y (n_1665));
INVX1 g68026(.A (g1395), .Y (n_26));
INVX1 g68149(.A (g4122), .Y (n_3135));
INVX1 g67159(.A (g17607), .Y (n_371));
INVX1 g67851(.A (n_1135), .Y (n_370));
INVX1 g67193(.A (n_1356), .Y (n_379));
INVX1 g67794(.A (g2259), .Y (n_5961));
INVX1 g68155(.A (g4621), .Y (n_23));
INVX1 g67741(.A (g_15740), .Y (n_708));
INVX1 g66972(.A (g1890), .Y (n_1688));
INVX1 g66961(.A (g23002), .Y (n_22));
INVX1 g67206(.A (g1361), .Y (n_297));
INVX1 g67883(.A (g4349), .Y (n_221));
INVX1 g67062(.A (g2102), .Y (n_5953));
CLKBUFX1 g67887(.A (g_4409), .Y (g12238));
INVX1 g67214(.A (g_13838), .Y (n_21));
INVX1 g68402(.A (g4821), .Y (n_20));
INVX1 g68258(.A (g4826), .Y (n_19));
INVX1 g68376(.A (g4831), .Y (n_1299));
INVX1 g68457(.A (g2307), .Y (n_2293));
INVX1 g67757(.A (g21292), .Y (g23612));
INVX1 g68414(.A (g2241), .Y (n_916));
INVX1 g67138(.A (g1913), .Y (n_17));
INVX1 g66910(.A (g1413), .Y (n_16));
INVX1 g67004(.A (g4489), .Y (n_13));
INVX1 g68107(.A (g2161), .Y (n_1528));
INVX1 g67804(.A (g1955), .Y (n_4187));
INVX1 g67926(.A (g2461), .Y (n_12));
INVX1 g67826(.A (g2735), .Y (n_11));
INVX1 g68059(.A (g5689), .Y (n_401));
INVX1 g67918(.A (g2661), .Y (n_5958));
INVX1 g67988(.A (g_5450), .Y (n_2566));
INVX1 g67772(.A (g4332), .Y (n_448));
INVX1 g65604(.A (g34028), .Y (n_987));
INVX2 g67036(.A (g6035), .Y (n_423));
INVX1 g68097(.A (g5489), .Y (n_3011));
INVX1 g67837(.A (g1748), .Y (n_2550));
INVX1 g68133(.A (g2283), .Y (n_5));
INVX1 g68136(.A (g6533), .Y (n_1794));
INVX1 g67055(.A (g5841), .Y (n_1807));
INVX1 g67003(.A (n_1216), .Y (n_261));
INVX1 g67996(.A (n_1210), .Y (n_365));
INVX1 g67024(.A (g5142), .Y (n_2718));
INVX1 g68139(.A (g4064), .Y (n_572));
INVX1 g68128(.A (g1700), .Y (n_5964));
INVX1 g68242(.A (g1384), .Y (n_2));
INVX1 g68299(.A (g6444), .Y (n_1));
INVX1 g67173(.A (g3125), .Y (n_0));
INVX1 g68443(.A (g5148), .Y (n_1813));
INVX1 g68032(.A (g6336), .Y (n_609));
INVX1 g68062(.A (g1825), .Y (n_827));
CLKBUFX1 g68446(.A (g_6165), .Y (g12422));
INVX1 g69642(.A (n_10306), .Y (n_6454));
INVX1 g69644(.A (n_6715), .Y (n_6457));
INVX1 g69646(.A (n_6464), .Y (n_6460));
INVX1 g69652(.A (n_6621), .Y (n_6468));
NOR2X1 g53(.A (n_6503), .B (n_10307), .Y (n_6479));
NAND3X1 g49(.A (n_6464), .B (n_6488), .C (n_6501), .Y (n_3661));
NOR2X1 g54(.A (n_10637), .B (n_7275), .Y (n_6464));
NOR2X1 g69656(.A (g_8896), .B (n_6552), .Y (n_6488));
NAND2X1 g69658(.A (n_10814), .B (n_10529), .Y (n_6490));
INVX1 g69664(.A (n_6490), .Y (n_6501));
OAI21X1 g41(.A0 (n_10313), .A1 (n_6504), .B0 (n_6507), .Y (n_6508));
NAND2X1 g69666(.A (n_9698), .B (n_6503), .Y (n_6504));
INVX1 g47(.A (g_9338), .Y (n_6503));
AOI21X1 g42(.A0 (n_7229), .A1 (n_10313), .B0 (n_6506), .Y (n_6507));
AND2X1 g69667(.A (n_7402), .B (g_9338), .Y (n_7229));
NOR2X1 g69668(.A (n_519), .B (n_9698), .Y (n_6506));
NAND2X1 g69670(.A (n_8793), .B (g_13871), .Y (n_6517));
OR2X1 g31(.A (n_6522), .B (n_6523), .Y (n_6524));
OR2X1 g34(.A (n_10311), .B (n_8792), .Y (n_6522));
NAND2X1 g32(.A (n_6610), .B (n_10863), .Y (n_6523));
INVX1 g12(.A (g_22021), .Y (n_6527));
OAI21X1 g69673(.A0 (g_21806), .A1 (g_22379), .B0 (n_11095), .Y(n_10142));
NAND2X1 g69676(.A (n_11094), .B (g_21806), .Y (n_6539));
AND2X1 g69677(.A (n_6548), .B (g_12922), .Y (n_11105));
INVX1 g26(.A (n_6547), .Y (n_6548));
NAND3X1 g21(.A (n_11120), .B (n_10494), .C (n_6690), .Y (n_6547));
NOR2X1 g24(.A (n_2566), .B (n_6545), .Y (n_10494));
NAND2X1 g25(.A (n_11064), .B (g_19659), .Y (n_6545));
CLKBUFX1 g69681(.A (n_6548), .Y (n_6549));
NOR2X1 g22(.A (n_2566), .B (n_7145), .Y (n_6551));
NOR2X1 g69685(.A (g_8896), .B (n_6552), .Y (n_6553));
NAND2X2 g69686(.A (n_417), .B (n_223), .Y (n_6552));
INVX1 g69693(.A (n_6800), .Y (n_6562));
NOR2X1 g69697(.A (n_447), .B (n_10309), .Y (n_6564));
NAND2X1 g69698(.A (n_7097), .B (g12184), .Y (n_6565));
NAND2X1 g23(.A (n_6565), .B (n_11118), .Y (n_6570));
NAND4X1 g69702(.A (n_6572), .B (n_7260), .C (n_662), .D (g4332), .Y(n_6574));
AND2X1 g69703(.A (g4349), .B (n_1627), .Y (n_6572));
NAND2X1 g69706(.A (n_6572), .B (n_7260), .Y (n_6578));
NOR2X1 g69707(.A (n_10402), .B (n_46), .Y (n_6582));
INVX1 g69713(.A (g1478), .Y (n_6584));
INVX1 g69730(.A (n_8546), .Y (n_6610));
NOR2X1 g69733(.A (g_20909), .B (n_5712), .Y (n_6612));
NOR2X1 g69734(.A (g_17086), .B (n_10311), .Y (n_6618));
AND2X1 g69740(.A (n_6618), .B (n_6620), .Y (n_6621));
NOR2X1 g69741(.A (n_5712), .B (n_8819), .Y (n_6620));
INVX1 g69742(.A (g_17086), .Y (n_6308));
AOI21X1 g69743(.A0 (n_6937), .A1 (n_6938), .B0 (n_9836), .Y (n_6631));
OR2X1 g69744(.A (n_4339), .B (n_4168), .Y (n_6938));
NAND2X1 g29(.A (n_10852), .B (g2421), .Y (n_6937));
AOI21X1 g69750(.A0 (n_6940), .A1 (n_6941), .B0 (n_9775), .Y (n_6639));
OR2X1 g69751(.A (g2361), .B (n_4169), .Y (n_6941));
NAND2X1 g69752(.A (n_10670), .B (g2287), .Y (n_6940));
NOR2X1 g18(.A (n_10264), .B (n_6801), .Y (n_6655));
INVX1 g69772(.A (n_6663), .Y (n_6664));
NAND2X1 g69773(.A (n_10981), .B (n_9453), .Y (n_6663));
INVX2 g69782(.A (n_10976), .Y (n_6666));
AOI21X1 g69786(.A0 (n_6668), .A1 (n_11097), .B0 (n_6669), .Y(n_6670));
NOR2X1 g69787(.A (g2704), .B (g2697), .Y (n_6668));
NOR2X1 g69788(.A (g1291), .B (n_6584), .Y (n_6669));
INVX1 g69790(.A (n_6669), .Y (n_6673));
INVX1 g69791(.A (n_6683), .Y (n_6684));
NAND2X1 g69792(.A (n_6680), .B (n_9717), .Y (n_6683));
OAI21X1 g69793(.A0 (n_3998), .A1 (g1936), .B0 (n_6679), .Y (n_6680));
NAND2X1 g69794(.A (n_6685), .B (g1862), .Y (n_6679));
CLKBUFX3 g69796(.A (n_6676), .Y (n_6677));
CLKBUFX3 g69797(.A (n_6789), .Y (n_6676));
INVX2 g69801(.A (n_6677), .Y (n_6685));
OAI21X1 g69802(.A0 (n_6687), .A1 (n_1183), .B0 (n_6689), .Y (n_6690));
OR4X1 g39(.A (g_22371), .B (g_13838), .C (n_70), .D (n_6923), .Y(n_6687));
NAND3X1 g40(.A (n_10566), .B (n_876), .C (n_6688), .Y (n_6689));
AND2X1 g69803(.A (g_22371), .B (g_13838), .Y (n_6688));
AOI21X1 g69804(.A0 (n_6692), .A1 (n_6693), .B0 (g_13838), .Y(n_6694));
NOR2X1 g69805(.A (n_6923), .B (n_6691), .Y (n_6692));
OR2X1 g69806(.A (g_22371), .B (n_70), .Y (n_6691));
INVX1 g69807(.A (n_1183), .Y (n_6693));
NAND3X1 g69808(.A (n_10566), .B (n_876), .C (g_22371), .Y (n_6695));
NOR2X1 g69812(.A (g2138), .B (g2145), .Y (n_6696));
NAND2X1 g69814(.A (n_10557), .B (g_11413), .Y (n_6697));
INVX1 g69818(.A (n_8846), .Y (n_6705));
CLKBUFX1 g3(.A (n_10678), .Y (n_6707));
NOR2X1 g69826(.A (n_6714), .B (n_6715), .Y (n_6716));
INVX1 g69827(.A (n_7043), .Y (n_6714));
NAND2X1 g69828(.A (n_7042), .B (n_10863), .Y (n_6715));
NAND2X1 g69838(.A (n_10399), .B (n_10401), .Y (n_6577));
NOR2X1 g69843(.A (n_3459), .B (n_6734), .Y (n_6735));
NOR2X1 g69845(.A (g1345), .B (n_10430), .Y (n_6734));
NOR3X1 g69852(.A (g2629), .B (n_6742), .C (n_6666), .Y (n_6746));
INVX1 g69853(.A (g2599), .Y (n_6742));
NOR2X1 g69858(.A (n_9019), .B (n_6756), .Y (n_6757));
AOI21X1 g69860(.A0 (n_6754), .A1 (g1996), .B0 (n_6755), .Y (n_6756));
CLKBUFX1 g69861(.A (n_6752), .Y (n_6754));
INVX1 g69863(.A (n_7099), .Y (n_6752));
NOR2X1 g69867(.A (g2070), .B (n_4516), .Y (n_6755));
INVX1 g69868(.A (n_6752), .Y (n_6758));
CLKBUFX1 g69869(.A (n_7099), .Y (n_6759));
NAND2X1 g69870(.A (n_6762), .B (n_10553), .Y (n_11081));
NAND4X1 g69871(.A (n_2451), .B (n_2452), .C (n_2150), .D (n_6760), .Y(n_10553));
NAND2X1 g69872(.A (g_19911), .B (g_16958), .Y (n_6760));
OR2X1 g69873(.A (n_10123), .B (g_15287), .Y (n_6762));
NOR2X1 g69874(.A (n_6764), .B (n_6766), .Y (n_6767));
INVX1 g69875(.A (n_6762), .Y (n_6764));
NOR2X1 g69876(.A (g_19911), .B (n_6765), .Y (n_6766));
NAND3X1 g69877(.A (n_2451), .B (n_2452), .C (n_2150), .Y (n_6765));
INVX1 g69888(.A (n_10803), .Y (n_6781));
CLKBUFX1 g15(.A (n_10801), .Y (n_6782));
CLKBUFX3 g69889(.A (n_6786), .Y (n_6787));
NOR2X1 g69890(.A (g4054), .B (n_6785), .Y (n_6786));
INVX1 g69891(.A (g3990), .Y (n_6785));
NAND2X1 g69892(.A (n_6789), .B (n_6790), .Y (n_6791));
NAND3X1 g69893(.A (n_898), .B (n_6788), .C (n_10986), .Y (n_6789));
OAI21X1 g69894(.A0 (n_698), .A1 (n_10829), .B0 (g17400), .Y (n_6788));
NOR2X1 g69895(.A (g1862), .B (g1936), .Y (n_6790));
AND2X1 g69897(.A (g3990), .B (g4054), .Y (n_8917));
AND2X1 g69898(.A (n_10495), .B (n_10261), .Y (n_6798));
NOR2X1 g69899(.A (g_18590), .B (n_6796), .Y (n_10495));
NAND3X1 g69900(.A (n_6794), .B (n_10142), .C (n_6057), .Y (n_6796));
AND2X1 g69901(.A (n_11120), .B (n_10628), .Y (n_6794));
NAND2X1 g19(.A (n_10261), .B (n_6799), .Y (n_6800));
INVX1 g69903(.A (n_6796), .Y (n_6799));
NAND2X1 g69904(.A (n_6794), .B (n_10142), .Y (n_6801));
NAND4X1 g69909(.A (n_6806), .B (n_6808), .C (g3945), .D (g16775), .Y(n_6809));
OAI21X1 g69910(.A0 (n_690), .A1 (g_3974), .B0 (n_802), .Y (n_6806));
NOR2X1 g69911(.A (g3990), .B (n_6807), .Y (n_6808));
INVX1 g69912(.A (g4054), .Y (n_6807));
NAND2X1 g63(.A (n_6821), .B (n_6822), .Y (n_6823));
NOR2X1 g66(.A (n_3764), .B (n_7168), .Y (n_6821));
INVX1 g67(.A (n_7354), .Y (n_6822));
OAI21X1 g69938(.A0 (n_6854), .A1 (n_6856), .B0 (n_6857), .Y (n_6858));
AOI21X1 g69939(.A0 (n_6848), .A1 (n_6849), .B0 (n_6853), .Y (n_6854));
INVX1 g69940(.A (n_4969), .Y (n_6848));
NOR2X1 g69941(.A (n_10271), .B (n_5471), .Y (n_6849));
OAI21X1 g69942(.A0 (n_6850), .A1 (n_6851), .B0 (n_6852), .Y (n_6853));
OR2X1 g50(.A (n_4968), .B (n_5471), .Y (n_6850));
CLKBUFX1 g69943(.A (n_4582), .Y (n_6851));
NAND2X1 g69944(.A (n_9693), .B (n_4120), .Y (n_6852));
AND2X1 g69945(.A (n_6852), .B (n_9129), .Y (n_6856));
NAND3X1 g69947(.A (n_5471), .B (n_9553), .C (n_4893), .Y (n_6857));
NOR2X1 g69949(.A (n_9019), .B (n_6865), .Y (n_6866));
AOI21X1 g69951(.A0 (n_10910), .A1 (g1728), .B0 (n_6864), .Y (n_6865));
NOR2X1 g69955(.A (n_4139), .B (n_4006), .Y (n_6864));
OAI21X1 g37(.A0 (n_8882), .A1 (n_8883), .B0 (n_6877), .Y (n_6878));
NAND3X1 g69961(.A (n_6872), .B (n_11207), .C (n_9359), .Y (n_8882));
NAND2X1 g69962(.A (n_6049), .B (n_6095), .Y (n_6872));
AOI22X1 g69965(.A0 (g3813), .A1 (n_9193), .B0 (n_9883), .B1 (n_6876),.Y (n_6877));
AND2X1 g69966(.A (n_6243), .B (n_3596), .Y (n_6876));
NAND2X1 g69970(.A (n_6696), .B (g2130), .Y (n_6880));
INVX2 g69974(.A (n_6891), .Y (n_6892));
INVX2 g7(.A (n_10609), .Y (n_6891));
INVX1 g69978(.A (n_6891), .Y (n_6893));
INVX2 g69980(.A (n_6891), .Y (n_6895));
NOR2X1 g69981(.A (n_10841), .B (n_6896), .Y (n_6897));
INVX1 g69982(.A (n_10607), .Y (n_6896));
NOR2X1 g69984(.A (n_6899), .B (n_6906), .Y (n_6907));
NAND2X1 g69985(.A (n_6553), .B (n_6898), .Y (n_6899));
NAND2X1 g69986(.A (n_584), .B (n_10108), .Y (n_6898));
NAND3X1 g69987(.A (n_6903), .B (n_10805), .C (n_10569), .Y (n_6906));
NOR2X1 g69988(.A (n_10637), .B (n_10639), .Y (n_6903));
NAND2X1 g6(.A (n_6922), .B (g_20208), .Y (n_6923));
INVX1 g70007(.A (g_21813), .Y (n_6922));
AOI21X1 g70008(.A0 (n_6925), .A1 (n_7144), .B0 (n_6926), .Y (n_6927));
AND2X1 g70009(.A (n_9521), .B (g_22605), .Y (n_6925));
NOR2X1 g70010(.A (n_9717), .B (g_22070), .Y (n_6926));
INVX1 g70011(.A (g_22070), .Y (n_6928));
AND2X1 g70021(.A (n_10936), .B (n_11034), .Y (n_6951));
AOI21X1 g70022(.A0 (n_3832), .A1 (g1242), .B0 (n_3831), .Y (n_6953));
AOI21X1 g61508_dup(.A0 (n_3832), .A1 (g1242), .B0 (n_3831), .Y(n_6954));
NOR2X1 g70023(.A (n_6823), .B (n_10974), .Y (n_7235));
NOR2X1 g59_dup(.A (n_10974), .B (n_6823), .Y (n_6956));
INVX1 g70025(.A (n_10708), .Y (n_6958));
CLKBUFX1 g70036(.A (n_6973), .Y (n_6972));
CLKBUFX1 g70039(.A (n_6979), .Y (n_6978));
CLKBUFX1 g70059(.A (n_7004), .Y (n_7003));
OR2X1 g70070(.A (g5046), .B (n_10768), .Y (n_7018));
NAND2X2 g70071(.A (n_7023), .B (n_7024), .Y (n_7025));
INVX1 g70072(.A (n_7022), .Y (n_7023));
NOR2X1 g29_dup(.A (n_10461), .B (n_8759), .Y (n_7022));
NAND3X1 g70075(.A (n_10827), .B (n_8832), .C (n_8796), .Y (n_8756));
NOR2X1 g70076(.A (g1728), .B (n_4139), .Y (n_7024));
INVX1 g71(.A (g_10903), .Y (n_7032));
NAND4X1 g70085(.A (n_7039), .B (n_7116), .C (n_8690), .D (n_10638),.Y (n_7040));
INVX1 g70086(.A (n_8691), .Y (n_7039));
NOR2X1 g70087(.A (n_8546), .B (n_7105), .Y (n_7042));
NOR2X1 g70(.A (n_153), .B (n_10311), .Y (n_7043));
NOR2X1 g70090(.A (n_7045), .B (n_7046), .Y (n_7047));
NAND3X1 g70091(.A (n_10577), .B (n_3740), .C (n_7044), .Y (n_7045));
NAND4X1 g70092(.A (n_10883), .B (n_10576), .C (g3590), .D (g13881),.Y (n_7044));
NAND4X1 g70093(.A (n_4107), .B (n_4683), .C (n_3542), .D (n_4996), .Y(n_7046));
AND2X1 g70094(.A (n_3761), .B (n_3541), .Y (n_7048));
AND2X1 g70095(.A (n_2652), .B (n_4101), .Y (n_7049));
XOR2X1 g70129(.A (n_7085), .B (n_11197), .Y (n_7093));
NOR2X1 g70130(.A (n_10443), .B (n_332), .Y (n_7085));
NOR2X1 g70132(.A (n_7086), .B (n_7087), .Y (n_7088));
NAND4X1 g70133(.A (n_2379), .B (n_2324), .C (n_2343), .D (n_2971), .Y(n_7086));
NAND4X1 g70134(.A (n_2326), .B (n_2659), .C (n_2130), .D (n_2414), .Y(n_7087));
NAND2X1 g70136(.A (n_2353), .B (n_2342), .Y (n_7089));
NAND4X1 g70137(.A (n_2141), .B (n_2030), .C (n_2132), .D (n_3267), .Y(n_7090));
INVX1 g70140(.A (g_15127), .Y (n_7094));
INVX1 g8(.A (g_17653), .Y (n_7097));
NAND2X2 g70141(.A (n_7099), .B (n_7101), .Y (n_7102));
NAND3X1 g70143(.A (n_8880), .B (n_1133), .C (n_2670), .Y (n_7099));
NAND2X1 g70144(.A (n_1709), .B (g_18330), .Y (n_8880));
NOR2X1 g70145(.A (g1996), .B (g2070), .Y (n_7101));
NAND2X1 g70146(.A (n_2670), .B (n_1133), .Y (n_7103));
OR2X1 g70150(.A (n_6517), .B (n_10309), .Y (n_7105));
AND2X1 g70159(.A (n_10569), .B (n_10805), .Y (n_7116));
NOR2X1 g70160(.A (n_10177), .B (n_10176), .Y (n_8909));
NAND3X1 g58(.A (n_7047), .B (n_7048), .C (n_7049), .Y (n_10176));
NAND3X1 g70161(.A (n_7119), .B (n_7120), .C (n_7124), .Y (n_10177));
INVX1 g59(.A (n_7118), .Y (n_7119));
NAND4X1 g70162(.A (n_2140), .B (n_1691), .C (n_5500), .D (n_1850), .Y(n_7118));
AND2X1 g70163(.A (n_2146), .B (n_2138), .Y (n_7120));
AOI21X1 g70164(.A0 (n_11126), .A1 (n_7122), .B0 (n_7123), .Y(n_7124));
INVX1 g70165(.A (n_7121), .Y (n_7122));
NAND3X1 g57(.A (n_10883), .B (g16722), .C (g3606), .Y (n_7121));
NAND2X1 g70166(.A (n_1587), .B (n_5425), .Y (n_7123));
NAND3X1 g70167(.A (n_7130), .B (n_7131), .C (n_7132), .Y (n_7133));
NAND3X1 g70168(.A (n_7127), .B (n_7128), .C (n_9558), .Y (n_7130));
INVX1 g70169(.A (n_6248), .Y (n_7127));
OAI22X1 g70170(.A0 (n_3779), .A1 (n_8909), .B0 (n_3779), .B1(n_6052), .Y (n_7128));
NAND2X1 g70172(.A (n_9300), .B (g3462), .Y (n_7131));
NAND3X1 g70173(.A (n_3779), .B (n_9139), .C (n_3601), .Y (n_7132));
AND2X1 g70179(.A (n_11105), .B (n_7143), .Y (n_7144));
NOR2X1 g70180(.A (n_7140), .B (n_7142), .Y (n_7143));
NAND3X1 g70181(.A (n_11055), .B (n_6928), .C (g_18308), .Y (n_7140));
INVX1 g70182(.A (n_7141), .Y (n_7142));
AND2X1 g70183(.A (n_6690), .B (n_11120), .Y (n_7141));
NAND2X1 g70184(.A (n_7141), .B (n_11055), .Y (n_7145));
AND2X1 g70185(.A (n_11105), .B (g_18308), .Y (n_7146));
NOR2X1 g70187(.A (n_10660), .B (n_191), .Y (n_7150));
NAND4X1 g70199(.A (n_8589), .B (n_7164), .C (n_7165), .D (n_7167), .Y(n_7168));
NAND4X1 g70201(.A (n_10941), .B (n_8588), .C (g16686), .D (g3247), .Y(n_7164));
NAND4X1 g70205(.A (n_11029), .B (n_8588), .C (g3187), .D (g14421), .Y(n_7165));
NAND4X1 g70206(.A (n_8572), .B (n_8588), .C (g3215), .D (g16874), .Y(n_7167));
AND2X1 g75(.A (n_2441), .B (n_2354), .Y (n_7208));
NAND3X1 g70249(.A (n_2966), .B (n_2327), .C (n_2336), .Y (n_7213));
NAND3X1 g72(.A (n_2598), .B (n_1293), .C (n_2149), .Y (n_7214));
NOR2X1 g70250(.A (n_356), .B (n_10341), .Y (n_7217));
NOR2X1 g70251(.A (n_7217), .B (n_7218), .Y (n_7219));
NAND4X1 g67_dup(.A (n_10238), .B (n_10239), .C (n_10240), .D(n_10241), .Y (n_7218));
INVX2 g70266(.A (n_7245), .Y (n_7242));
INVX1 g70267(.A (n_7245), .Y (n_7243));
INVX2 g70269(.A (n_3829), .Y (n_7245));
NOR2X1 g70292(.A (n_7032), .B (n_153), .Y (n_7268));
INVX1 g70296(.A (n_10569), .Y (n_7275));
AOI22X1 g70339(.A0 (n_7330), .A1 (n_7332), .B0 (n_7329), .B1(n_7331), .Y (n_7333));
INVX1 g70340(.A (n_7329), .Y (n_7330));
NAND4X1 g70341(.A (n_7322), .B (n_7325), .C (n_7328), .D (n_3693), .Y(n_7329));
NOR2X1 g70342(.A (n_7320), .B (n_7321), .Y (n_7322));
NAND4X1 g70343(.A (n_2436), .B (n_2334), .C (n_2323), .D (n_2349), .Y(n_7320));
NAND3X1 g70344(.A (n_3265), .B (n_2434), .C (n_2431), .Y (n_7321));
INVX1 g70345(.A (n_7324), .Y (n_7325));
NAND3X1 g70346(.A (n_2601), .B (n_7323), .C (n_3276), .Y (n_7324));
AND2X1 g78(.A (n_1292), .B (n_2148), .Y (n_7323));
NOR2X1 g70347(.A (n_7326), .B (n_7327), .Y (n_7328));
NAND2X1 g70348(.A (n_2388), .B (n_2964), .Y (n_7326));
NAND2X1 g77(.A (n_2338), .B (n_2321), .Y (n_7327));
INVX1 g70349(.A (n_7331), .Y (n_7332));
NOR2X1 g70350(.A (n_247), .B (n_2039), .Y (n_7331));
NAND3X1 g70360(.A (n_7343), .B (n_7344), .C (n_7353), .Y (n_7354));
NAND4X1 g70361(.A (n_1499), .B (n_10941), .C (g3235), .D (g16718), .Y(n_7343));
NAND4X1 g70362(.A (n_1499), .B (n_8586), .C (g3219), .D (g13895), .Y(n_7344));
AND2X1 g70363(.A (n_7348), .B (n_7352), .Y (n_7353));
NAND4X1 g70364(.A (n_11030), .B (n_8588), .C (g3195), .D (g3329), .Y(n_7348));
NAND4X1 g70368(.A (n_8572), .B (n_8588), .C (g_4050), .D (g3191), .Y(n_7352));
INVX4 g70397(.A (n_8588), .Y (n_7383));
CLKBUFX3 g70409(.A (n_7402), .Y (n_7395));
CLKBUFX1 g71109(.A (n_8509), .Y (n_8508));
NAND2X1 g71126(.A (n_10379), .B (n_8534), .Y (n_10101));
OAI21X1 g71130(.A0 (n_1180), .A1 (n_2108), .B0 (g17320), .Y (n_8532));
NOR2X1 g71131(.A (g2153), .B (g2227), .Y (n_8534));
NAND2X2 g71132(.A (n_8864), .B (n_8537), .Y (n_10829));
NOR2X1 g71134(.A (n_10129), .B (n_8800), .Y (n_8537));
NAND3X1 g71137(.A (n_10308), .B (n_7268), .C (n_10806), .Y (n_8540));
NAND2X1 g71139(.A (n_10308), .B (g_16296), .Y (n_8546));
NAND4X1 g71140(.A (n_8548), .B (n_8572), .C (g3243), .D (g16718), .Y(n_8552));
NAND2X2 g71141(.A (n_800), .B (n_8547), .Y (n_8548));
OR2X1 g71142(.A (g_4050), .B (n_8587), .Y (n_8547));
INVX2 g71148(.A (n_8556), .Y (n_8557));
INVX1 g71149(.A (n_8555), .Y (n_8556));
NOR2X1 g71150(.A (g2724), .B (n_10656), .Y (n_8555));
INVX2 g71164(.A (n_8571), .Y (n_8572));
NAND2X1 g71165(.A (n_10839), .B (n_7004), .Y (n_8571));
INVX1 g71172(.A (n_8582), .Y (n_8583));
NAND4X1 g71173(.A (n_10262), .B (n_10263), .C (n_11119), .D(n_10142), .Y (n_8582));
NAND4X1 g71175(.A (n_8586), .B (n_8588), .C (g3231), .D (g13865), .Y(n_8589));
INVX2 g71176(.A (n_8585), .Y (n_8586));
NAND2X1 g71177(.A (n_8584), .B (n_10834), .Y (n_8585));
INVX1 g71178(.A (n_7004), .Y (n_8584));
INVX2 g71179(.A (n_8587), .Y (n_8588));
INVX2 g71180(.A (g3338), .Y (n_8587));
NOR2X1 g71181(.A (n_8770), .B (g1183), .Y (n_8591));
INVX2 g71186(.A (g_13091), .Y (n_8594));
NAND2X1 g71190(.A (n_8601), .B (n_8604), .Y (n_8605));
NAND3X1 g71191(.A (n_8599), .B (n_8600), .C (n_9453), .Y (n_8601));
OAI22X1 g71192(.A0 (n_3775), .A1 (n_7235), .B0 (n_3775), .B1(n_6051), .Y (n_8599));
INVX1 g71193(.A (n_6250), .Y (n_8600));
AOI22X1 g71194(.A0 (g3111), .A1 (n_9772), .B0 (n_3775), .B1 (n_8603),.Y (n_8604));
AND2X1 g43(.A (n_10385), .B (n_3609), .Y (n_8603));
NAND2X2 g71198(.A (n_8615), .B (n_8619), .Y (n_8620));
NAND2X1 g71199(.A (n_8611), .B (n_9717), .Y (n_8615));
INVX1 g71200(.A (n_8610), .Y (n_8611));
AOI21X1 g71201(.A0 (n_8768), .A1 (n_3855), .B0 (n_8609), .Y (n_8610));
AND2X1 g71203(.A (g7916), .B (n_8591), .Y (n_8609));
NAND2X2 g71207(.A (n_8616), .B (n_8618), .Y (n_8619));
OR2X1 g71208(.A (n_9466), .B (n_8768), .Y (n_8616));
NAND3X1 g71209(.A (n_3854), .B (n_3841), .C (n_10005), .Y (n_8618));
NAND2X2 g71214(.A (n_10937), .B (n_8627), .Y (n_8628));
NOR2X1 g71217(.A (g2287), .B (g2361), .Y (n_8627));
AND2X1 g71218(.A (n_10936), .B (n_11034), .Y (n_8629));
NAND2X2 g71219(.A (n_10961), .B (n_8632), .Y (n_8633));
NOR2X1 g71222(.A (g2421), .B (n_4339), .Y (n_8632));
AND2X1 g71223(.A (n_10960), .B (n_11035), .Y (n_8634));
INVX2 g71224(.A (n_8638), .Y (n_8639));
NAND2X1 g71225(.A (n_11210), .B (n_8637), .Y (n_8638));
INVX2 g71228(.A (g4793), .Y (n_8637));
NAND2X1 g71255(.A (n_6880), .B (n_10316), .Y (n_10173));
NOR2X1 g71257(.A (n_10228), .B (n_10175), .Y (n_8810));
INVX2 g71261(.A (n_8675), .Y (n_8676));
NAND3X1 g71262(.A (n_10192), .B (g4966), .C (n_598), .Y (n_8675));
AND2X1 g71265(.A (n_10192), .B (g4966), .Y (n_8677));
NOR2X1 g71267(.A (n_8678), .B (n_7105), .Y (n_8679));
NAND3X1 g71268(.A (n_10638), .B (n_10569), .C (g_16296), .Y (n_8678));
INVX1 g71269(.A (n_8681), .Y (n_8682));
NAND2X1 g71270(.A (n_8680), .B (n_6564), .Y (n_8681));
AND2X1 g56_dup(.A (n_6565), .B (n_6898), .Y (n_8680));
NOR2X1 g71271(.A (n_8686), .B (n_8540), .Y (n_8687));
NAND2X1 g71272(.A (n_6553), .B (n_10308), .Y (n_8686));
AND2X1 g71277(.A (n_6565), .B (n_6898), .Y (n_8690));
NAND2X1 g71278(.A (n_6564), .B (n_6553), .Y (n_8691));
CLKBUFX1 g71279(.A (n_8693), .Y (n_8694));
NOR2X1 g71280(.A (g4785), .B (n_10225), .Y (n_8693));
OAI21X1 g71284(.A0 (n_8702), .A1 (n_8703), .B0 (n_8705), .Y (n_8706));
NAND3X1 g71285(.A (n_8697), .B (g28753), .C (n_9521), .Y (n_8702));
OR2X1 g71286(.A (n_10684), .B (n_2078), .Y (n_8697));
AND2X1 g71289(.A (n_2078), .B (n_10684), .Y (n_8703));
AOI22X1 g71290(.A0 (g5120), .A1 (n_9454), .B0 (n_8704), .B1 (n_3244),.Y (n_8705));
AND2X1 g71291(.A (n_9698), .B (n_3618), .Y (n_8704));
INVX1 g45(.A (g28753), .Y (n_8707));
NAND2X1 g71314(.A (n_8731), .B (n_8735), .Y (n_8736));
INVX1 g71315(.A (n_8730), .Y (n_8731));
NAND4X1 g71316(.A (n_11194), .B (n_1575), .C (n_11195), .D (n_1855),.Y (n_8730));
INVX1 g71317(.A (n_8734), .Y (n_8735));
NAND4X1 g71318(.A (n_3286), .B (n_10368), .C (n_8733), .D (n_1859),.Y (n_8734));
NAND4X1 g71320(.A (n_2339), .B (n_1695), .C (g5264), .D (g17639), .Y(n_8733));
NOR2X1 g71335(.A (n_262), .B (n_8885), .Y (n_8757));
NOR2X1 g62211_dup(.A (n_262), .B (n_8886), .Y (n_8758));
AND2X1 g71336(.A (g17316), .B (n_8756), .Y (n_8759));
AOI21X1 g71337(.A0 (n_6951), .A1 (g1585), .B0 (n_3873), .Y (n_8761));
AOI21X1 g61378_dup(.A0 (n_6951), .A1 (g1585), .B0 (n_3873), .Y(n_8762));
AOI21X1 g71338(.A0 (n_11211), .A1 (n_10764), .B0 (n_3870), .Y(n_8763));
AOI21X1 g61379_dup(.A0 (n_11212), .A1 (n_10764), .B0 (n_3870), .Y(n_8764));
CLKBUFX1 g71342(.A (n_8769), .Y (n_8768));
INVX2 g71343(.A (n_8770), .Y (n_8769));
INVX2 g71344(.A (g1171), .Y (n_8770));
INVX1 g71349(.A (n_8777), .Y (n_8776));
CLKBUFX3 g71350(.A (n_8778), .Y (n_8777));
INVX1 g71363(.A (n_8793), .Y (n_8792));
CLKBUFX1 g71368(.A (n_8800), .Y (n_8799));
CLKBUFX1 g71372(.A (n_8807), .Y (n_8806));
CLKBUFX1 g71374(.A (n_8810), .Y (n_8809));
NAND4X1 g71375(.A (n_8679), .B (n_8682), .C (n_8687), .D (n_8818), .Y(n_8819));
NOR2X1 g71376(.A (n_8816), .B (n_8817), .Y (n_8818));
NAND2X1 g71377(.A (n_10310), .B (g_21799), .Y (n_8816));
OR2X1 g71382(.A (n_86), .B (n_10309), .Y (n_8817));
OR2X1 g71384(.A (n_8817), .B (n_8820), .Y (n_8821));
NAND3X1 g71385(.A (n_8679), .B (n_8682), .C (n_8687), .Y (n_8820));
NOR2X1 g71394(.A (g7916), .B (n_8835), .Y (n_8836));
NAND2X2 g71395(.A (n_8831), .B (n_8834), .Y (n_8835));
NAND2X2 g71396(.A (n_1833), .B (n_1255), .Y (n_8831));
AOI21X1 g71397(.A0 (n_8833), .A1 (n_10647), .B0 (n_1636), .Y(n_8834));
INVX1 g71398(.A (n_8832), .Y (n_8833));
AND2X1 g71399(.A (g1183), .B (n_8770), .Y (n_8832));
INVX1 g71400(.A (g7916), .Y (n_8837));
NOR2X1 g71402(.A (n_1636), .B (n_8839), .Y (n_8840));
INVX1 g71403(.A (n_8831), .Y (n_8839));
AND2X1 g71409(.A (n_10724), .B (n_10647), .Y (n_8846));
NAND2X1 g71414(.A (n_8848), .B (n_10286), .Y (n_8850));
NAND2X1 g71415(.A (n_10956), .B (g1300), .Y (n_8848));
INVX1 g71419(.A (n_8848), .Y (n_8855));
NOR2X1 g71426(.A (n_10120), .B (g1221), .Y (n_8864));
OR2X1 g71439(.A (n_512), .B (n_10395), .Y (n_8885));
OR2X1 g63195_dup(.A (n_512), .B (n_10395), .Y (n_8886));
INVX1 g71440(.A (n_10225), .Y (n_10175));
CLKBUFX3 g71446(.A (n_8898), .Y (n_8895));
CLKBUFX1 g71452(.A (n_10227), .Y (n_8906));
CLKBUFX1 g71453(.A (n_8909), .Y (n_8908));
CLKBUFX1 g71458(.A (n_8915), .Y (n_8913));
CLKBUFX1 g71463(.A (g35), .Y (n_8921));
INVX8 g71489(.A (n_9107), .Y (n_8955));
INVX8 g71515(.A (n_9107), .Y (n_9000));
INVX2 g71522(.A (n_10385), .Y (n_9019));
INVX8 g71571(.A (n_9129), .Y (n_9091));
INVX4 g71584(.A (n_10687), .Y (n_9107));
INVX8 g71600(.A (n_10687), .Y (n_9129));
INVX1 g71609(.A (n_9139), .Y (n_9141));
INVX2 g71610(.A (n_9107), .Y (n_9139));
INVX1 g71618(.A (n_9129), .Y (n_9156));
INVX4 g71628(.A (n_9176), .Y (n_9172));
INVX1 g71630(.A (n_9167), .Y (n_9176));
INVX4 g71640(.A (n_9209), .Y (n_9193));
BUFX3 g71654(.A (n_10687), .Y (n_9209));
INVX4 g71655(.A (n_9269), .Y (n_9218));
INVX4 g71664(.A (n_9269), .Y (n_9234));
INVX4 g71668(.A (n_9269), .Y (n_9240));
INVX4 g71677(.A (n_9269), .Y (n_9256));
INVX4 g71686(.A (n_9279), .Y (n_9269));
INVX4 g71699(.A (n_9129), .Y (n_9279));
INVX1 g71705(.A (g35), .Y (n_9297));
INVX8 g71713(.A (n_9300), .Y (n_9311));
INVX2 g71723(.A (n_9300), .Y (n_9333));
INVX8 g71730(.A (n_9358), .Y (n_9300));
INVX2 g71739(.A (n_9351), .Y (n_9353));
CLKBUFX1 g71740(.A (n_9358), .Y (n_9351));
INVX8 g71747(.A (n_9371), .Y (n_9359));
INVX4 g71767(.A (n_9358), .Y (n_9371));
INVX1 g71770(.A (n_9398), .Y (n_9404));
BUFX3 g71773(.A (n_9358), .Y (n_9398));
BUFX3 g71775(.A (n_10949), .Y (n_9358));
INVX2 g71780(.A (n_9425), .Y (n_9419));
INVX4 g71782(.A (n_9419), .Y (n_9422));
INVX8 g71784(.A (n_9491), .Y (n_9425));
INVX2 g71788(.A (n_9425), .Y (n_9431));
INVX1 g71796(.A (n_9448), .Y (n_9443));
CLKBUFX1 g71799(.A (n_9493), .Y (n_9448));
INVX1 g71802(.A (n_9453), .Y (n_9454));
CLKBUFX3 g71804(.A (n_9493), .Y (n_9453));
INVX1 g71807(.A (n_9466), .Y (n_9461));
BUFX3 g71810(.A (n_9493), .Y (n_9466));
INVX1 g71812(.A (n_10952), .Y (n_9469));
INVX2 g71824(.A (n_9493), .Y (n_9491));
INVX4 g71828(.A (n_10716), .Y (n_9493));
INVX2 g71836(.A (n_9501), .Y (n_9505));
INVX2 g71837(.A (n_10716), .Y (n_9501));
INVX1 g71854(.A (n_9521), .Y (n_9526));
INVX4 g71863(.A (n_10376), .Y (n_9521));
INVX8 g71895(.A (n_9599), .Y (n_9558));
INVX8 g71898(.A (n_9553), .Y (n_9599));
INVX4 g71899(.A (n_10376), .Y (n_9553));
INVX1 g71917(.A (n_9628), .Y (n_9630));
INVX8 g71918(.A (n_9627), .Y (n_9628));
INVX4 g71931(.A (n_10782), .Y (n_9627));
INVX2 g71941(.A (n_10782), .Y (n_9651));
INVX4 g71953(.A (n_9672), .Y (n_9681));
INVX4 g71956(.A (n_9664), .Y (n_9672));
INVX2 g71961(.A (n_9664), .Y (n_9693));
BUFX3 g71962(.A (n_10950), .Y (n_9664));
INVX1 g71964(.A (n_9698), .Y (n_9697));
CLKBUFX1 g71972(.A (n_10949), .Y (n_9698));
INVX8 g72006(.A (n_9772), .Y (n_9750));
INVX4 g72018(.A (n_9717), .Y (n_9772));
CLKBUFX3 g72019(.A (n_10949), .Y (n_9717));
INVX8 g72031(.A (n_9775), .Y (n_9797));
INVX4 g72034(.A (n_9834), .Y (n_9775));
INVX8 g72036(.A (n_9775), .Y (n_9811));
INVX2 g72047(.A (n_9836), .Y (n_9830));
INVX4 g72052(.A (n_9834), .Y (n_9836));
BUFX3 g72060(.A (n_10949), .Y (n_9834));
INVX2 g72068(.A (n_9874), .Y (n_9856));
BUFX3 g72069(.A (n_9874), .Y (n_9862));
INVX1 g72071(.A (n_9862), .Y (n_9871));
INVX2 g72074(.A (n_10376), .Y (n_9874));
INVX1 g72080(.A (n_9884), .Y (n_9883));
CLKBUFX3 g72086(.A (n_10376), .Y (n_9884));
INVX8 g72088(.A (n_9928), .Y (n_9894));
INVX8 g72097(.A (n_9894), .Y (n_9903));
INVX4 g72120(.A (n_9903), .Y (n_9940));
CLKBUFX3 g72129(.A (n_10376), .Y (n_9928));
CLKBUFX1 g72132(.A (n_10376), .Y (n_9952));
INVX2 g72146(.A (n_9664), .Y (n_9976));
INVX1 g72148(.A (n_9952), .Y (n_9978));
INVX8 g72159(.A (n_10078), .Y (n_9992));
INVX8 g72169(.A (n_10078), .Y (n_10005));
INVX4 g72203(.A (n_10078), .Y (n_10063));
INVX8 g72221(.A (n_10013), .Y (n_10078));
BUFX3 g72222(.A (n_10949), .Y (n_10013));
INVX2 g72224(.A (n_10100), .Y (n_10097));
INVX2 g72225(.A (n_10100), .Y (n_10099));
INVX2 g72226(.A (n_10101), .Y (n_10100));
INVX1 g72228(.A (n_10107), .Y (n_10103));
INVX1 g72232(.A (n_10108), .Y (n_10107));
INVX2 g72233(.A (n_10631), .Y (n_10108));
CLKBUFX1 g72237(.A (n_10113), .Y (n_10112));
CLKBUFX1 g72239(.A (n_10532), .Y (n_10115));
CLKBUFX1 g72242(.A (n_10120), .Y (n_10119));
CLKBUFX1 g72245(.A (n_10125), .Y (n_10123));
CLKBUFX1 g72249(.A (n_10129), .Y (n_10128));
INVX1 g72253(.A (n_10139), .Y (n_10134));
INVX1 g72259(.A (g5016), .Y (n_10139));
CLKBUFX1 g72292(.A (n_10185), .Y (n_10184));
INVX1 g72294(.A (n_10192), .Y (n_10188));
INVX1 g72299(.A (g4991), .Y (n_10192));
CLKBUFX1 g72301(.A (n_10197), .Y (n_10196));
INVX1 g72303(.A (n_10200), .Y (n_10199));
CLKBUFX2 g72304(.A (n_10202), .Y (n_10200));
INVX1 g72305(.A (n_10202), .Y (n_10201));
CLKBUFX1 g72306(.A (n_10804), .Y (n_10202));
INVX2 g72307(.A (n_10804), .Y (n_10203));
CLKBUFX1 g72308(.A (n_10206), .Y (n_10205));
AND2X1 g72314(.A (n_10213), .B (n_11129), .Y (n_10214));
INVX2 g72315(.A (n_10997), .Y (n_10213));
INVX1 g72321(.A (n_10771), .Y (n_10216));
INVX1 g72322(.A (g5046), .Y (n_10217));
NOR2X1 g72326(.A (n_10224), .B (n_10226), .Y (n_10227));
CLKBUFX1 g72327(.A (g4785), .Y (n_10224));
INVX1 g72328(.A (n_10225), .Y (n_10226));
INVX2 g72329(.A (g4709), .Y (n_10225));
INVX1 g72330(.A (g4785), .Y (n_10228));
AND2X1 g51(.A (n_2444), .B (n_2331), .Y (n_10229));
NOR2X1 g72337(.A (n_10516), .B (n_10512), .Y (n_10238));
INVX1 g72338(.A (n_10514), .Y (n_10239));
NOR2X1 g72339(.A (n_7213), .B (n_7214), .Y (n_10240));
NOR2X1 g72340(.A (n_2442), .B (n_3326), .Y (n_10241));
OR2X1 g72343(.A (n_3364), .B (n_11077), .Y (n_10242));
NAND3X1 g72344(.A (n_11076), .B (n_1275), .C (n_3365), .Y (n_10243));
AOI21X1 g72345(.A0 (g1345), .A1 (g1361), .B0 (n_2177), .Y (n_10247));
CLKBUFX1 g72347(.A (n_10802), .Y (n_10245));
NOR2X1 g72356(.A (n_10257), .B (n_10260), .Y (n_10261));
NAND2X1 g72357(.A (n_11120), .B (n_10142), .Y (n_10257));
NAND4X1 g72358(.A (n_10628), .B (n_11094), .C (n_10259), .D(g_16311), .Y (n_10260));
AND2X1 g72360(.A (g_11293), .B (g_15691), .Y (n_10259));
AND2X1 g72361(.A (n_10628), .B (g_11293), .Y (n_10262));
AND2X1 g72362(.A (n_11094), .B (g_15691), .Y (n_10263));
INVX1 g72363(.A (n_10263), .Y (n_10264));
NAND2X1 g72367(.A (n_10270), .B (n_10271), .Y (n_10901));
NAND2X1 g72368(.A (n_10268), .B (n_10322), .Y (n_10270));
OAI21X1 g72369(.A0 (n_1298), .A1 (n_10829), .B0 (g17291), .Y(n_10268));
NOR2X1 g72371(.A (n_4120), .B (g1592), .Y (n_10271));
NAND2X1 g72379(.A (n_10283), .B (n_11122), .Y (n_10285));
AOI21X1 g72380(.A0 (n_10281), .A1 (n_10282), .B0 (n_8855), .Y(n_10283));
NOR2X1 g72381(.A (n_10867), .B (n_10280), .Y (n_10281));
INVX1 g72382(.A (g2697), .Y (n_10280));
AND2X1 g72384(.A (g2704), .B (n_11099), .Y (n_10282));
AND2X1 g72386(.A (n_10289), .B (g1585), .Y (n_10290));
AND2X1 g72387(.A (n_10288), .B (n_11122), .Y (n_10289));
NOR2X1 g72388(.A (n_10287), .B (n_8855), .Y (n_10288));
INVX1 g72389(.A (n_10286), .Y (n_10287));
NAND2X1 g72390(.A (n_10282), .B (g2697), .Y (n_10286));
CLKBUFX1 g72391(.A (n_10998), .Y (n_10296));
NAND2X1 g72402(.A (n_10306), .B (n_10312), .Y (n_10313));
NOR2X1 g72403(.A (n_10304), .B (n_8819), .Y (n_10306));
NAND3X1 g72404(.A (n_6612), .B (n_6618), .C (n_10303), .Y (n_10304));
NOR2X1 g72405(.A (n_10311), .B (g_5342), .Y (n_10303));
NOR2X1 g72407(.A (n_10307), .B (n_10311), .Y (n_10312));
INVX2 g72408(.A (g_10233), .Y (n_10307));
INVX2 g72409(.A (n_10310), .Y (n_10311));
INVX2 g72410(.A (n_10309), .Y (n_10310));
INVX2 g44(.A (n_10308), .Y (n_10309));
NAND2X2 g72411(.A (n_7094), .B (g_17653), .Y (n_10308));
INVX1 g72412(.A (n_10307), .Y (n_10314));
NAND3X1 g72413(.A (n_11138), .B (n_6612), .C (n_6618), .Y (n_10315));
AOI21X1 g72414(.A0 (n_10319), .A1 (n_10871), .B0 (n_10320), .Y(n_10321));
NOR2X1 g72415(.A (n_10317), .B (n_10318), .Y (n_10319));
INVX1 g72416(.A (n_10316), .Y (n_10317));
AND2X1 g72417(.A (n_11065), .B (n_10708), .Y (n_10316));
NAND3X1 g72418(.A (n_6697), .B (n_10723), .C (n_10649), .Y (n_10318));
NOR2X1 g72419(.A (n_10318), .B (n_10173), .Y (n_10320));
CLKBUFX1 g72420(.A (n_10322), .Y (n_10323));
NOR2X1 g72421(.A (n_10318), .B (n_10173), .Y (n_10322));
AOI21X1 g72422(.A0 (n_10327), .A1 (n_10328), .B0 (n_10329), .Y(n_10330));
NAND4X1 g72423(.A (n_11076), .B (n_10325), .C (n_10426), .D (g7946),.Y (n_10327));
INVX1 g72425(.A (n_1276), .Y (n_10325));
OR2X1 g72427(.A (n_3849), .B (n_6781), .Y (n_10328));
OR2X1 g72428(.A (g1532), .B (n_461), .Y (n_10329));
AOI21X1 g72436(.A0 (n_10342), .A1 (g5485), .B0 (n_10345), .Y(n_10346));
NAND2X1 g72437(.A (n_10781), .B (n_10341), .Y (n_10342));
AND2X1 g72439(.A (n_1484), .B (n_2443), .Y (n_10341));
NOR2X1 g72440(.A (n_10344), .B (n_10342), .Y (n_10345));
OAI21X1 g72441(.A0 (g5481), .A1 (g5475), .B0 (n_10343), .Y (n_10344));
NAND2X1 g72442(.A (g5481), .B (g5475), .Y (n_10343));
INVX1 g72443(.A (n_10342), .Y (n_10347));
NOR2X1 g72452(.A (n_10357), .B (n_10362), .Y (n_10363));
NOR2X1 g72453(.A (n_10687), .B (g5619), .Y (n_10357));
AOI21X1 g72455(.A0 (n_10948), .A1 (n_10519), .B0 (n_10361), .Y(n_10362));
OAI21X1 g72459(.A0 (n_10948), .A1 (g4821), .B0 (n_10687), .Y(n_10361));
NAND4X1 g72461(.A (g5248), .B (n_1695), .C (n_10833), .D (g14597), .Y(n_10368));
CLKBUFX3 g72463(.A (g5343), .Y (g25219));
INVX1 g72465(.A (g5343), .Y (n_10369));
AOI21X1 g72467(.A0 (n_10371), .A1 (n_10374), .B0 (n_10376), .Y(n_10377));
OR2X1 g72468(.A (g2227), .B (n_4699), .Y (n_10371));
NAND2X1 g72469(.A (g2153), .B (n_10373), .Y (n_10374));
INVX1 g72470(.A (n_10372), .Y (n_10373));
NAND2X1 g35_dup(.A (n_8532), .B (n_10763), .Y (n_10372));
INVX4 g72471(.A (n_10949), .Y (n_10376));
CLKBUFX1 g72473(.A (n_10372), .Y (n_10378));
INVX2 g72474(.A (n_10379), .Y (n_10380));
NAND2X2 g72475(.A (n_10763), .B (n_8532), .Y (n_10379));
NAND2X1 g72476(.A (n_10386), .B (n_10387), .Y (n_10388));
OAI21X1 g72477(.A0 (n_4840), .A1 (n_10383), .B0 (n_10385), .Y(n_10386));
NOR2X1 g72478(.A (n_10381), .B (n_10382), .Y (n_10383));
INVX1 g72479(.A (n_4839), .Y (n_10381));
INVX1 g72480(.A (n_1592), .Y (n_10382));
BUFX3 g72481(.A (n_10687), .Y (n_10385));
NAND2X1 g20(.A (n_10078), .B (g20049), .Y (n_10387));
NAND4X1 g72484(.A (n_10390), .B (n_10391), .C (n_10392), .D(n_10394), .Y (n_10395));
INVX1 g72485(.A (n_6574), .Y (n_10390));
NOR2X1 g72486(.A (n_23), .B (n_6578), .Y (n_10391));
NOR2X1 g72487(.A (n_7247), .B (n_46), .Y (n_10392));
NOR2X1 g72488(.A (n_3624), .B (n_46), .Y (n_10394));
NOR2X1 g72490(.A (n_10396), .B (n_10397), .Y (n_10398));
NAND2X1 g72491(.A (n_10391), .B (n_10392), .Y (n_10396));
OR2X1 g72492(.A (n_46), .B (n_6574), .Y (n_10397));
INVX1 g72493(.A (n_10397), .Y (n_10399));
INVX1 g72494(.A (n_10396), .Y (n_10400));
NOR2X1 g72495(.A (n_7247), .B (n_23), .Y (n_10401));
INVX1 g72496(.A (n_10401), .Y (n_10402));
NOR2X1 g72497(.A (n_10504), .B (g_18739), .Y (n_10404));
OR2X1 g72502(.A (n_10412), .B (n_10415), .Y (n_10416));
NAND4X1 g72503(.A (n_11218), .B (n_11219), .C (n_2968), .D (n_10411),.Y (n_10412));
NAND4X1 g72504(.A (n_6787), .B (n_690), .C (g4031), .D (g3913), .Y(n_11218));
NAND3X1 g73(.A (g3909), .B (n_803), .C (n_8917), .Y (n_10411));
NAND4X1 g72506(.A (n_6809), .B (n_10413), .C (n_10414), .D (n_1851),.Y (n_10415));
NAND4X1 g72507(.A (n_3894), .B (n_6808), .C (g3957), .D (g16748), .Y(n_10413));
NAND4X1 g72508(.A (n_3894), .B (n_4988), .C (g3941), .D (g13906), .Y(n_10414));
AND2X1 g72510(.A (n_11037), .B (n_8807), .Y (g25114));
AND2X1 g72514(.A (n_10425), .B (n_10426), .Y (n_10427));
NAND3X1 g72515(.A (n_10242), .B (n_10424), .C (n_10243), .Y(n_10425));
INVX1 g72516(.A (n_10423), .Y (n_10424));
AOI21X1 g72517(.A0 (n_10245), .A1 (n_10422), .B0 (n_10247), .Y(n_10423));
INVX1 g72518(.A (g1367), .Y (n_10422));
OR2X1 g72519(.A (g1322), .B (g1333), .Y (n_10426));
NAND2X1 g72520(.A (n_10428), .B (n_10426), .Y (n_10429));
NAND3X1 g72521(.A (n_10242), .B (n_10243), .C (n_10247), .Y(n_10428));
INVX1 g72522(.A (n_10430), .Y (n_10431));
NAND3X1 g72523(.A (n_10242), .B (n_10243), .C (n_10245), .Y(n_10430));
AOI21X1 g28(.A0 (n_10445), .A1 (n_10446), .B0 (n_10447), .Y(n_10448));
INVX2 g72533(.A (n_10444), .Y (n_10445));
NAND3X1 g72534(.A (n_2391), .B (n_10443), .C (n_69), .Y (n_10444));
AND2X1 g72535(.A (n_2352), .B (n_1457), .Y (n_10443));
XOR2X1 g72536(.A (g6167), .B (g6173), .Y (n_10446));
AND2X1 g72537(.A (n_10444), .B (g6177), .Y (n_10447));
NAND2X2 g72538(.A (n_2391), .B (n_69), .Y (n_3784));
NAND2X1 g72549(.A (n_10460), .B (n_10466), .Y (n_10467));
NAND2X1 g72550(.A (n_7025), .B (n_4190), .Y (n_10460));
NAND3X1 g72551(.A (n_10913), .B (n_7024), .C (g1816), .Y (n_10466));
NAND2X1 g72553(.A (n_10462), .B (n_10463), .Y (n_10464));
INVX1 g72554(.A (n_10461), .Y (n_10462));
NAND2X2 g72555(.A (n_2983), .B (n_1241), .Y (n_10461));
NAND2X1 g72556(.A (n_8756), .B (g17316), .Y (n_10463));
INVX1 g72559(.A (n_10472), .Y (n_10473));
NAND4X1 g72560(.A (n_10470), .B (n_1458), .C (n_10623), .D (g34028),.Y (n_10472));
NAND4X1 g72561(.A (n_8639), .B (n_8694), .C (n_10905), .D (g4754), .Y(n_10470));
NAND2X2 g72563(.A (n_10470), .B (g34028), .Y (n_3612));
AND2X1 g72564(.A (n_1458), .B (n_10623), .Y (n_10475));
INVX2 g72583(.A (n_10503), .Y (n_10499));
CLKBUFX1 g72586(.A (n_10504), .Y (n_10503));
CLKBUFX1 g72587(.A (n_10505), .Y (n_10504));
INVX2 g72588(.A (g_15838), .Y (n_10505));
CLKBUFX1 g72589(.A (n_10508), .Y (n_10506));
NAND4X1 g72593(.A (n_10513), .B (n_10515), .C (n_10517), .D(n_10518), .Y (n_10519));
NOR2X1 g72594(.A (n_2442), .B (n_10512), .Y (n_10513));
NAND2X1 g72595(.A (n_2438), .B (n_2329), .Y (n_10512));
NOR2X1 g72596(.A (n_3326), .B (n_10514), .Y (n_10515));
NAND2X1 g72597(.A (n_2382), .B (n_3281), .Y (n_10514));
INVX1 g72598(.A (n_10516), .Y (n_10517));
NAND3X1 g72599(.A (n_7208), .B (n_10229), .C (n_3268), .Y (n_10516));
NOR2X1 g72600(.A (n_7213), .B (n_7214), .Y (n_10518));
NAND4X1 g72601(.A (n_10526), .B (n_10527), .C (n_10528), .D (n_3388),.Y (n_10532));
INVX1 g72602(.A (n_10525), .Y (n_10526));
NAND3X1 g72603(.A (n_10520), .B (g_20951), .C (n_10524), .Y(n_10525));
AND2X1 g72604(.A (g_20952), .B (n_11116), .Y (n_10520));
INVX1 g72606(.A (n_10522), .Y (n_10524));
INVX1 g72608(.A (g_5029), .Y (n_10522));
NOR2X1 g72609(.A (g_8896), .B (n_780), .Y (n_10527));
INVX1 g72610(.A (g_18996), .Y (n_10528));
INVX1 g72611(.A (n_10529), .Y (n_3388));
INVX1 g72613(.A (g_19789), .Y (n_10529));
NOR2X1 g72614(.A (n_10534), .B (n_10520), .Y (n_10535));
NOR2X1 g72615(.A (n_11113), .B (g_20952), .Y (n_10534));
NOR2X1 g72628(.A (g_7563), .B (n_11027), .Y (n_11095));
INVX2 g72630(.A (g_22349), .Y (n_10557));
NAND4X1 g72631(.A (n_10558), .B (n_10708), .C (n_11065), .D(n_10649), .Y (n_10560));
NAND2X2 g26_dup(.A (n_10505), .B (n_8594), .Y (n_10558));
NOR2X1 g72634(.A (n_10564), .B (n_10565), .Y (n_10566));
OR2X1 g17(.A (n_11110), .B (n_10563), .Y (n_10564));
INVX1 g72635(.A (g_19515), .Y (n_10563));
OR2X1 g72636(.A (g_22600), .B (g_21318), .Y (n_10565));
NOR2X1 g72637(.A (g_21318), .B (n_11110), .Y (n_10567));
INVX1 g72638(.A (n_10563), .Y (n_10568));
AND2X1 g72639(.A (g_20952), .B (n_11116), .Y (n_10569));
NAND4X1 g72641(.A (n_10573), .B (n_10576), .C (g16627), .D (g3602),.Y (n_10577));
MX2X1 g72644(.A (g_9298), .B (n_11091), .S0 (n_10898), .Y (n_10573));
NOR2X1 g72646(.A (n_6979), .B (g3639), .Y (n_10576));
NAND2X1 g72647(.A (n_10883), .B (g11388), .Y (n_10578));
NAND3X1 g72648(.A (n_10587), .B (n_10588), .C (n_10589), .Y(n_10590));
NAND2X1 g72649(.A (n_10582), .B (n_9091), .Y (n_10587));
OAI21X1 g72650(.A0 (n_4805), .A1 (n_10579), .B0 (n_10581), .Y(n_10582));
OR2X1 g72651(.A (n_11055), .B (n_3177), .Y (n_10579));
OR2X1 g72652(.A (n_1286), .B (n_10580), .Y (n_10581));
OR2X1 g72653(.A (n_284), .B (n_3177), .Y (n_10580));
NAND3X1 g72658(.A (n_9894), .B (n_3177), .C (n_11055), .Y (n_10588));
NAND2X1 g72659(.A (n_9884), .B (g20899), .Y (n_10589));
NAND2X2 g72661(.A (n_9493), .B (n_10600), .Y (n_10601));
OAI21X1 g72665(.A0 (n_10596), .A1 (n_10597), .B0 (n_10599), .Y(n_10600));
NOR2X1 g72666(.A (n_10595), .B (n_4213), .Y (n_10596));
AND2X1 g72667(.A (n_3409), .B (n_685), .Y (n_10595));
NAND3X1 g72668(.A (n_1578), .B (n_477), .C (g4878), .Y (n_10597));
INVX1 g72669(.A (n_10598), .Y (n_10599));
AOI21X1 g72670(.A0 (n_1819), .A1 (n_844), .B0 (n_1830), .Y (n_10598));
NOR2X1 g72671(.A (n_8807), .B (n_11037), .Y (n_10833));
NAND3X1 g72676(.A (n_10607), .B (n_10846), .C (g2735), .Y (n_10609));
NOR2X1 g72677(.A (n_11013), .B (g2748), .Y (n_10607));
NOR2X1 g72682(.A (n_10613), .B (n_10617), .Y (n_10618));
XOR2X1 g72683(.A (n_6027), .B (n_878), .Y (n_10613));
NAND2X2 g72684(.A (n_5799), .B (n_10616), .Y (n_10617));
NAND2X2 g72686(.A (n_5617), .B (n_5705), .Y (n_10614));
AND2X1 g72687(.A (g1657), .B (g1624), .Y (n_10616));
INVX2 g72688(.A (n_10620), .Y (n_10621));
OR2X1 g72689(.A (n_8807), .B (n_11038), .Y (n_10620));
AND2X1 g72691(.A (n_11198), .B (g5990), .Y (n_10622));
CLKBUFX1 g72692(.A (n_10622), .Y (n_10623));
AND2X1 g72693(.A (n_10626), .B (n_11064), .Y (n_10628));
OR2X1 g72694(.A (n_10625), .B (n_11028), .Y (n_10626));
NAND2X1 g72695(.A (n_10624), .B (g_20837), .Y (n_10625));
INVX1 g72696(.A (g_7563), .Y (n_10624));
AOI21X1 g72699(.A0 (n_10633), .A1 (n_10634), .B0 (n_10637), .Y(n_10638));
INVX1 g72700(.A (n_10632), .Y (n_10633));
NAND2X2 g72701(.A (n_10630), .B (n_10631), .Y (n_10632));
INVX2 g72702(.A (g_22034), .Y (n_10630));
INVX2 g72703(.A (g_18238), .Y (n_10631));
INVX2 g72706(.A (g_22038), .Y (n_10634));
NAND2X1 g72707(.A (n_10522), .B (g_20951), .Y (n_10637));
NOR2X1 g72708(.A (n_552), .B (n_10632), .Y (n_10639));
INVX1 g72713(.A (n_10647), .Y (n_10644));
CLKBUFX1 g72717(.A (n_10649), .Y (n_10647));
CLKBUFX1 g72722(.A (n_10656), .Y (n_10650));
CLKBUFX2 g72727(.A (n_10657), .Y (n_10660));
INVX1 g72728(.A (n_10667), .Y (n_10664));
INVX1 g72731(.A (n_10404), .Y (n_10667));
INVX1 g72732(.A (n_10670), .Y (n_10669));
INVX2 g72733(.A (n_10671), .Y (n_10670));
CLKBUFX3 g72734(.A (n_10672), .Y (n_10671));
CLKBUFX3 g72735(.A (n_10937), .Y (n_10672));
INVX1 g72737(.A (n_10675), .Y (n_10674));
CLKBUFX2 g72738(.A (n_10937), .Y (n_10675));
XOR2X1 g72739(.A (g_20614), .B (n_10125), .Y (n_10678));
AOI21X1 g72741(.A0 (n_10686), .A1 (n_9167), .B0 (n_10689), .Y(n_10690));
OAI21X1 g72742(.A0 (g28753), .A1 (g21245), .B0 (n_10685), .Y(n_10686));
AND2X1 g43_dup(.A (n_2416), .B (g34026), .Y (g28753));
OR2X1 g72744(.A (n_3244), .B (n_10684), .Y (n_10685));
NAND2X1 g72746(.A (n_10682), .B (n_10683), .Y (n_10684));
NOR2X1 g72747(.A (n_3990), .B (n_3385), .Y (n_10682));
NOR2X1 g72748(.A (n_8736), .B (n_3044), .Y (n_10683));
BUFX3 g72749(.A (n_10687), .Y (n_9167));
BUFX3 g72750(.A (g35), .Y (n_10687));
NOR2X1 g72751(.A (n_9167), .B (g5272), .Y (n_10689));
AND2X1 g72754(.A (n_2416), .B (g34026), .Y (n_10693));
INVX2 g72755(.A (n_10699), .Y (n_10700));
NAND2X1 g72756(.A (n_10696), .B (n_10698), .Y (n_10699));
NAND3X1 g72757(.A (n_10216), .B (n_10695), .C (n_10217), .Y(n_10696));
AND2X1 g72758(.A (n_10766), .B (n_10694), .Y (n_10695));
INVX1 g72759(.A (g5052), .Y (n_10694));
OR2X1 g72760(.A (n_10694), .B (n_10697), .Y (n_10698));
NAND3X1 g72761(.A (n_10765), .B (g5046), .C (g5041), .Y (n_10697));
CLKBUFX2 g72769(.A (n_10709), .Y (n_10710));
AND2X1 g72770(.A (n_11065), .B (n_10708), .Y (n_10709));
INVX2 g72771(.A (g_18635), .Y (n_10708));
OAI21X1 g72772(.A0 (g_19913), .A1 (n_9664), .B0 (n_10714), .Y(n_10715));
NAND3X1 g72775(.A (n_10713), .B (n_9651), .C (n_7144), .Y (n_10714));
INVX1 g72776(.A (g_22605), .Y (n_10713));
INVX1 g72777(.A (n_10949), .Y (n_10716));
NAND2X2 g72778(.A (n_10720), .B (n_10976), .Y (n_10874));
NOR2X1 g72780(.A (n_11121), .B (n_8850), .Y (n_10717));
OAI21X1 g72781(.A0 (n_900), .A1 (n_2108), .B0 (g1430), .Y (n_10718));
NOR2X1 g72782(.A (g2629), .B (g2555), .Y (n_10720));
XOR2X1 g72783(.A (g1322), .B (g1339), .Y (n_11077));
CLKBUFX1 g72786(.A (n_10723), .Y (n_10724));
NAND2X1 g72787(.A (n_10505), .B (n_8594), .Y (n_10723));
NAND2X2 g72788(.A (n_1559), .B (n_6762), .Y (n_10725));
XOR2X1 g72806(.A (n_10745), .B (n_10751), .Y (n_10752));
OR4X1 g72807(.A (g_15287), .B (g13259), .C (g19334), .D (n_923), .Y(n_10745));
OR2X1 g72808(.A (n_10750), .B (n_10725), .Y (n_10751));
AOI21X1 g72809(.A0 (n_10123), .A1 (n_10746), .B0 (n_10749), .Y(n_10750));
NOR2X1 g72810(.A (n_10724), .B (g1236), .Y (n_10746));
NOR2X1 g72811(.A (n_10748), .B (n_10123), .Y (n_10749));
NAND2X1 g72812(.A (n_10747), .B (g1236), .Y (n_10748));
INVX1 g72813(.A (n_10724), .Y (n_10747));
NOR2X1 g72814(.A (n_10724), .B (n_10725), .Y (n_10753));
INVX2 g72815(.A (n_10760), .Y (n_10761));
OAI21X1 g72816(.A0 (g1585), .A1 (n_10755), .B0 (n_10759), .Y(n_10760));
CLKBUFX1 g72817(.A (n_10754), .Y (n_10755));
NAND3X1 g72818(.A (n_10201), .B (n_6670), .C (n_10710), .Y (n_10754));
NAND2X2 g72819(.A (n_10758), .B (n_10755), .Y (n_10759));
NAND4X1 g72820(.A (n_10199), .B (n_10756), .C (n_6673), .D (n_10871),.Y (n_10758));
CLKBUFX1 g72821(.A (n_10710), .Y (n_10756));
INVX1 g72823(.A (n_10759), .Y (n_10762));
INVX2 g72824(.A (n_10754), .Y (n_10763));
INVX1 g72825(.A (g1585), .Y (n_10764));
AOI21X1 g72826(.A0 (n_10765), .A1 (g5041), .B0 (n_10769), .Y(n_10770));
NOR2X1 g72827(.A (n_281), .B (n_1493), .Y (n_10765));
INVX1 g72828(.A (n_10768), .Y (n_10769));
NAND2X1 g72829(.A (n_10766), .B (n_10767), .Y (n_10768));
INVX1 g72830(.A (g5041), .Y (n_10766));
NOR2X1 g72831(.A (g5037), .B (n_6970), .Y (n_10767));
INVX1 g72832(.A (n_10767), .Y (n_10771));
INVX1 g72835(.A (n_7219), .Y (n_10772));
NAND2X1 g72836(.A (n_10519), .B (n_7217), .Y (n_10773));
AND2X1 g72839(.A (g34027), .B (n_2385), .Y (n_10781));
INVX1 g72840(.A (n_10949), .Y (n_10782));
NAND2X2 g72843(.A (n_5944), .B (n_10789), .Y (n_10790));
NAND2X2 g72845(.A (n_10785), .B (n_10993), .Y (n_10787));
OAI21X1 g72846(.A0 (n_6893), .A1 (g2819), .B0 (n_8557), .Y (n_10785));
AND2X1 g72848(.A (g2619), .B (g2587), .Y (n_10789));
NAND2X2 g72859(.A (n_10803), .B (g1536), .Y (n_10804));
NAND2X2 g72860(.A (n_10801), .B (n_10802), .Y (n_10803));
INVX1 g14(.A (g1351), .Y (n_10801));
INVX2 g72861(.A (g1312), .Y (n_10802));
NOR2X1 g72862(.A (n_6490), .B (n_6479), .Y (n_10805));
NOR2X1 g69657_dup(.A (n_6490), .B (n_6479), .Y (n_10806));
CLKBUFX1 g72864(.A (n_10809), .Y (n_10808));
INVX1 g72867(.A (n_10814), .Y (n_10813));
INVX1 g72868(.A (g_14843), .Y (n_10814));
INVX1 g72872(.A (n_10823), .Y (n_10818));
CLKBUFX1 g72879(.A (n_10826), .Y (n_10823));
INVX1 g72880(.A (g4776), .Y (n_10826));
INVX1 g72881(.A (n_10829), .Y (n_10827));
INVX1 g72883(.A (n_10831), .Y (n_10830));
CLKBUFX1 g72884(.A (n_10833), .Y (n_10831));
INVX1 g72885(.A (n_10839), .Y (n_10834));
INVX1 g72889(.A (g3288), .Y (n_10839));
INVX1 g72891(.A (n_10846), .Y (n_10841));
INVX1 g72899(.A (g2756), .Y (n_10846));
INVX1 g72901(.A (n_10853), .Y (n_10852));
CLKBUFX3 g72902(.A (n_10854), .Y (n_10853));
CLKBUFX3 g72903(.A (n_10961), .Y (n_10854));
INVX1 g72905(.A (n_10857), .Y (n_10856));
CLKBUFX1 g72906(.A (n_10961), .Y (n_10857));
INVX1 g72908(.A (n_10863), .Y (n_10861));
INVX1 g72910(.A (n_7040), .Y (n_10863));
CLKBUFX1 g72915(.A (n_10871), .Y (n_10867));
INVX1 g72916(.A (n_10874), .Y (n_10873));
INVX1 g72918(.A (n_10879), .Y (n_10877));
INVX2 g72920(.A (n_10573), .Y (n_10879));
INVX2 g72930(.A (n_10894), .Y (n_10889));
INVX1 g72932(.A (n_10894), .Y (n_10893));
INVX2 g72933(.A (n_10883), .Y (n_10894));
INVX2 g72934(.A (n_10883), .Y (n_10895));
INVX4 g72935(.A (n_10897), .Y (n_10883));
INVX2 g72936(.A (n_10898), .Y (n_10897));
INVX2 g72937(.A (g3689), .Y (n_10898));
INVX2 g72938(.A (n_10903), .Y (n_10899));
INVX1 g72940(.A (n_10901), .Y (n_10903));
INVX1 g72941(.A (n_10907), .Y (n_10906));
INVX1 g72942(.A (n_10905), .Y (n_10907));
INVX1 g72943(.A (n_10913), .Y (n_10910));
INVX1 g72944(.A (n_10912), .Y (n_10911));
INVX1 g72945(.A (n_10913), .Y (n_10912));
CLKBUFX3 g72946(.A (n_10915), .Y (n_10913));
INVX1 g72947(.A (n_10917), .Y (n_10916));
INVX2 g72948(.A (n_10915), .Y (n_10917));
CLKBUFX3 g72949(.A (n_10464), .Y (n_10915));
INVX1 g72950(.A (n_10920), .Y (n_10921));
CLKBUFX3 g72951(.A (n_6791), .Y (n_10920));
NAND3X1 g72959(.A (n_10932), .B (n_11033), .C (n_10936), .Y(n_10937));
OAI21X1 g33(.A0 (n_1166), .A1 (n_2108), .B0 (g17404), .Y (n_10932));
NAND2X1 g36_dup(.A (n_10709), .B (n_10203), .Y (n_10934));
NAND3X1 g72962(.A (n_10280), .B (g2704), .C (n_11097), .Y (n_10936));
NAND2X1 g72964(.A (n_10939), .B (n_10943), .Y (n_10944));
AND2X1 g16_dup(.A (g34035), .B (n_10181), .Y (n_10939));
INVX1 g13(.A (n_10942), .Y (n_10943));
NAND2X1 g72965(.A (n_10940), .B (n_10941), .Y (n_10942));
AND2X1 g72966(.A (n_8588), .B (g16624), .Y (n_10940));
AND2X1 g72967(.A (g3288), .B (n_7004), .Y (n_10941));
AND2X1 g16(.A (g34035), .B (n_10181), .Y (n_3249));
NAND2X1 g72968(.A (n_10951), .B (n_10954), .Y (n_10955));
NAND4X1 g72969(.A (n_10772), .B (n_10773), .C (n_10948), .D(n_10950), .Y (n_10951));
INVX1 g72970(.A (n_10947), .Y (n_10948));
NAND2X1 g72971(.A (n_2385), .B (g34027), .Y (n_10947));
CLKBUFX3 g72973(.A (n_10949), .Y (n_10950));
BUFX3 g1(.A (g35), .Y (n_10949));
AOI22X1 g72974(.A0 (n_10952), .A1 (g5467), .B0 (n_10953), .B1(n_10947), .Y (n_10954));
INVX2 g72975(.A (n_10950), .Y (n_10952));
AND2X1 g72976(.A (n_3616), .B (n_9862), .Y (n_10953));
NAND3X1 g72977(.A (n_11035), .B (n_10959), .C (n_10960), .Y(n_10961));
INVX1 g72979(.A (g1291), .Y (n_10956));
NAND2X2 g72980(.A (n_10203), .B (n_10709), .Y (n_11121));
OAI21X1 g72981(.A0 (n_909), .A1 (n_2108), .B0 (g17423), .Y (n_10959));
NAND3X1 g72982(.A (n_169), .B (g2697), .C (n_11097), .Y (n_10960));
NAND4X1 g98(.A (n_10968), .B (n_10972), .C (n_10973), .D (n_1586), .Y(n_10974));
NOR2X1 g99(.A (n_10964), .B (n_10967), .Y (n_10968));
NAND2X1 g101(.A (n_10962), .B (n_10963), .Y (n_10964));
NAND4X1 g107(.A (n_1499), .B (n_11030), .C (g3251), .D (g16603), .Y(n_10962));
NAND4X1 g105(.A (n_8586), .B (n_7383), .C (g3199), .D (g14421), .Y(n_10963));
NAND3X1 g100(.A (n_6948), .B (n_10965), .C (n_10966), .Y (n_10967));
NAND4X1 g104(.A (n_7383), .B (n_10941), .C (g16874), .D (g3223), .Y(n_10965));
NAND4X1 g103(.A (n_8572), .B (n_8587), .C (g16624), .D (g3203), .Y(n_10966));
AOI21X1 g102(.A0 (n_10970), .A1 (n_8572), .B0 (n_10971), .Y(n_10972));
INVX1 g108(.A (n_10969), .Y (n_10970));
NAND3X1 g109(.A (n_7383), .B (g16686), .C (g3255), .Y (n_10969));
NAND2X1 g110(.A (n_8552), .B (n_5501), .Y (n_10971));
NAND4X1 g106(.A (n_11029), .B (n_7383), .C (g3239), .D (g13865), .Y(n_10973));
OAI21X1 g72983(.A0 (n_10975), .A1 (g2629), .B0 (n_10980), .Y(n_10981));
AOI21X1 g72984(.A0 (n_10976), .A1 (n_6742), .B0 (g2555), .Y(n_10975));
NAND2X1 g72985(.A (n_10982), .B (g2555), .Y (n_10980));
CLKBUFX1 g72987(.A (n_10976), .Y (n_10978));
NAND2X2 g72989(.A (n_10718), .B (n_10717), .Y (n_10976));
INVX1 g72990(.A (n_10978), .Y (n_10982));
INVX2 g72991(.A (n_10983), .Y (n_10984));
NAND3X1 g72992(.A (g4849), .B (g4843), .C (n_11216), .Y (n_10983));
INVX1 g72994(.A (g1242), .Y (g23683));
AND2X1 g26_dup72995(.A (n_898), .B (n_10986), .Y (n_10987));
AOI21X1 g72996(.A0 (n_10557), .A1 (g_20563), .B0 (n_10560), .Y(n_10986));
AOI21X1 g72997(.A0 (n_10871), .A1 (n_10986), .B0 (n_10988), .Y(n_10989));
AND2X1 g72998(.A (n_10986), .B (n_898), .Y (n_10988));
OR2X1 g72999(.A (n_10991), .B (n_10994), .Y (n_10995));
NAND2X1 g73000(.A (g2060), .B (g2028), .Y (n_10991));
NAND2X1 g73001(.A (n_10992), .B (n_10993), .Y (n_10994));
OAI21X1 g73002(.A0 (g2787), .A1 (n_6892), .B0 (n_8557), .Y (n_10992));
AND2X1 g73003(.A (n_3679), .B (n_8895), .Y (n_10993));
INVX1 g73004(.A (n_10991), .Y (n_10996));
NOR2X1 g73005(.A (n_11129), .B (n_10997), .Y (n_10998));
INVX2 g73006(.A (g4899), .Y (n_10997));
CLKBUFX1 g73019(.A (n_11013), .Y (n_11012));
NOR2X1 g73027(.A (g1319), .B (n_10200), .Y (n_11025));
NOR2X1 g61156_dup(.A (g1319), .B (n_10200), .Y (n_11026));
NAND2X1 g73028(.A (n_10813), .B (n_6527), .Y (n_11027));
NAND2X1 g10_dup(.A (n_10813), .B (n_6527), .Y (n_11028));
NOR2X1 g73029(.A (n_10834), .B (n_7004), .Y (n_11029));
NOR2X1 g71188_dup(.A (n_10834), .B (n_7004), .Y (n_11030));
AOI21X1 g73030(.A0 (n_2479), .A1 (n_3713), .B0 (n_3718), .Y(n_11031));
AOI21X1 g62838_dup(.A0 (n_2479), .A1 (n_3713), .B0 (n_3718), .Y(n_11032));
AOI21X1 g73031(.A0 (n_10956), .A1 (g1448), .B0 (n_10934), .Y(n_11033));
AOI21X1 g72960_dup(.A0 (n_10956), .A1 (g1448), .B0 (n_10934), .Y(n_11034));
AOI21X1 g73032(.A0 (n_10956), .A1 (g1472), .B0 (n_11121), .Y(n_11035));
AOI21X1 g72978_dup(.A0 (n_10956), .A1 (g1472), .B0 (n_11121), .Y(n_11036));
INVX2 g73033(.A (n_11038), .Y (n_11037));
INVX1 g73034(.A (g5297), .Y (n_11038));
AOI21X1 g73035(.A0 (g23683), .A1 (n_10987), .B0 (n_10989), .Y(n_11039));
AOI21X1 g72993_dup(.A0 (g23683), .A1 (n_10987), .B0 (n_10989), .Y(n_11040));
NOR2X1 g73036(.A (n_11073), .B (n_3459), .Y (n_11041));
NOR2X1 g61208_dup(.A (n_11076), .B (n_3459), .Y (n_11042));
INVX1 g73039(.A (g12350), .Y (n_11045));
CLKBUFX1 g73042(.A (n_11050), .Y (g12350));
INVX1 g73044(.A (n_11064), .Y (n_11051));
INVX1 g73048(.A (n_11055), .Y (n_11056));
CLKBUFX3 g73052(.A (n_11064), .Y (n_11055));
CLKBUFX1 g73055(.A (n_11065), .Y (n_11064));
CLKBUFX1 g73058(.A (n_11071), .Y (n_11070));
CLKBUFX1 g73061(.A (n_11076), .Y (n_11073));
CLKBUFX2 g73062(.A (n_11077), .Y (n_11076));
CLKBUFX1 g73064(.A (n_11081), .Y (n_11080));
INVX2 g73070(.A (n_11088), .Y (g11388));
CLKBUFX1 g73073(.A (n_11091), .Y (n_11088));
INVX1 g73074(.A (g_9298), .Y (n_11091));
CLKBUFX1 g73076(.A (n_11095), .Y (n_11094));
CLKBUFX1 g73079(.A (n_11099), .Y (n_11097));
CLKBUFX1 g73082(.A (n_11105), .Y (n_11104));
INVX1 g73083(.A (n_11110), .Y (n_11106));
INVX1 g73088(.A (g_20244), .Y (n_11110));
CLKBUFX1 g73091(.A (n_11116), .Y (n_11113));
INVX1 g73093(.A (n_11119), .Y (n_11118));
CLKBUFX1 g73094(.A (n_11120), .Y (n_11119));
INVX2 g73095(.A (n_6907), .Y (n_11120));
INVX1 g73096(.A (n_11121), .Y (n_11122));
INVX1 g73097(.A (n_11126), .Y (n_11124));
CLKBUFX2 g73099(.A (n_11128), .Y (n_11126));
INVX1 g73103(.A (n_11134), .Y (n_11133));
CLKBUFX1 g73104(.A (n_11129), .Y (n_11134));
INVX1 g73106(.A (n_11129), .Y (n_11187));
INVX1 g73107(.A (n_8819), .Y (n_11138));
INVX4 g73122(.A (n_11150), .Y (n_11157));
BUFX3 g73124(.A (n_11160), .Y (n_11150));
INVX1 g73125(.A (g6381), .Y (n_11160));
CLKBUFX1 g73127(.A (n_11163), .Y (n_11162));
INVX1 g73128(.A (n_11186), .Y (n_11165));
INVX1 g73135(.A (n_11173), .Y (n_11171));
INVX2 g73137(.A (n_11177), .Y (n_11173));
CLKBUFX3 g73139(.A (n_11185), .Y (n_11177));
INVX1 g73140(.A (n_11184), .Y (n_11178));
CLKBUFX1 g73146(.A (n_11185), .Y (n_11184));
CLKBUFX1 g73147(.A (n_11186), .Y (n_11185));
NOR2X1 g73148(.A (n_10285), .B (n_10290), .Y (n_11190));
NOR2X1 g72378_dup(.A (n_10285), .B (n_10290), .Y (n_11191));
NAND3X1 g73149(.A (n_4206), .B (n_7088), .C (n_11205), .Y (n_11196));
NAND3X1 g70131_dup(.A (n_4206), .B (n_7088), .C (n_11206), .Y(n_11197));
CLKBUFX1 g73153(.A (n_11203), .Y (n_11201));
CLKBUFX1 g73154(.A (n_11198), .Y (n_11203));
NOR2X1 g73155(.A (n_7089), .B (n_7090), .Y (n_11205));
NOR2X1 g70135_dup(.A (n_7089), .B (n_7090), .Y (n_11206));
AOI21X1 g73156(.A0 (n_1564), .A1 (n_1747), .B0 (g4878), .Y (n_11207));
AOI21X1 g64564_dup(.A0 (n_1564), .A1 (n_1747), .B0 (g4878), .Y(n_11208));
NOR2X1 g73157(.A (n_8915), .B (n_10826), .Y (n_11209));
NOR2X1 g71226_dup(.A (n_8915), .B (n_10826), .Y (n_11210));
AND2X1 g73158(.A (n_10960), .B (n_11036), .Y (n_11211));
AND2X1 g70020_dup(.A (n_10960), .B (n_11036), .Y (n_11212));
endmodule
