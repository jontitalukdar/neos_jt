module sha1_exec ( clk, reset, start, data_in, load_in, cv, use_prev_cv, busy,out_valid, cv_next );
input [31:0] data_in;
input [159:0] cv;
output [159:0] cv_next;
input clk, reset, start, load_in, use_prev_cv;
output busy, out_valid;
wire   N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70,N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84,N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,N188, n4654, n4655, n4656, n4658, n4660, n4661, n4662, n4663, n4664,n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,n4715, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,n6096, n6117, n6118, n6139, n6140, n6145, n6146, n6147, n6148, n6149,n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6569,n6570, n6571, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,n6852, n6853, n6856, n6859, n6862, n6865, n6868, n6871, n6874, n6877,n6880, n6883, n6884, n6885, n6886, n6889, n6892, n6895, n6898, n6901,n6904, n6907, n6910, n6913, n6916, n6917, n6918, n6919, n6922, n6925,n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,n7046, n7047, n7048, n7049, n7050, n7052, n7053, n7054, n7055, n7056,n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,n7397, n7398, n7399, n7400, n7401, n7402, n7403, _sha1_round_n825 ,_sha1_round_n824 , _sha1_round_n823 , _sha1_round_n822 ,_sha1_round_n821 , _sha1_round_n820 , _sha1_round_n819 ,_sha1_round_n818 , _sha1_round_n817 , _sha1_round_n816 ,_sha1_round_n815 , _sha1_round_n814 , _sha1_round_n813 ,_sha1_round_n812 , _sha1_round_n811 , _sha1_round_n810 ,_sha1_round_n809 , _sha1_round_n808 , _sha1_round_n807 ,_sha1_round_n806 , _sha1_round_n805 , _sha1_round_n804 ,_sha1_round_n803 , _sha1_round_n802 , _sha1_round_n801 ,_sha1_round_n800 , _sha1_round_n799 , _sha1_round_n798 ,_sha1_round_n797 , _sha1_round_n796 , _sha1_round_n795 ,_sha1_round_n794 , _sha1_round_n793 , _sha1_round_n792 ,_sha1_round_n791 , _sha1_round_n790 , _sha1_round_n789 ,_sha1_round_n788 , _sha1_round_n787 , _sha1_round_n786 ,_sha1_round_n785 , _sha1_round_n784 , _sha1_round_n783 ,_sha1_round_n782 , _sha1_round_n781 , _sha1_round_n780 ,_sha1_round_n779 , _sha1_round_n778 , _sha1_round_n777 ,_sha1_round_n776 , _sha1_round_n775 , _sha1_round_n774 ,_sha1_round_n773 , _sha1_round_n772 , _sha1_round_n771 ,_sha1_round_n770 , _sha1_round_n769 , _sha1_round_n768 ,_sha1_round_n767 , _sha1_round_n766 , _sha1_round_n765 ,_sha1_round_n764 , _sha1_round_n763 , _sha1_round_n762 ,_sha1_round_n761 , _sha1_round_n760 , _sha1_round_n759 ,_sha1_round_n758 , _sha1_round_n757 , _sha1_round_n756 ,_sha1_round_n755 , _sha1_round_n754 , _sha1_round_n753 ,_sha1_round_n752 , _sha1_round_n751 , _sha1_round_n750 ,_sha1_round_n749 , _sha1_round_n748 , _sha1_round_n747 ,_sha1_round_n746 , _sha1_round_n745 , _sha1_round_n744 ,_sha1_round_n743 , _sha1_round_n742 , _sha1_round_n741 ,_sha1_round_n740 , _sha1_round_n739 , _sha1_round_n738 ,_sha1_round_n737 , _sha1_round_n736 , _sha1_round_n735 ,_sha1_round_n734 , _sha1_round_n733 , _sha1_round_n732 ,_sha1_round_n731 , _sha1_round_n730 , _sha1_round_n729 ,_sha1_round_n728 , _sha1_round_n727 , _sha1_round_n726 ,_sha1_round_n725 , _sha1_round_n724 , _sha1_round_n723 ,_sha1_round_n722 , _sha1_round_n721 , _sha1_round_n720 ,_sha1_round_n719 , _sha1_round_n718 , _sha1_round_n717 ,_sha1_round_n716 , _sha1_round_n715 , _sha1_round_n714 ,_sha1_round_n713 , _sha1_round_n712 , _sha1_round_n711 ,_sha1_round_n710 , _sha1_round_n709 , _sha1_round_n708 ,_sha1_round_n707 , _sha1_round_n706 , _sha1_round_n705 ,_sha1_round_n704 , _sha1_round_n703 , _sha1_round_n702 ,_sha1_round_n701 , _sha1_round_n700 , _sha1_round_n699 ,_sha1_round_n698 , _sha1_round_n697 , _sha1_round_n696 ,_sha1_round_n695 , _sha1_round_n694 , _sha1_round_n693 ,_sha1_round_n692 , _sha1_round_n691 , _sha1_round_n690 ,_sha1_round_n689 , _sha1_round_n688 , _sha1_round_n687 ,_sha1_round_n686 , _sha1_round_n685 , _sha1_round_n684 ,_sha1_round_n683 , _sha1_round_n682 , _sha1_round_n681 ,_sha1_round_n680 , _sha1_round_n679 , _sha1_round_n678 ,_sha1_round_n677 , _sha1_round_n676 , _sha1_round_n675 ,_sha1_round_n674 , _sha1_round_n673 , _sha1_round_n672 ,_sha1_round_n671 , _sha1_round_n670 , _sha1_round_n669 ,_sha1_round_n668 , _sha1_round_n667 , _sha1_round_n666 ,_sha1_round_n665 , _sha1_round_n664 , _sha1_round_n663 ,_sha1_round_n662 , _sha1_round_n661 , _sha1_round_n660 ,_sha1_round_n659 , _sha1_round_n658 , _sha1_round_n657 ,_sha1_round_n656 , _sha1_round_n655 , _sha1_round_n654 ,_sha1_round_n653 , _sha1_round_n652 , _sha1_round_n651 ,_sha1_round_n650 , _sha1_round_n649 , _sha1_round_n648 ,_sha1_round_n647 , _sha1_round_n646 , _sha1_round_n645 ,_sha1_round_n644 , _sha1_round_n643 , _sha1_round_n642 ,_sha1_round_n641 , _sha1_round_n640 , _sha1_round_n639 ,_sha1_round_n638 , _sha1_round_n637 , _sha1_round_n636 ,_sha1_round_n635 , _sha1_round_n634 , _sha1_round_n633 ,_sha1_round_n632 , _sha1_round_n631 , _sha1_round_n630 ,_sha1_round_n629 , _sha1_round_n628 , _sha1_round_n627 ,_sha1_round_n626 , _sha1_round_n625 , _sha1_round_n624 ,_sha1_round_n623 , _sha1_round_n622 , _sha1_round_n621 ,_sha1_round_n620 , _sha1_round_n619 , _sha1_round_n618 ,_sha1_round_n617 , _sha1_round_n616 , _sha1_round_n615 ,_sha1_round_n614 , _sha1_round_n613 , _sha1_round_n612 ,_sha1_round_n611 , _sha1_round_n610 , _sha1_round_n609 ,_sha1_round_n608 , _sha1_round_n607 , _sha1_round_n606 ,_sha1_round_n605 , _sha1_round_n604 , _sha1_round_n603 ,_sha1_round_n602 , _sha1_round_n601 , _sha1_round_n600 ,_sha1_round_n599 , _sha1_round_n598 , _sha1_round_n597 ,_sha1_round_n596 , _sha1_round_n595 , _sha1_round_n594 ,_sha1_round_n593 , _sha1_round_n592 , _sha1_round_n591 ,_sha1_round_n590 , _sha1_round_n589 , _sha1_round_n588 ,_sha1_round_n587 , _sha1_round_n586 , _sha1_round_n585 ,_sha1_round_n584 , _sha1_round_n583 , _sha1_round_n582 ,_sha1_round_n581 , _sha1_round_n580 , _sha1_round_n579 ,_sha1_round_n578 , _sha1_round_n577 , _sha1_round_n576 ,_sha1_round_n575 , _sha1_round_n574 , _sha1_round_n573 ,_sha1_round_n572 , _sha1_round_n571 , _sha1_round_n570 ,_sha1_round_n569 , _sha1_round_n568 , _sha1_round_n567 ,_sha1_round_n566 , _sha1_round_n565 , _sha1_round_n564 ,_sha1_round_n563 , _sha1_round_n562 , _sha1_round_n561 ,_sha1_round_n560 , _sha1_round_n559 , _sha1_round_n558 ,_sha1_round_n557 , _sha1_round_n556 , _sha1_round_n555 ,_sha1_round_n554 , _sha1_round_n553 , _sha1_round_n552 ,_sha1_round_n551 , _sha1_round_n550 , _sha1_round_n549 ,_sha1_round_n548 , _sha1_round_n547 , _sha1_round_n546 ,_sha1_round_n545 , _sha1_round_n544 , _sha1_round_n543 ,_sha1_round_n542 , _sha1_round_n541 , _sha1_round_n540 ,_sha1_round_n539 , _sha1_round_n538 , _sha1_round_n537 ,_sha1_round_n536 , _sha1_round_n535 , _sha1_round_n534 ,_sha1_round_n533 , _sha1_round_n532 , _sha1_round_n531 ,_sha1_round_n530 , _sha1_round_n529 , _sha1_round_n528 ,_sha1_round_n527 , _sha1_round_n526 , _sha1_round_n525 ,_sha1_round_n524 , _sha1_round_n523 , _sha1_round_n522 ,_sha1_round_n521 , _sha1_round_n520 , _sha1_round_n519 ,_sha1_round_n518 , _sha1_round_n517 , _sha1_round_n516 ,_sha1_round_n515 , _sha1_round_n514 , _sha1_round_n513 ,_sha1_round_n512 , _sha1_round_n511 , _sha1_round_n510 ,_sha1_round_n509 , _sha1_round_n508 , _sha1_round_n380 ,_sha1_round_n379 , _sha1_round_n378 , _sha1_round_n377 ,_sha1_round_n376 , _sha1_round_n375 , _sha1_round_n374 ,_sha1_round_n373 , _sha1_round_n372 , _sha1_round_n371 ,_sha1_round_n370 , _sha1_round_n369 , _sha1_round_n368 ,_sha1_round_n367 , _sha1_round_n366 , _sha1_round_n365 ,_sha1_round_n364 , _sha1_round_n363 , _sha1_round_n362 ,_sha1_round_n361 , _sha1_round_n360 , _sha1_round_n359 ,_sha1_round_n358 , _sha1_round_n357 , _sha1_round_n356 ,_sha1_round_n355 , _sha1_round_n354 , _sha1_round_n353 ,_sha1_round_n352 , _sha1_round_n351 , _sha1_round_n350 ,_sha1_round_n349 , _sha1_round_n348 , _sha1_round_n3470 ,_sha1_round_n3460 , _sha1_round_n3450 , _sha1_round_n3440 ,_sha1_round_n3430 , _sha1_round_n3420 , _sha1_round_n3410 ,_sha1_round_n3400 , _sha1_round_n3390 , _sha1_round_n3380 ,_sha1_round_n3370 , _sha1_round_n3360 , _sha1_round_n3350 ,_sha1_round_n3340 , _sha1_round_n3330 , _sha1_round_n3320 ,_sha1_round_n3300 , _sha1_round_n3290 , _sha1_round_n3280 ,_sha1_round_n3270 , _sha1_round_n3260 , _sha1_round_n3250 ,_sha1_round_n3240 , _sha1_round_n3230 , _sha1_round_n3220 ,_sha1_round_n3210 , _sha1_round_n3200 , _sha1_round_n3190 ,_sha1_round_n3180 , _sha1_round_n3160 , _sha1_round_n3150 ,_sha1_round_n3140 , _sha1_round_n3130 , _sha1_round_n3120 ,_sha1_round_n3170 , _sha1_round_n168 , _sha1_round_n167 ,_sha1_round_n159 , _sha1_round_n158 , _sha1_round_n150 ,_sha1_round_n149 , _sha1_round_n141 , _sha1_round_n140 ,_sha1_round_n132 , _sha1_round_n131 , _sha1_round_n123 ,_sha1_round_n122 , _sha1_round_n114 , _sha1_round_n113 ,_sha1_round_n96 , _sha1_round_n95 , _sha1_round_n87 ,_sha1_round_n86 , _sha1_round_n2 , _sha1_round_N252 ,_sha1_round_N253 , _sha1_round_N254 , _sha1_round_N255 ,_sha1_round_N256 , _sha1_round_N257 , _sha1_round_N258 ,_sha1_round_N259 , _sha1_round_N260 , _sha1_round_N261 ,_sha1_round_N262 , _sha1_round_N263 , _sha1_round_N264 ,_sha1_round_N265 , _sha1_round_N266 , _sha1_round_N267 ,_sha1_round_N268 , _sha1_round_N269 , _sha1_round_N270 ,_sha1_round_N271 , _sha1_round_N272 , _sha1_round_N273 ,_sha1_round_N274 , _sha1_round_N275 , _sha1_round_N276 ,_sha1_round_N277 , _sha1_round_N278 , _sha1_round_N279 ,_sha1_round_N280 , _sha1_round_N281 , _sha1_round_N282 ,_sha1_round_N283 , _sha1_round_N284 , _sha1_round_N285 ,_sha1_round_N286 , _sha1_round_N287 , _sha1_round_N288 ,_sha1_round_N289 , _sha1_round_N290 , _sha1_round_N291 ,_sha1_round_N292 , _sha1_round_N293 , _sha1_round_N294 ,_sha1_round_N295 , _sha1_round_N296 , _sha1_round_N297 ,_sha1_round_N298 , _sha1_round_N299 , _sha1_round_N300 ,_sha1_round_N301 , _sha1_round_N302 , _sha1_round_N303 ,_sha1_round_N304 , _sha1_round_N305 , _sha1_round_N306 ,_sha1_round_N307 , _sha1_round_N308 , _sha1_round_N309 ,_sha1_round_N310 , _sha1_round_N311 , _sha1_round_N312 ,_sha1_round_N313 , _sha1_round_N314 , _sha1_round_N315 ,_sha1_round_N316 , _sha1_round_N317 , _sha1_round_N318 ,_sha1_round_N319 , _sha1_round_N320 , _sha1_round_N321 ,_sha1_round_N322 , _sha1_round_N323 , _sha1_round_N324 ,_sha1_round_N325 , _sha1_round_N326 , _sha1_round_N327 ,_sha1_round_N328 , _sha1_round_N329 , _sha1_round_N330 ,_sha1_round_N331 , _sha1_round_N332 , _sha1_round_N333 ,_sha1_round_N334 , _sha1_round_N335 , _sha1_round_N336 ,_sha1_round_N337 , _sha1_round_N338 , _sha1_round_N339 ,_sha1_round_N340 , _sha1_round_N341 , _sha1_round_N342 ,_sha1_round_N343 , _sha1_round_N344 , _sha1_round_N345 ,_sha1_round_N346 , _sha1_round_N347 , _sha1_round_k[3] ,_sha1_round_k[13] , _sha1_round_k[15] , _sha1_round_k_23 ,_sha1_round_k_26 , _sha1_round_k_27 , _sha1_round_k_30 ,_sha1_round_add_79_4_n345 , _sha1_round_add_79_4_n344 ,_sha1_round_add_79_4_n343 , _sha1_round_add_79_4_n342 ,_sha1_round_add_79_4_n341 , _sha1_round_add_79_4_n340 ,_sha1_round_add_79_4_n339 , _sha1_round_add_79_4_n338 ,_sha1_round_add_79_4_n337 , _sha1_round_add_79_4_n336 ,_sha1_round_add_79_4_n335 , _sha1_round_add_79_4_n334 ,_sha1_round_add_79_4_n333 , _sha1_round_add_79_4_n332 ,_sha1_round_add_79_4_n331 , _sha1_round_add_79_4_n330 ,_sha1_round_add_79_4_n329 , _sha1_round_add_79_4_n328 ,_sha1_round_add_79_4_n327 , _sha1_round_add_79_4_n326 ,_sha1_round_add_79_4_n325 , _sha1_round_add_79_4_n324 ,_sha1_round_add_79_4_n323 , _sha1_round_add_79_4_n322 ,_sha1_round_add_79_4_n321 , _sha1_round_add_79_4_n320 ,_sha1_round_add_79_4_n319 , _sha1_round_add_79_4_n318 ,_sha1_round_add_79_4_n317 , _sha1_round_add_79_4_n316 ,_sha1_round_add_79_4_n315 , _sha1_round_add_79_4_n314 ,_sha1_round_add_79_4_n313 , _sha1_round_add_79_4_n312 ,_sha1_round_add_79_4_n311 , _sha1_round_add_79_4_n310 ,_sha1_round_add_79_4_n309 , _sha1_round_add_79_4_n308 ,_sha1_round_add_79_4_n307 , _sha1_round_add_79_4_n306 ,_sha1_round_add_79_4_n305 , _sha1_round_add_79_4_n304 ,_sha1_round_add_79_4_n303 , _sha1_round_add_79_4_n302 ,_sha1_round_add_79_4_n301 , _sha1_round_add_79_4_n300 ,_sha1_round_add_79_4_n299 , _sha1_round_add_79_4_n298 ,_sha1_round_add_79_4_n297 , _sha1_round_add_79_4_n296 ,_sha1_round_add_79_4_n295 , _sha1_round_add_79_4_n294 ,_sha1_round_add_79_4_n293 , _sha1_round_add_79_4_n292 ,_sha1_round_add_79_4_n291 , _sha1_round_add_79_4_n290 ,_sha1_round_add_79_4_n289 , _sha1_round_add_79_4_n288 ,_sha1_round_add_79_4_n287 , _sha1_round_add_79_4_n286 ,_sha1_round_add_79_4_n285 , _sha1_round_add_79_4_n284 ,_sha1_round_add_79_4_n283 , _sha1_round_add_79_4_n282 ,_sha1_round_add_79_4_n281 , _sha1_round_add_79_4_n280 ,_sha1_round_add_79_4_n279 , _sha1_round_add_79_4_n278 ,_sha1_round_add_79_4_n277 , _sha1_round_add_79_4_n276 ,_sha1_round_add_79_4_n275 , _sha1_round_add_79_4_n274 ,_sha1_round_add_79_4_n273 , _sha1_round_add_79_4_n272 ,_sha1_round_add_79_4_n271 , _sha1_round_add_79_4_n270 ,_sha1_round_add_79_4_n269 , _sha1_round_add_79_4_n268 ,_sha1_round_add_79_4_n267 , _sha1_round_add_79_4_n266 ,_sha1_round_add_79_4_n265 , _sha1_round_add_79_4_n264 ,_sha1_round_add_79_4_n263 , _sha1_round_add_79_4_n262 ,_sha1_round_add_79_4_n261 , _sha1_round_add_79_4_n260 ,_sha1_round_add_79_4_n259 , _sha1_round_add_79_4_n258 ,_sha1_round_add_79_4_n257 , _sha1_round_add_79_4_n256 ,_sha1_round_add_79_4_n255 , _sha1_round_add_79_4_n254 ,_sha1_round_add_79_4_n253 , _sha1_round_add_79_4_n252 ,_sha1_round_add_79_4_n251 , _sha1_round_add_79_4_n250 ,_sha1_round_add_79_4_n249 , _sha1_round_add_79_4_n248 ,_sha1_round_add_79_4_n247 , _sha1_round_add_79_4_n246 ,_sha1_round_add_79_4_n245 , _sha1_round_add_79_4_n244 ,_sha1_round_add_79_4_n243 , _sha1_round_add_79_4_n242 ,_sha1_round_add_79_4_n241 , _sha1_round_add_79_4_n240 ,_sha1_round_add_79_4_n239 , _sha1_round_add_79_4_n238 ,_sha1_round_add_79_4_n237 , _sha1_round_add_79_4_n236 ,_sha1_round_add_79_4_n235 , _sha1_round_add_79_4_n234 ,_sha1_round_add_79_4_n233 , _sha1_round_add_79_4_n232 ,_sha1_round_add_79_4_n231 , _sha1_round_add_79_4_n230 ,_sha1_round_add_79_4_n229 , _sha1_round_add_79_4_n228 ,_sha1_round_add_79_4_n227 , _sha1_round_add_79_4_n226 ,_sha1_round_add_79_4_n225 , _sha1_round_add_79_4_n224 ,_sha1_round_add_79_4_n223 , _sha1_round_add_79_4_n222 ,_sha1_round_add_79_4_n221 , _sha1_round_add_79_4_n220 ,_sha1_round_add_79_4_n219 , _sha1_round_add_79_4_n218 ,_sha1_round_add_79_4_n217 , _sha1_round_add_79_4_n216 ,_sha1_round_add_79_4_n215 , _sha1_round_add_79_4_n214 ,_sha1_round_add_79_4_n213 , _sha1_round_add_79_4_n212 ,_sha1_round_add_79_4_n211 , _sha1_round_add_79_4_n210 ,_sha1_round_add_79_4_n209 , _sha1_round_add_79_4_n208 ,_sha1_round_add_79_4_n207 , _sha1_round_add_79_4_n206 ,_sha1_round_add_79_4_n205 , _sha1_round_add_79_4_n204 ,_sha1_round_add_79_4_n203 , _sha1_round_add_79_4_n202 ,_sha1_round_add_79_4_n201 , _sha1_round_add_79_4_n200 ,_sha1_round_add_79_4_n199 , _sha1_round_add_79_4_n198 ,_sha1_round_add_79_4_n197 , _sha1_round_add_79_4_n196 ,_sha1_round_add_79_4_n195 , _sha1_round_add_79_4_n194 ,_sha1_round_add_79_4_n193 , _sha1_round_add_79_4_n192 ,_sha1_round_add_79_4_n191 , _sha1_round_add_79_4_n190 ,_sha1_round_add_79_4_n189 , _sha1_round_add_79_4_n188 ,_sha1_round_add_79_4_n187 , _sha1_round_add_79_4_n186 ,_sha1_round_add_79_4_n185 , _sha1_round_add_79_4_n184 ,_sha1_round_add_79_4_n183 , _sha1_round_add_79_4_n182 ,_sha1_round_add_79_4_n181 , _sha1_round_add_79_4_n180 ,_sha1_round_add_79_4_n179 , _sha1_round_add_79_4_n178 ,_sha1_round_add_79_4_n177 , _sha1_round_add_79_4_n176 ,_sha1_round_add_79_4_n175 , _sha1_round_add_79_4_n174 ,_sha1_round_add_79_4_n173 , _sha1_round_add_79_4_n172 ,_sha1_round_add_79_4_n171 , _sha1_round_add_79_4_n170 ,_sha1_round_add_79_4_n169 , _sha1_round_add_79_4_n168 ,_sha1_round_add_79_4_n167 , _sha1_round_add_79_4_n166 ,_sha1_round_add_79_4_n165 , _sha1_round_add_79_4_n164 ,_sha1_round_add_79_4_n163 , _sha1_round_add_79_4_n162 ,_sha1_round_add_79_4_n161 , _sha1_round_add_79_4_n160 ,_sha1_round_add_79_4_n159 , _sha1_round_add_79_4_n158 ,_sha1_round_add_79_4_n157 , _sha1_round_add_79_4_n156 ,_sha1_round_add_79_4_n155 , _sha1_round_add_79_4_n154 ,_sha1_round_add_79_4_n153 , _sha1_round_add_79_4_n152 ,_sha1_round_add_79_4_n151 , _sha1_round_add_79_4_n150 ,_sha1_round_add_79_4_n149 , _sha1_round_add_79_4_n148 ,_sha1_round_add_79_4_n147 , _sha1_round_add_79_4_n146 ,_sha1_round_add_79_4_n145 , _sha1_round_add_79_4_n144 ,_sha1_round_add_79_4_n143 , _sha1_round_add_79_4_n142 ,_sha1_round_add_79_4_n141 , _sha1_round_add_79_4_n140 ,_sha1_round_add_79_4_n139 , _sha1_round_add_79_4_n138 ,_sha1_round_add_79_4_n137 , _sha1_round_add_79_4_n136 ,_sha1_round_add_79_4_n135 , _sha1_round_add_79_4_n134 ,_sha1_round_add_79_4_n133 , _sha1_round_add_79_4_n132 ,_sha1_round_add_79_4_n131 , _sha1_round_add_79_4_n130 ,_sha1_round_add_79_4_n129 , _sha1_round_add_79_4_n128 ,_sha1_round_add_79_4_n127 , _sha1_round_add_79_4_n126 ,_sha1_round_add_79_4_n125 , _sha1_round_add_79_4_n124 ,_sha1_round_add_79_4_n123 , _sha1_round_add_79_4_n122 ,_sha1_round_add_79_4_n121 , _sha1_round_add_79_4_n120 ,_sha1_round_add_79_4_n119 , _sha1_round_add_79_4_n118 ,_sha1_round_add_79_4_n117 , _sha1_round_add_79_4_n116 ,_sha1_round_add_79_4_n115 , _sha1_round_add_79_4_n114 ,_sha1_round_add_79_4_n113 , _sha1_round_add_79_4_n112 ,_sha1_round_add_79_4_n111 , _sha1_round_add_79_4_n110 ,_sha1_round_add_79_4_n109 , _sha1_round_add_79_4_n108 ,_sha1_round_add_79_4_n107 , _sha1_round_add_79_4_n106 ,_sha1_round_add_79_4_n105 , _sha1_round_add_79_4_n104 ,_sha1_round_add_79_4_n103 , _sha1_round_add_79_4_n102 ,_sha1_round_add_79_4_n101 , _sha1_round_add_79_4_n100 ,_sha1_round_add_79_4_n99 , _sha1_round_add_79_4_n98 ,_sha1_round_add_79_4_n97 , _sha1_round_add_79_4_n96 ,_sha1_round_add_79_4_n95 , _sha1_round_add_79_4_n94 ,_sha1_round_add_79_4_n93 , _sha1_round_add_79_4_n92 ,_sha1_round_add_79_4_n91 , _sha1_round_add_79_4_n90 ,_sha1_round_add_79_4_n89 , _sha1_round_add_79_4_n88 ,_sha1_round_add_79_4_n87 , _sha1_round_add_79_4_n86 ,_sha1_round_add_79_4_n85 , _sha1_round_add_79_4_n84 ,_sha1_round_add_79_4_n83 , _sha1_round_add_79_4_n82 ,_sha1_round_add_79_4_n81 , _sha1_round_add_79_4_n80 ,_sha1_round_add_79_4_n79 , _sha1_round_add_79_4_n78 ,_sha1_round_add_79_4_n77 , _sha1_round_add_79_4_n76 ,_sha1_round_add_79_4_n75 , _sha1_round_add_79_4_n74 ,_sha1_round_add_79_4_n73 , _sha1_round_add_79_4_n72 ,_sha1_round_add_79_4_n71 , _sha1_round_add_79_4_n70 ,_sha1_round_add_79_4_n69 , _sha1_round_add_79_4_n68 ,_sha1_round_add_79_4_n67 , _sha1_round_add_79_4_n66 ,_sha1_round_add_79_4_n65 , _sha1_round_add_79_4_n64 ,_sha1_round_add_79_4_n63 , _sha1_round_add_79_4_n62 ,_sha1_round_add_79_4_n61 , _sha1_round_add_79_4_n60 ,_sha1_round_add_79_4_n59 , _sha1_round_add_79_4_n58 ,_sha1_round_add_79_4_n57 , _sha1_round_add_79_4_n56 ,_sha1_round_add_79_4_n55 , _sha1_round_add_79_4_n54 ,_sha1_round_add_79_4_n53 , _sha1_round_add_79_4_n52 ,_sha1_round_add_79_4_n51 , _sha1_round_add_79_4_n50 ,_sha1_round_add_79_4_n49 , _sha1_round_add_79_4_n48 ,_sha1_round_add_79_4_n47 , _sha1_round_add_79_4_n46 ,_sha1_round_add_79_4_n45 , _sha1_round_add_79_4_n44 ,_sha1_round_add_79_4_n43 , _sha1_round_add_79_4_n42 ,_sha1_round_add_79_4_n41 , _sha1_round_add_79_4_n40 ,_sha1_round_add_79_4_n39 , _sha1_round_add_79_4_n38 ,_sha1_round_add_79_4_n37 , _sha1_round_add_79_4_n36 ,_sha1_round_add_79_4_n35 , _sha1_round_add_79_4_n34 ,_sha1_round_add_79_4_n33 , _sha1_round_add_79_4_n32 ,_sha1_round_add_79_4_n31 , _sha1_round_add_79_4_n30 ,_sha1_round_add_79_4_n29 , _sha1_round_add_79_4_n28 ,_sha1_round_add_79_4_n27 , _sha1_round_add_79_4_n26 ,_sha1_round_add_79_4_n25 , _sha1_round_add_79_4_n24 ,_sha1_round_add_79_4_n23 , _sha1_round_add_79_4_n22 ,_sha1_round_add_79_4_n21 , _sha1_round_add_79_4_n20 ,_sha1_round_add_79_4_n19 , _sha1_round_add_79_4_n18 ,_sha1_round_add_79_4_n17 , _sha1_round_add_79_4_n15 ,_sha1_round_add_79_4_n14 , _sha1_round_add_79_4_n13 ,_sha1_round_add_79_4_n12 , _sha1_round_add_79_4_n11 ,_sha1_round_add_79_4_n10 , _sha1_round_add_79_4_n9 ,_sha1_round_add_79_4_n8 , _sha1_round_add_79_4_n7 ,_sha1_round_add_79_4_n6 , _sha1_round_add_79_4_n5 ,_sha1_round_add_79_4_n4 , _sha1_round_add_79_4_n3 ,_sha1_round_add_79_4_n2 , _sha1_round_add_79_4_n1 ,_sha1_round_add_79_3_n387 , _sha1_round_add_79_3_n386 ,_sha1_round_add_79_3_n385 , _sha1_round_add_79_3_n384 ,_sha1_round_add_79_3_n383 , _sha1_round_add_79_3_n382 ,_sha1_round_add_79_3_n381 , _sha1_round_add_79_3_n380 ,_sha1_round_add_79_3_n379 , _sha1_round_add_79_3_n378 ,_sha1_round_add_79_3_n377 , _sha1_round_add_79_3_n376 ,_sha1_round_add_79_3_n375 , _sha1_round_add_79_3_n374 ,_sha1_round_add_79_3_n373 , _sha1_round_add_79_3_n372 ,_sha1_round_add_79_3_n371 , _sha1_round_add_79_3_n370 ,_sha1_round_add_79_3_n369 , _sha1_round_add_79_3_n368 ,_sha1_round_add_79_3_n367 , _sha1_round_add_79_3_n366 ,_sha1_round_add_79_3_n365 , _sha1_round_add_79_3_n364 ,_sha1_round_add_79_3_n363 , _sha1_round_add_79_3_n362 ,_sha1_round_add_79_3_n361 , _sha1_round_add_79_3_n360 ,_sha1_round_add_79_3_n359 , _sha1_round_add_79_3_n358 ,_sha1_round_add_79_3_n357 , _sha1_round_add_79_3_n356 ,_sha1_round_add_79_3_n355 , _sha1_round_add_79_3_n354 ,_sha1_round_add_79_3_n353 , _sha1_round_add_79_3_n352 ,_sha1_round_add_79_3_n351 , _sha1_round_add_79_3_n350 ,_sha1_round_add_79_3_n349 , _sha1_round_add_79_3_n348 ,_sha1_round_add_79_3_n347 , _sha1_round_add_79_3_n346 ,_sha1_round_add_79_3_n345 , _sha1_round_add_79_3_n344 ,_sha1_round_add_79_3_n343 , _sha1_round_add_79_3_n342 ,_sha1_round_add_79_3_n341 , _sha1_round_add_79_3_n340 ,_sha1_round_add_79_3_n339 , _sha1_round_add_79_3_n338 ,_sha1_round_add_79_3_n337 , _sha1_round_add_79_3_n336 ,_sha1_round_add_79_3_n335 , _sha1_round_add_79_3_n334 ,_sha1_round_add_79_3_n333 , _sha1_round_add_79_3_n332 ,_sha1_round_add_79_3_n331 , _sha1_round_add_79_3_n330 ,_sha1_round_add_79_3_n329 , _sha1_round_add_79_3_n328 ,_sha1_round_add_79_3_n327 , _sha1_round_add_79_3_n326 ,_sha1_round_add_79_3_n325 , _sha1_round_add_79_3_n324 ,_sha1_round_add_79_3_n323 , _sha1_round_add_79_3_n322 ,_sha1_round_add_79_3_n321 , _sha1_round_add_79_3_n320 ,_sha1_round_add_79_3_n319 , _sha1_round_add_79_3_n318 ,_sha1_round_add_79_3_n317 , _sha1_round_add_79_3_n316 ,_sha1_round_add_79_3_n315 , _sha1_round_add_79_3_n314 ,_sha1_round_add_79_3_n313 , _sha1_round_add_79_3_n312 ,_sha1_round_add_79_3_n311 , _sha1_round_add_79_3_n310 ,_sha1_round_add_79_3_n309 , _sha1_round_add_79_3_n308 ,_sha1_round_add_79_3_n307 , _sha1_round_add_79_3_n306 ,_sha1_round_add_79_3_n305 , _sha1_round_add_79_3_n304 ,_sha1_round_add_79_3_n303 , _sha1_round_add_79_3_n302 ,_sha1_round_add_79_3_n301 , _sha1_round_add_79_3_n300 ,_sha1_round_add_79_3_n299 , _sha1_round_add_79_3_n298 ,_sha1_round_add_79_3_n297 , _sha1_round_add_79_3_n296 ,_sha1_round_add_79_3_n295 , _sha1_round_add_79_3_n294 ,_sha1_round_add_79_3_n293 , _sha1_round_add_79_3_n292 ,_sha1_round_add_79_3_n291 , _sha1_round_add_79_3_n290 ,_sha1_round_add_79_3_n289 , _sha1_round_add_79_3_n288 ,_sha1_round_add_79_3_n287 , _sha1_round_add_79_3_n286 ,_sha1_round_add_79_3_n285 , _sha1_round_add_79_3_n284 ,_sha1_round_add_79_3_n283 , _sha1_round_add_79_3_n282 ,_sha1_round_add_79_3_n281 , _sha1_round_add_79_3_n280 ,_sha1_round_add_79_3_n279 , _sha1_round_add_79_3_n278 ,_sha1_round_add_79_3_n277 , _sha1_round_add_79_3_n276 ,_sha1_round_add_79_3_n275 , _sha1_round_add_79_3_n274 ,_sha1_round_add_79_3_n273 , _sha1_round_add_79_3_n272 ,_sha1_round_add_79_3_n271 , _sha1_round_add_79_3_n270 ,_sha1_round_add_79_3_n269 , _sha1_round_add_79_3_n268 ,_sha1_round_add_79_3_n267 , _sha1_round_add_79_3_n266 ,_sha1_round_add_79_3_n265 , _sha1_round_add_79_3_n264 ,_sha1_round_add_79_3_n263 , _sha1_round_add_79_3_n262 ,_sha1_round_add_79_3_n261 , _sha1_round_add_79_3_n260 ,_sha1_round_add_79_3_n259 , _sha1_round_add_79_3_n258 ,_sha1_round_add_79_3_n257 , _sha1_round_add_79_3_n256 ,_sha1_round_add_79_3_n255 , _sha1_round_add_79_3_n254 ,_sha1_round_add_79_3_n253 , _sha1_round_add_79_3_n252 ,_sha1_round_add_79_3_n251 , _sha1_round_add_79_3_n250 ,_sha1_round_add_79_3_n249 , _sha1_round_add_79_3_n248 ,_sha1_round_add_79_3_n247 , _sha1_round_add_79_3_n246 ,_sha1_round_add_79_3_n245 , _sha1_round_add_79_3_n244 ,_sha1_round_add_79_3_n243 , _sha1_round_add_79_3_n242 ,_sha1_round_add_79_3_n241 , _sha1_round_add_79_3_n240 ,_sha1_round_add_79_3_n239 , _sha1_round_add_79_3_n238 ,_sha1_round_add_79_3_n237 , _sha1_round_add_79_3_n236 ,_sha1_round_add_79_3_n235 , _sha1_round_add_79_3_n234 ,_sha1_round_add_79_3_n233 , _sha1_round_add_79_3_n232 ,_sha1_round_add_79_3_n231 , _sha1_round_add_79_3_n230 ,_sha1_round_add_79_3_n229 , _sha1_round_add_79_3_n228 ,_sha1_round_add_79_3_n227 , _sha1_round_add_79_3_n226 ,_sha1_round_add_79_3_n225 , _sha1_round_add_79_3_n224 ,_sha1_round_add_79_3_n223 , _sha1_round_add_79_3_n222 ,_sha1_round_add_79_3_n221 , _sha1_round_add_79_3_n220 ,_sha1_round_add_79_3_n219 , _sha1_round_add_79_3_n218 ,_sha1_round_add_79_3_n217 , _sha1_round_add_79_3_n216 ,_sha1_round_add_79_3_n215 , _sha1_round_add_79_3_n214 ,_sha1_round_add_79_3_n213 , _sha1_round_add_79_3_n212 ,_sha1_round_add_79_3_n211 , _sha1_round_add_79_3_n210 ,_sha1_round_add_79_3_n209 , _sha1_round_add_79_3_n208 ,_sha1_round_add_79_3_n207 , _sha1_round_add_79_3_n206 ,_sha1_round_add_79_3_n205 , _sha1_round_add_79_3_n204 ,_sha1_round_add_79_3_n203 , _sha1_round_add_79_3_n202 ,_sha1_round_add_79_3_n201 , _sha1_round_add_79_3_n200 ,_sha1_round_add_79_3_n199 , _sha1_round_add_79_3_n198 ,_sha1_round_add_79_3_n197 , _sha1_round_add_79_3_n196 ,_sha1_round_add_79_3_n195 , _sha1_round_add_79_3_n194 ,_sha1_round_add_79_3_n193 , _sha1_round_add_79_3_n192 ,_sha1_round_add_79_3_n191 , _sha1_round_add_79_3_n190 ,_sha1_round_add_79_3_n189 , _sha1_round_add_79_3_n188 ,_sha1_round_add_79_3_n187 , _sha1_round_add_79_3_n186 ,_sha1_round_add_79_3_n185 , _sha1_round_add_79_3_n184 ,_sha1_round_add_79_3_n183 , _sha1_round_add_79_3_n182 ,_sha1_round_add_79_3_n181 , _sha1_round_add_79_3_n180 ,_sha1_round_add_79_3_n179 , _sha1_round_add_79_3_n178 ,_sha1_round_add_79_3_n177 , _sha1_round_add_79_3_n176 ,_sha1_round_add_79_3_n175 , _sha1_round_add_79_3_n174 ,_sha1_round_add_79_3_n173 , _sha1_round_add_79_3_n172 ,_sha1_round_add_79_3_n171 , _sha1_round_add_79_3_n170 ,_sha1_round_add_79_3_n169 , _sha1_round_add_79_3_n168 ,_sha1_round_add_79_3_n167 , _sha1_round_add_79_3_n166 ,_sha1_round_add_79_3_n165 , _sha1_round_add_79_3_n164 ,_sha1_round_add_79_3_n163 , _sha1_round_add_79_3_n162 ,_sha1_round_add_79_3_n161 , _sha1_round_add_79_3_n160 ,_sha1_round_add_79_3_n159 , _sha1_round_add_79_3_n158 ,_sha1_round_add_79_3_n157 , _sha1_round_add_79_3_n156 ,_sha1_round_add_79_3_n155 , _sha1_round_add_79_3_n154 ,_sha1_round_add_79_3_n153 , _sha1_round_add_79_3_n152 ,_sha1_round_add_79_3_n151 , _sha1_round_add_79_3_n150 ,_sha1_round_add_79_3_n149 , _sha1_round_add_79_3_n148 ,_sha1_round_add_79_3_n147 , _sha1_round_add_79_3_n146 ,_sha1_round_add_79_3_n145 , _sha1_round_add_79_3_n144 ,_sha1_round_add_79_3_n143 , _sha1_round_add_79_3_n142 ,_sha1_round_add_79_3_n141 , _sha1_round_add_79_3_n140 ,_sha1_round_add_79_3_n139 , _sha1_round_add_79_3_n138 ,_sha1_round_add_79_3_n137 , _sha1_round_add_79_3_n136 ,_sha1_round_add_79_3_n135 , _sha1_round_add_79_3_n134 ,_sha1_round_add_79_3_n133 , _sha1_round_add_79_3_n132 ,_sha1_round_add_79_3_n131 , _sha1_round_add_79_3_n130 ,_sha1_round_add_79_3_n129 , _sha1_round_add_79_3_n128 ,_sha1_round_add_79_3_n127 , _sha1_round_add_79_3_n126 ,_sha1_round_add_79_3_n125 , _sha1_round_add_79_3_n124 ,_sha1_round_add_79_3_n123 , _sha1_round_add_79_3_n122 ,_sha1_round_add_79_3_n121 , _sha1_round_add_79_3_n120 ,_sha1_round_add_79_3_n119 , _sha1_round_add_79_3_n118 ,_sha1_round_add_79_3_n117 , _sha1_round_add_79_3_n116 ,_sha1_round_add_79_3_n115 , _sha1_round_add_79_3_n114 ,_sha1_round_add_79_3_n113 , _sha1_round_add_79_3_n112 ,_sha1_round_add_79_3_n111 , _sha1_round_add_79_3_n110 ,_sha1_round_add_79_3_n109 , _sha1_round_add_79_3_n108 ,_sha1_round_add_79_3_n107 , _sha1_round_add_79_3_n106 ,_sha1_round_add_79_3_n105 , _sha1_round_add_79_3_n104 ,_sha1_round_add_79_3_n103 , _sha1_round_add_79_3_n102 ,_sha1_round_add_79_3_n101 , _sha1_round_add_79_3_n100 ,_sha1_round_add_79_3_n99 , _sha1_round_add_79_3_n98 ,_sha1_round_add_79_3_n97 , _sha1_round_add_79_3_n96 ,_sha1_round_add_79_3_n95 , _sha1_round_add_79_3_n94 ,_sha1_round_add_79_3_n93 , _sha1_round_add_79_3_n92 ,_sha1_round_add_79_3_n91 , _sha1_round_add_79_3_n90 ,_sha1_round_add_79_3_n89 , _sha1_round_add_79_3_n88 ,_sha1_round_add_79_3_n87 , _sha1_round_add_79_3_n86 ,_sha1_round_add_79_3_n85 , _sha1_round_add_79_3_n84 ,_sha1_round_add_79_3_n83 , _sha1_round_add_79_3_n82 ,_sha1_round_add_79_3_n81 , _sha1_round_add_79_3_n80 ,_sha1_round_add_79_3_n79 , _sha1_round_add_79_3_n78 ,_sha1_round_add_79_3_n77 , _sha1_round_add_79_3_n76 ,_sha1_round_add_79_3_n75 , _sha1_round_add_79_3_n74 ,_sha1_round_add_79_3_n73 , _sha1_round_add_79_3_n72 ,_sha1_round_add_79_3_n71 , _sha1_round_add_79_3_n70 ,_sha1_round_add_79_3_n69 , _sha1_round_add_79_3_n68 ,_sha1_round_add_79_3_n67 , _sha1_round_add_79_3_n66 ,_sha1_round_add_79_3_n65 , _sha1_round_add_79_3_n64 ,_sha1_round_add_79_3_n63 , _sha1_round_add_79_3_n62 ,_sha1_round_add_79_3_n61 , _sha1_round_add_79_3_n60 ,_sha1_round_add_79_3_n58 , _sha1_round_add_79_3_n57 ,_sha1_round_add_79_3_n56 , _sha1_round_add_79_3_n55 ,_sha1_round_add_79_3_n54 , _sha1_round_add_79_3_n53 ,_sha1_round_add_79_3_n52 , _sha1_round_add_79_3_n51 ,_sha1_round_add_79_3_n50 , _sha1_round_add_79_3_n49 ,_sha1_round_add_79_3_n48 , _sha1_round_add_79_3_n47 ,_sha1_round_add_79_3_n46 , _sha1_round_add_79_3_n45 ,_sha1_round_add_79_3_n44 , _sha1_round_add_79_3_n43 ,_sha1_round_add_79_3_n42 , _sha1_round_add_79_3_n41 ,_sha1_round_add_79_3_n40 , _sha1_round_add_79_3_n39 ,_sha1_round_add_79_3_n38 , _sha1_round_add_79_3_n37 ,_sha1_round_add_79_3_n36 , _sha1_round_add_79_3_n35 ,_sha1_round_add_79_3_n34 , _sha1_round_add_79_3_n33 ,_sha1_round_add_79_3_n32 , _sha1_round_add_79_3_n31 ,_sha1_round_add_79_3_n30 , _sha1_round_add_79_3_n29 ,_sha1_round_add_79_3_n28 , _sha1_round_add_79_3_n27 ,_sha1_round_add_79_3_n26 , _sha1_round_add_79_3_n25 ,_sha1_round_add_79_3_n24 , _sha1_round_add_79_3_n23 ,_sha1_round_add_79_3_n22 , _sha1_round_add_79_3_n21 ,_sha1_round_add_79_3_n20 , _sha1_round_add_79_3_n19 ,_sha1_round_add_79_3_n18 , _sha1_round_add_79_3_n17 ,_sha1_round_add_79_3_n16 , _sha1_round_add_79_3_n15 ,_sha1_round_add_79_3_n14 , _sha1_round_add_79_3_n13 ,_sha1_round_add_79_3_n12 , _sha1_round_add_79_3_n11 ,_sha1_round_add_79_3_n10 , _sha1_round_add_79_3_n9 ,_sha1_round_add_79_3_n8 , _sha1_round_add_79_3_n7 ,_sha1_round_add_79_3_n6 , _sha1_round_add_79_3_n5 ,_sha1_round_add_79_3_n4 , _sha1_round_add_79_3_n3 ,_sha1_round_add_79_3_n1 , _sha1_round_add_79_n381 ,_sha1_round_add_79_n380 , _sha1_round_add_79_n379 ,_sha1_round_add_79_n378 , _sha1_round_add_79_n377 ,_sha1_round_add_79_n376 , _sha1_round_add_79_n375 ,_sha1_round_add_79_n374 , _sha1_round_add_79_n373 ,_sha1_round_add_79_n372 , _sha1_round_add_79_n371 ,_sha1_round_add_79_n370 , _sha1_round_add_79_n369 ,_sha1_round_add_79_n368 , _sha1_round_add_79_n367 ,_sha1_round_add_79_n366 , _sha1_round_add_79_n365 ,_sha1_round_add_79_n364 , _sha1_round_add_79_n363 ,_sha1_round_add_79_n362 , _sha1_round_add_79_n361 ,_sha1_round_add_79_n360 , _sha1_round_add_79_n359 ,_sha1_round_add_79_n358 , _sha1_round_add_79_n357 ,_sha1_round_add_79_n356 , _sha1_round_add_79_n355 ,_sha1_round_add_79_n354 , _sha1_round_add_79_n353 ,_sha1_round_add_79_n352 , _sha1_round_add_79_n351 ,_sha1_round_add_79_n350 , _sha1_round_add_79_n349 ,_sha1_round_add_79_n348 , _sha1_round_add_79_n347 ,_sha1_round_add_79_n346 , _sha1_round_add_79_n345 ,_sha1_round_add_79_n344 , _sha1_round_add_79_n343 ,_sha1_round_add_79_n342 , _sha1_round_add_79_n341 ,_sha1_round_add_79_n340 , _sha1_round_add_79_n339 ,_sha1_round_add_79_n338 , _sha1_round_add_79_n337 ,_sha1_round_add_79_n336 , _sha1_round_add_79_n335 ,_sha1_round_add_79_n334 , _sha1_round_add_79_n333 ,_sha1_round_add_79_n332 , _sha1_round_add_79_n331 ,_sha1_round_add_79_n330 , _sha1_round_add_79_n329 ,_sha1_round_add_79_n328 , _sha1_round_add_79_n327 ,_sha1_round_add_79_n326 , _sha1_round_add_79_n325 ,_sha1_round_add_79_n324 , _sha1_round_add_79_n323 ,_sha1_round_add_79_n322 , _sha1_round_add_79_n321 ,_sha1_round_add_79_n320 , _sha1_round_add_79_n319 ,_sha1_round_add_79_n318 , _sha1_round_add_79_n317 ,_sha1_round_add_79_n316 , _sha1_round_add_79_n315 ,_sha1_round_add_79_n314 , _sha1_round_add_79_n313 ,_sha1_round_add_79_n312 , _sha1_round_add_79_n311 ,_sha1_round_add_79_n310 , _sha1_round_add_79_n309 ,_sha1_round_add_79_n308 , _sha1_round_add_79_n307 ,_sha1_round_add_79_n306 , _sha1_round_add_79_n305 ,_sha1_round_add_79_n304 , _sha1_round_add_79_n303 ,_sha1_round_add_79_n302 , _sha1_round_add_79_n301 ,_sha1_round_add_79_n300 , _sha1_round_add_79_n299 ,_sha1_round_add_79_n298 , _sha1_round_add_79_n297 ,_sha1_round_add_79_n296 , _sha1_round_add_79_n295 ,_sha1_round_add_79_n294 , _sha1_round_add_79_n293 ,_sha1_round_add_79_n292 , _sha1_round_add_79_n291 ,_sha1_round_add_79_n290 , _sha1_round_add_79_n289 ,_sha1_round_add_79_n288 , _sha1_round_add_79_n287 ,_sha1_round_add_79_n286 , _sha1_round_add_79_n285 ,_sha1_round_add_79_n284 , _sha1_round_add_79_n283 ,_sha1_round_add_79_n282 , _sha1_round_add_79_n281 ,_sha1_round_add_79_n280 , _sha1_round_add_79_n279 ,_sha1_round_add_79_n278 , _sha1_round_add_79_n277 ,_sha1_round_add_79_n276 , _sha1_round_add_79_n275 ,_sha1_round_add_79_n274 , _sha1_round_add_79_n273 ,_sha1_round_add_79_n272 , _sha1_round_add_79_n271 ,_sha1_round_add_79_n270 , _sha1_round_add_79_n269 ,_sha1_round_add_79_n268 , _sha1_round_add_79_n267 ,_sha1_round_add_79_n266 , _sha1_round_add_79_n265 ,_sha1_round_add_79_n264 , _sha1_round_add_79_n263 ,_sha1_round_add_79_n262 , _sha1_round_add_79_n261 ,_sha1_round_add_79_n260 , _sha1_round_add_79_n259 ,_sha1_round_add_79_n258 , _sha1_round_add_79_n257 ,_sha1_round_add_79_n256 , _sha1_round_add_79_n255 ,_sha1_round_add_79_n254 , _sha1_round_add_79_n253 ,_sha1_round_add_79_n252 , _sha1_round_add_79_n251 ,_sha1_round_add_79_n250 , _sha1_round_add_79_n249 ,_sha1_round_add_79_n248 , _sha1_round_add_79_n247 ,_sha1_round_add_79_n246 , _sha1_round_add_79_n245 ,_sha1_round_add_79_n244 , _sha1_round_add_79_n243 ,_sha1_round_add_79_n242 , _sha1_round_add_79_n241 ,_sha1_round_add_79_n240 , _sha1_round_add_79_n239 ,_sha1_round_add_79_n238 , _sha1_round_add_79_n237 ,_sha1_round_add_79_n236 , _sha1_round_add_79_n235 ,_sha1_round_add_79_n234 , _sha1_round_add_79_n233 ,_sha1_round_add_79_n232 , _sha1_round_add_79_n231 ,_sha1_round_add_79_n230 , _sha1_round_add_79_n229 ,_sha1_round_add_79_n228 , _sha1_round_add_79_n227 ,_sha1_round_add_79_n226 , _sha1_round_add_79_n225 ,_sha1_round_add_79_n224 , _sha1_round_add_79_n223 ,_sha1_round_add_79_n222 , _sha1_round_add_79_n221 ,_sha1_round_add_79_n220 , _sha1_round_add_79_n219 ,_sha1_round_add_79_n218 , _sha1_round_add_79_n217 ,_sha1_round_add_79_n216 , _sha1_round_add_79_n215 ,_sha1_round_add_79_n214 , _sha1_round_add_79_n213 ,_sha1_round_add_79_n212 , _sha1_round_add_79_n211 ,_sha1_round_add_79_n210 , _sha1_round_add_79_n209 ,_sha1_round_add_79_n208 , _sha1_round_add_79_n207 ,_sha1_round_add_79_n206 , _sha1_round_add_79_n205 ,_sha1_round_add_79_n204 , _sha1_round_add_79_n203 ,_sha1_round_add_79_n202 , _sha1_round_add_79_n201 ,_sha1_round_add_79_n200 , _sha1_round_add_79_n199 ,_sha1_round_add_79_n198 , _sha1_round_add_79_n197 ,_sha1_round_add_79_n196 , _sha1_round_add_79_n195 ,_sha1_round_add_79_n194 , _sha1_round_add_79_n193 ,_sha1_round_add_79_n192 , _sha1_round_add_79_n191 ,_sha1_round_add_79_n190 , _sha1_round_add_79_n189 ,_sha1_round_add_79_n188 , _sha1_round_add_79_n187 ,_sha1_round_add_79_n186 , _sha1_round_add_79_n185 ,_sha1_round_add_79_n184 , _sha1_round_add_79_n183 ,_sha1_round_add_79_n182 , _sha1_round_add_79_n181 ,_sha1_round_add_79_n180 , _sha1_round_add_79_n179 ,_sha1_round_add_79_n178 , _sha1_round_add_79_n177 ,_sha1_round_add_79_n176 , _sha1_round_add_79_n175 ,_sha1_round_add_79_n174 , _sha1_round_add_79_n173 ,_sha1_round_add_79_n172 , _sha1_round_add_79_n171 ,_sha1_round_add_79_n170 , _sha1_round_add_79_n169 ,_sha1_round_add_79_n168 , _sha1_round_add_79_n167 ,_sha1_round_add_79_n166 , _sha1_round_add_79_n165 ,_sha1_round_add_79_n164 , _sha1_round_add_79_n163 ,_sha1_round_add_79_n162 , _sha1_round_add_79_n161 ,_sha1_round_add_79_n160 , _sha1_round_add_79_n159 ,_sha1_round_add_79_n158 , _sha1_round_add_79_n157 ,_sha1_round_add_79_n156 , _sha1_round_add_79_n155 ,_sha1_round_add_79_n154 , _sha1_round_add_79_n153 ,_sha1_round_add_79_n152 , _sha1_round_add_79_n151 ,_sha1_round_add_79_n150 , _sha1_round_add_79_n149 ,_sha1_round_add_79_n148 , _sha1_round_add_79_n147 ,_sha1_round_add_79_n146 , _sha1_round_add_79_n145 ,_sha1_round_add_79_n144 , _sha1_round_add_79_n143 ,_sha1_round_add_79_n142 , _sha1_round_add_79_n141 ,_sha1_round_add_79_n140 , _sha1_round_add_79_n139 ,_sha1_round_add_79_n138 , _sha1_round_add_79_n137 ,_sha1_round_add_79_n136 , _sha1_round_add_79_n135 ,_sha1_round_add_79_n134 , _sha1_round_add_79_n133 ,_sha1_round_add_79_n132 , _sha1_round_add_79_n131 ,_sha1_round_add_79_n130 , _sha1_round_add_79_n129 ,_sha1_round_add_79_n128 , _sha1_round_add_79_n127 ,_sha1_round_add_79_n126 , _sha1_round_add_79_n125 ,_sha1_round_add_79_n124 , _sha1_round_add_79_n123 ,_sha1_round_add_79_n122 , _sha1_round_add_79_n121 ,_sha1_round_add_79_n120 , _sha1_round_add_79_n119 ,_sha1_round_add_79_n118 , _sha1_round_add_79_n117 ,_sha1_round_add_79_n116 , _sha1_round_add_79_n115 ,_sha1_round_add_79_n114 , _sha1_round_add_79_n113 ,_sha1_round_add_79_n112 , _sha1_round_add_79_n111 ,_sha1_round_add_79_n110 , _sha1_round_add_79_n109 ,_sha1_round_add_79_n108 , _sha1_round_add_79_n107 ,_sha1_round_add_79_n106 , _sha1_round_add_79_n105 ,_sha1_round_add_79_n104 , _sha1_round_add_79_n103 ,_sha1_round_add_79_n102 , _sha1_round_add_79_n101 ,_sha1_round_add_79_n100 , _sha1_round_add_79_n99 ,_sha1_round_add_79_n98 , _sha1_round_add_79_n97 ,_sha1_round_add_79_n96 , _sha1_round_add_79_n95 ,_sha1_round_add_79_n94 , _sha1_round_add_79_n93 ,_sha1_round_add_79_n92 , _sha1_round_add_79_n91 ,_sha1_round_add_79_n90 , _sha1_round_add_79_n89 ,_sha1_round_add_79_n88 , _sha1_round_add_79_n87 ,_sha1_round_add_79_n86 , _sha1_round_add_79_n85 ,_sha1_round_add_79_n84 , _sha1_round_add_79_n83 ,_sha1_round_add_79_n82 , _sha1_round_add_79_n81 ,_sha1_round_add_79_n80 , _sha1_round_add_79_n79 ,_sha1_round_add_79_n78 , _sha1_round_add_79_n77 ,_sha1_round_add_79_n75 , _sha1_round_add_79_n74 ,_sha1_round_add_79_n73 , _sha1_round_add_79_n71 ,_sha1_round_add_79_n70 , _sha1_round_add_79_n69 ,_sha1_round_add_79_n68 , _sha1_round_add_79_n67 ,_sha1_round_add_79_n64 , _sha1_round_add_79_n63 ,_sha1_round_add_79_n62 , _sha1_round_add_79_n61 ,_sha1_round_add_79_n60 , _sha1_round_add_79_n59 ,_sha1_round_add_79_n58 , _sha1_round_add_79_n57 ,_sha1_round_add_79_n56 , _sha1_round_add_79_n55 ,_sha1_round_add_79_n54 , _sha1_round_add_79_n53 ,_sha1_round_add_79_n52 , _sha1_round_add_79_n51 ,_sha1_round_add_79_n50 , _sha1_round_add_79_n49 ,_sha1_round_add_79_n48 , _sha1_round_add_79_n47 ,_sha1_round_add_79_n46 , _sha1_round_add_79_n45 ,_sha1_round_add_79_n44 , _sha1_round_add_79_n43 ,_sha1_round_add_79_n42 , _sha1_round_add_79_n41 ,_sha1_round_add_79_n40 , _sha1_round_add_79_n39 ,_sha1_round_add_79_n38 , _sha1_round_add_79_n37 ,_sha1_round_add_79_n36 , _sha1_round_add_79_n35 ,_sha1_round_add_79_n34 , _sha1_round_add_79_n33 ,_sha1_round_add_79_n32 , _sha1_round_add_79_n31 ,_sha1_round_add_79_n30 , _sha1_round_add_79_n29 ,_sha1_round_add_79_n28 , _sha1_round_add_79_n27 ,_sha1_round_add_79_n26 , _sha1_round_add_79_n25 ,_sha1_round_add_79_n24 , _sha1_round_add_79_n23 ,_sha1_round_add_79_n22 , _sha1_round_add_79_n21 ,_sha1_round_add_79_n20 , _sha1_round_add_79_n19 ,_sha1_round_add_79_n18 , _sha1_round_add_79_n17 ,_sha1_round_add_79_n16 , _sha1_round_add_79_n15 ,_sha1_round_add_79_n14 , _sha1_round_add_79_n13 ,_sha1_round_add_79_n12 , _sha1_round_add_79_n11 ,_sha1_round_add_79_n8 , _sha1_round_add_79_n5 ,_sha1_round_add_79_n4 , _sha1_round_add_79_n2 ,_sha1_round_add_79_n1 , _sha1_round_add_79_2_n374 ,_sha1_round_add_79_2_n373 , _sha1_round_add_79_2_n372 ,_sha1_round_add_79_2_n371 , _sha1_round_add_79_2_n370 ,_sha1_round_add_79_2_n369 , _sha1_round_add_79_2_n368 ,_sha1_round_add_79_2_n367 , _sha1_round_add_79_2_n366 ,_sha1_round_add_79_2_n365 , _sha1_round_add_79_2_n364 ,_sha1_round_add_79_2_n363 , _sha1_round_add_79_2_n362 ,_sha1_round_add_79_2_n361 , _sha1_round_add_79_2_n360 ,_sha1_round_add_79_2_n359 , _sha1_round_add_79_2_n358 ,_sha1_round_add_79_2_n357 , _sha1_round_add_79_2_n356 ,_sha1_round_add_79_2_n355 , _sha1_round_add_79_2_n354 ,_sha1_round_add_79_2_n353 , _sha1_round_add_79_2_n352 ,_sha1_round_add_79_2_n351 , _sha1_round_add_79_2_n350 ,_sha1_round_add_79_2_n349 , _sha1_round_add_79_2_n348 ,_sha1_round_add_79_2_n347 , _sha1_round_add_79_2_n346 ,_sha1_round_add_79_2_n345 , _sha1_round_add_79_2_n344 ,_sha1_round_add_79_2_n343 , _sha1_round_add_79_2_n342 ,_sha1_round_add_79_2_n341 , _sha1_round_add_79_2_n340 ,_sha1_round_add_79_2_n339 , _sha1_round_add_79_2_n338 ,_sha1_round_add_79_2_n337 , _sha1_round_add_79_2_n336 ,_sha1_round_add_79_2_n335 , _sha1_round_add_79_2_n334 ,_sha1_round_add_79_2_n333 , _sha1_round_add_79_2_n332 ,_sha1_round_add_79_2_n331 , _sha1_round_add_79_2_n330 ,_sha1_round_add_79_2_n329 , _sha1_round_add_79_2_n328 ,_sha1_round_add_79_2_n327 , _sha1_round_add_79_2_n326 ,_sha1_round_add_79_2_n325 , _sha1_round_add_79_2_n324 ,_sha1_round_add_79_2_n323 , _sha1_round_add_79_2_n322 ,_sha1_round_add_79_2_n321 , _sha1_round_add_79_2_n320 ,_sha1_round_add_79_2_n319 , _sha1_round_add_79_2_n318 ,_sha1_round_add_79_2_n317 , _sha1_round_add_79_2_n316 ,_sha1_round_add_79_2_n315 , _sha1_round_add_79_2_n314 ,_sha1_round_add_79_2_n313 , _sha1_round_add_79_2_n312 ,_sha1_round_add_79_2_n311 , _sha1_round_add_79_2_n310 ,_sha1_round_add_79_2_n309 , _sha1_round_add_79_2_n308 ,_sha1_round_add_79_2_n307 , _sha1_round_add_79_2_n306 ,_sha1_round_add_79_2_n305 , _sha1_round_add_79_2_n304 ,_sha1_round_add_79_2_n303 , _sha1_round_add_79_2_n302 ,_sha1_round_add_79_2_n301 , _sha1_round_add_79_2_n300 ,_sha1_round_add_79_2_n299 , _sha1_round_add_79_2_n298 ,_sha1_round_add_79_2_n297 , _sha1_round_add_79_2_n296 ,_sha1_round_add_79_2_n295 , _sha1_round_add_79_2_n294 ,_sha1_round_add_79_2_n293 , _sha1_round_add_79_2_n292 ,_sha1_round_add_79_2_n291 , _sha1_round_add_79_2_n290 ,_sha1_round_add_79_2_n289 , _sha1_round_add_79_2_n288 ,_sha1_round_add_79_2_n287 , _sha1_round_add_79_2_n286 ,_sha1_round_add_79_2_n285 , _sha1_round_add_79_2_n284 ,_sha1_round_add_79_2_n283 , _sha1_round_add_79_2_n282 ,_sha1_round_add_79_2_n281 , _sha1_round_add_79_2_n280 ,_sha1_round_add_79_2_n279 , _sha1_round_add_79_2_n278 ,_sha1_round_add_79_2_n277 , _sha1_round_add_79_2_n276 ,_sha1_round_add_79_2_n275 , _sha1_round_add_79_2_n274 ,_sha1_round_add_79_2_n273 , _sha1_round_add_79_2_n272 ,_sha1_round_add_79_2_n271 , _sha1_round_add_79_2_n270 ,_sha1_round_add_79_2_n269 , _sha1_round_add_79_2_n268 ,_sha1_round_add_79_2_n267 , _sha1_round_add_79_2_n266 ,_sha1_round_add_79_2_n265 , _sha1_round_add_79_2_n264 ,_sha1_round_add_79_2_n263 , _sha1_round_add_79_2_n262 ,_sha1_round_add_79_2_n261 , _sha1_round_add_79_2_n260 ,_sha1_round_add_79_2_n259 , _sha1_round_add_79_2_n258 ,_sha1_round_add_79_2_n257 , _sha1_round_add_79_2_n256 ,_sha1_round_add_79_2_n255 , _sha1_round_add_79_2_n254 ,_sha1_round_add_79_2_n253 , _sha1_round_add_79_2_n252 ,_sha1_round_add_79_2_n251 , _sha1_round_add_79_2_n250 ,_sha1_round_add_79_2_n249 , _sha1_round_add_79_2_n248 ,_sha1_round_add_79_2_n247 , _sha1_round_add_79_2_n246 ,_sha1_round_add_79_2_n245 , _sha1_round_add_79_2_n244 ,_sha1_round_add_79_2_n243 , _sha1_round_add_79_2_n242 ,_sha1_round_add_79_2_n241 , _sha1_round_add_79_2_n240 ,_sha1_round_add_79_2_n239 , _sha1_round_add_79_2_n238 ,_sha1_round_add_79_2_n237 , _sha1_round_add_79_2_n236 ,_sha1_round_add_79_2_n235 , _sha1_round_add_79_2_n234 ,_sha1_round_add_79_2_n233 , _sha1_round_add_79_2_n232 ,_sha1_round_add_79_2_n231 , _sha1_round_add_79_2_n230 ,_sha1_round_add_79_2_n229 , _sha1_round_add_79_2_n228 ,_sha1_round_add_79_2_n227 , _sha1_round_add_79_2_n226 ,_sha1_round_add_79_2_n225 , _sha1_round_add_79_2_n224 ,_sha1_round_add_79_2_n223 , _sha1_round_add_79_2_n222 ,_sha1_round_add_79_2_n221 , _sha1_round_add_79_2_n220 ,_sha1_round_add_79_2_n219 , _sha1_round_add_79_2_n218 ,_sha1_round_add_79_2_n217 , _sha1_round_add_79_2_n216 ,_sha1_round_add_79_2_n215 , _sha1_round_add_79_2_n214 ,_sha1_round_add_79_2_n213 , _sha1_round_add_79_2_n212 ,_sha1_round_add_79_2_n211 , _sha1_round_add_79_2_n210 ,_sha1_round_add_79_2_n209 , _sha1_round_add_79_2_n208 ,_sha1_round_add_79_2_n207 , _sha1_round_add_79_2_n206 ,_sha1_round_add_79_2_n205 , _sha1_round_add_79_2_n204 ,_sha1_round_add_79_2_n203 , _sha1_round_add_79_2_n202 ,_sha1_round_add_79_2_n201 , _sha1_round_add_79_2_n200 ,_sha1_round_add_79_2_n199 , _sha1_round_add_79_2_n198 ,_sha1_round_add_79_2_n197 , _sha1_round_add_79_2_n196 ,_sha1_round_add_79_2_n195 , _sha1_round_add_79_2_n194 ,_sha1_round_add_79_2_n193 , _sha1_round_add_79_2_n192 ,_sha1_round_add_79_2_n191 , _sha1_round_add_79_2_n190 ,_sha1_round_add_79_2_n189 , _sha1_round_add_79_2_n188 ,_sha1_round_add_79_2_n187 , _sha1_round_add_79_2_n186 ,_sha1_round_add_79_2_n185 , _sha1_round_add_79_2_n184 ,_sha1_round_add_79_2_n183 , _sha1_round_add_79_2_n182 ,_sha1_round_add_79_2_n181 , _sha1_round_add_79_2_n180 ,_sha1_round_add_79_2_n179 , _sha1_round_add_79_2_n178 ,_sha1_round_add_79_2_n177 , _sha1_round_add_79_2_n176 ,_sha1_round_add_79_2_n175 , _sha1_round_add_79_2_n174 ,_sha1_round_add_79_2_n173 , _sha1_round_add_79_2_n172 ,_sha1_round_add_79_2_n171 , _sha1_round_add_79_2_n170 ,_sha1_round_add_79_2_n169 , _sha1_round_add_79_2_n168 ,_sha1_round_add_79_2_n167 , _sha1_round_add_79_2_n166 ,_sha1_round_add_79_2_n165 , _sha1_round_add_79_2_n164 ,_sha1_round_add_79_2_n163 , _sha1_round_add_79_2_n162 ,_sha1_round_add_79_2_n161 , _sha1_round_add_79_2_n160 ,_sha1_round_add_79_2_n159 , _sha1_round_add_79_2_n158 ,_sha1_round_add_79_2_n157 , _sha1_round_add_79_2_n156 ,_sha1_round_add_79_2_n155 , _sha1_round_add_79_2_n154 ,_sha1_round_add_79_2_n153 , _sha1_round_add_79_2_n152 ,_sha1_round_add_79_2_n151 , _sha1_round_add_79_2_n150 ,_sha1_round_add_79_2_n149 , _sha1_round_add_79_2_n148 ,_sha1_round_add_79_2_n147 , _sha1_round_add_79_2_n146 ,_sha1_round_add_79_2_n145 , _sha1_round_add_79_2_n144 ,_sha1_round_add_79_2_n143 , _sha1_round_add_79_2_n142 ,_sha1_round_add_79_2_n141 , _sha1_round_add_79_2_n140 ,_sha1_round_add_79_2_n139 , _sha1_round_add_79_2_n138 ,_sha1_round_add_79_2_n137 , _sha1_round_add_79_2_n136 ,_sha1_round_add_79_2_n135 , _sha1_round_add_79_2_n134 ,_sha1_round_add_79_2_n133 , _sha1_round_add_79_2_n132 ,_sha1_round_add_79_2_n131 , _sha1_round_add_79_2_n130 ,_sha1_round_add_79_2_n129 , _sha1_round_add_79_2_n128 ,_sha1_round_add_79_2_n127 , _sha1_round_add_79_2_n126 ,_sha1_round_add_79_2_n125 , _sha1_round_add_79_2_n124 ,_sha1_round_add_79_2_n123 , _sha1_round_add_79_2_n122 ,_sha1_round_add_79_2_n121 , _sha1_round_add_79_2_n120 ,_sha1_round_add_79_2_n119 , _sha1_round_add_79_2_n118 ,_sha1_round_add_79_2_n117 , _sha1_round_add_79_2_n116 ,_sha1_round_add_79_2_n115 , _sha1_round_add_79_2_n114 ,_sha1_round_add_79_2_n113 , _sha1_round_add_79_2_n112 ,_sha1_round_add_79_2_n111 , _sha1_round_add_79_2_n110 ,_sha1_round_add_79_2_n109 , _sha1_round_add_79_2_n108 ,_sha1_round_add_79_2_n107 , _sha1_round_add_79_2_n106 ,_sha1_round_add_79_2_n105 , _sha1_round_add_79_2_n104 ,_sha1_round_add_79_2_n103 , _sha1_round_add_79_2_n102 ,_sha1_round_add_79_2_n101 , _sha1_round_add_79_2_n100 ,_sha1_round_add_79_2_n99 , _sha1_round_add_79_2_n98 ,_sha1_round_add_79_2_n97 , _sha1_round_add_79_2_n96 ,_sha1_round_add_79_2_n95 , _sha1_round_add_79_2_n94 ,_sha1_round_add_79_2_n93 , _sha1_round_add_79_2_n92 ,_sha1_round_add_79_2_n91 , _sha1_round_add_79_2_n90 ,_sha1_round_add_79_2_n89 , _sha1_round_add_79_2_n88 ,_sha1_round_add_79_2_n87 , _sha1_round_add_79_2_n86 ,_sha1_round_add_79_2_n85 , _sha1_round_add_79_2_n84 ,_sha1_round_add_79_2_n83 , _sha1_round_add_79_2_n82 ,_sha1_round_add_79_2_n81 , _sha1_round_add_79_2_n80 ,_sha1_round_add_79_2_n79 , _sha1_round_add_79_2_n78 ,_sha1_round_add_79_2_n77 , _sha1_round_add_79_2_n76 ,_sha1_round_add_79_2_n75 , _sha1_round_add_79_2_n74 ,_sha1_round_add_79_2_n73 , _sha1_round_add_79_2_n72 ,_sha1_round_add_79_2_n71 , _sha1_round_add_79_2_n70 ,_sha1_round_add_79_2_n69 , _sha1_round_add_79_2_n68 ,_sha1_round_add_79_2_n67 , _sha1_round_add_79_2_n66 ,_sha1_round_add_79_2_n65 , _sha1_round_add_79_2_n64 ,_sha1_round_add_79_2_n63 , _sha1_round_add_79_2_n62 ,_sha1_round_add_79_2_n61 , _sha1_round_add_79_2_n60 ,_sha1_round_add_79_2_n59 , _sha1_round_add_79_2_n58 ,_sha1_round_add_79_2_n57 , _sha1_round_add_79_2_n56 ,_sha1_round_add_79_2_n55 , _sha1_round_add_79_2_n54 ,_sha1_round_add_79_2_n53 , _sha1_round_add_79_2_n52 ,_sha1_round_add_79_2_n51 , _sha1_round_add_79_2_n50 ,_sha1_round_add_79_2_n49 , _sha1_round_add_79_2_n48 ,_sha1_round_add_79_2_n47 , _sha1_round_add_79_2_n46 ,_sha1_round_add_79_2_n45 , _sha1_round_add_79_2_n44 ,_sha1_round_add_79_2_n43 , _sha1_round_add_79_2_n42 ,_sha1_round_add_79_2_n41 , _sha1_round_add_79_2_n40 ,_sha1_round_add_79_2_n39 , _sha1_round_add_79_2_n38 ,_sha1_round_add_79_2_n37 , _sha1_round_add_79_2_n36 ,_sha1_round_add_79_2_n35 , _sha1_round_add_79_2_n34 ,_sha1_round_add_79_2_n33 , _sha1_round_add_79_2_n32 ,_sha1_round_add_79_2_n31 , _sha1_round_add_79_2_n29 ,_sha1_round_add_79_2_n28 , _sha1_round_add_79_2_n27 ,_sha1_round_add_79_2_n25 , _sha1_round_add_79_2_n24 ,_sha1_round_add_79_2_n23 , _sha1_round_add_79_2_n22 ,_sha1_round_add_79_2_n21 , _sha1_round_add_79_2_n20 ,_sha1_round_add_79_2_n19 , _sha1_round_add_79_2_n18 ,_sha1_round_add_79_2_n17 , _sha1_round_add_79_2_n16 ,_sha1_round_add_79_2_n15 , _sha1_round_add_79_2_n14 ,_sha1_round_add_79_2_n13 , _sha1_round_add_79_2_n12 ,_sha1_round_add_79_2_n11 , _sha1_round_add_79_2_n10 ,_sha1_round_add_79_2_n9 , _sha1_round_add_79_2_n8 ,_sha1_round_add_79_2_n7 , _sha1_round_add_79_2_n6 ,_sha1_round_add_79_2_n5 , _sha1_round_add_79_2_n4 ,_sha1_round_add_79_2_n3 , _sha1_round_add_79_2_n2 ,_sha1_round_add_79_2_n1 , _rnd_cnt_reg_n12 , _rnd_cnt_reg_n10 ,_rnd_cnt_reg_n70 , _rnd_cnt_reg_n60 , _rnd_cnt_reg_n40 ,_rnd_cnt_reg_n2 , _rnd_cnt_reg_N9 , _rnd_cnt_reg_N8 ,_rnd_cnt_reg_N7 , _rnd_cnt_reg_N6 , _rnd_cnt_reg_N5 ,_rnd_cnt_reg_N4 , _rnd_cnt_reg_N3 , _state_reg_n2 , _state_reg_N4 ,_state_reg_N3 , _w_reg_n1070 , _w_reg_n1060 , _w_reg_n1050 ,_w_reg_n1040 , _w_reg_n1030 , _w_reg_n1020 , _w_reg_n1010 ,_w_reg_n1000 , _w_reg_n990 , _w_reg_n980 , _w_reg_n970 , _w_reg_n960 ,_w_reg_n950 , _w_reg_n940 , _w_reg_n930 , _w_reg_n920 , _w_reg_n910 ,_w_reg_n900 , _w_reg_n890 , _w_reg_n880 , _w_reg_n870 , _w_reg_n860 ,_w_reg_n850 , _w_reg_n840 , _w_reg_n830 , _w_reg_n820 , _w_reg_n810 ,_w_reg_n800 , _w_reg_n790 , _w_reg_n780 , _w_reg_n770 , _w_reg_n760 ,_w_reg_n750 , _w_reg_n740 , _w_reg_n730 , _w_reg_n720 , _w_reg_n710 ,_w_reg_n700 , _w_reg_n690 , _w_reg_n680 , _w_reg_n670 , _w_reg_n660 ,_w_reg_n650 , _w_reg_n640 , _w_reg_n630 , _w_reg_n620 , _w_reg_n610 ,_w_reg_n600 , _w_reg_N514 , _w_reg_N513 , _w_reg_N512 , _w_reg_N511 ,_w_reg_N510 , _w_reg_N509 , _w_reg_N508 , _w_reg_N507 , _w_reg_N506 ,_w_reg_N505 , _w_reg_N504 , _w_reg_N503 , _w_reg_N502 , _w_reg_N501 ,_w_reg_N500 , _w_reg_N499 , _w_reg_N498 , _w_reg_N497 , _w_reg_N496 ,_w_reg_N495 , _w_reg_N494 , _w_reg_N493 , _w_reg_N492 , _w_reg_N491 ,_w_reg_N490 , _w_reg_N489 , _w_reg_N488 , _w_reg_N487 , _w_reg_N486 ,_w_reg_N485 , _w_reg_N484 , _w_reg_N483 , _w_reg_N482 , _w_reg_N481 ,_w_reg_N480 , _w_reg_N479 , _w_reg_N478 , _w_reg_N477 , _w_reg_N476 ,_w_reg_N475 , _w_reg_N474 , _w_reg_N473 , _w_reg_N472 , _w_reg_N471 ,_w_reg_N470 , _w_reg_N469 , _w_reg_N468 , _w_reg_N467 , _w_reg_N466 ,_w_reg_N465 , _w_reg_N464 , _w_reg_N463 , _w_reg_N462 , _w_reg_N461 ,_w_reg_N460 , _w_reg_N459 , _w_reg_N458 , _w_reg_N457 , _w_reg_N456 ,_w_reg_N455 , _w_reg_N454 , _w_reg_N453 , _w_reg_N452 , _w_reg_N451 ,_w_reg_N450 , _w_reg_N449 , _w_reg_N448 , _w_reg_N447 , _w_reg_N446 ,_w_reg_N445 , _w_reg_N444 , _w_reg_N443 , _w_reg_N442 , _w_reg_N441 ,_w_reg_N440 , _w_reg_N439 , _w_reg_N438 , _w_reg_N437 , _w_reg_N436 ,_w_reg_N435 , _w_reg_N434 , _w_reg_N433 , _w_reg_N432 , _w_reg_N431 ,_w_reg_N430 , _w_reg_N429 , _w_reg_N428 , _w_reg_N427 , _w_reg_N426 ,_w_reg_N425 , _w_reg_N424 , _w_reg_N423 , _w_reg_N422 , _w_reg_N421 ,_w_reg_N420 , _w_reg_N419 , _w_reg_N418 , _w_reg_N417 , _w_reg_N416 ,_w_reg_N415 , _w_reg_N414 , _w_reg_N413 , _w_reg_N412 , _w_reg_N411 ,_w_reg_N410 , _w_reg_N409 , _w_reg_N408 , _w_reg_N407 , _w_reg_N406 ,_w_reg_N405 , _w_reg_N404 , _w_reg_N403 , _w_reg_N402 , _w_reg_N401 ,_w_reg_N400 , _w_reg_N399 , _w_reg_N398 , _w_reg_N397 , _w_reg_N396 ,_w_reg_N395 , _w_reg_N394 , _w_reg_N393 , _w_reg_N392 , _w_reg_N391 ,_w_reg_N390 , _w_reg_N389 , _w_reg_N388 , _w_reg_N387 , _w_reg_N386 ,_w_reg_N385 , _w_reg_N384 , _w_reg_N383 , _w_reg_N382 , _w_reg_N381 ,_w_reg_N380 , _w_reg_N379 , _w_reg_N378 , _w_reg_N377 , _w_reg_N376 ,_w_reg_N375 , _w_reg_N374 , _w_reg_N373 , _w_reg_N372 , _w_reg_N371 ,_w_reg_N370 , _w_reg_N369 , _w_reg_N368 , _w_reg_N367 , _w_reg_N366 ,_w_reg_N365 , _w_reg_N364 , _w_reg_N363 , _w_reg_N362 , _w_reg_N361 ,_w_reg_N360 , _w_reg_N359 , _w_reg_N358 , _w_reg_N357 , _w_reg_N356 ,_w_reg_N355 , _w_reg_N354 , _w_reg_N353 , _w_reg_N352 , _w_reg_N351 ,_w_reg_N350 , _w_reg_N349 , _w_reg_N348 , _w_reg_N347 , _w_reg_N346 ,_w_reg_N345 , _w_reg_N344 , _w_reg_N343 , _w_reg_N342 , _w_reg_N341 ,_w_reg_N340 , _w_reg_N339 , _w_reg_N338 , _w_reg_N337 , _w_reg_N336 ,_w_reg_N335 , _w_reg_N334 , _w_reg_N333 , _w_reg_N332 , _w_reg_N331 ,_w_reg_N330 , _w_reg_N329 , _w_reg_N328 , _w_reg_N327 , _w_reg_N326 ,_w_reg_N325 , _w_reg_N324 , _w_reg_N323 , _w_reg_N322 , _w_reg_N321 ,_w_reg_N320 , _w_reg_N319 , _w_reg_N318 , _w_reg_N317 , _w_reg_N316 ,_w_reg_N315 , _w_reg_N314 , _w_reg_N313 , _w_reg_N312 , _w_reg_N311 ,_w_reg_N310 , _w_reg_N309 , _w_reg_N308 , _w_reg_N307 , _w_reg_N306 ,_w_reg_N305 , _w_reg_N304 , _w_reg_N303 , _w_reg_N302 , _w_reg_N301 ,_w_reg_N300 , _w_reg_N299 , _w_reg_N298 , _w_reg_N297 , _w_reg_N296 ,_w_reg_N295 , _w_reg_N294 , _w_reg_N293 , _w_reg_N292 , _w_reg_N291 ,_w_reg_N290 , _w_reg_N289 , _w_reg_N288 , _w_reg_N287 , _w_reg_N286 ,_w_reg_N285 , _w_reg_N284 , _w_reg_N283 , _w_reg_N282 , _w_reg_N281 ,_w_reg_N280 , _w_reg_N279 , _w_reg_N278 , _w_reg_N277 , _w_reg_N276 ,_w_reg_N275 , _w_reg_N274 , _w_reg_N273 , _w_reg_N272 , _w_reg_N271 ,_w_reg_N270 , _w_reg_N269 , _w_reg_N268 , _w_reg_N267 , _w_reg_N266 ,_w_reg_N265 , _w_reg_N264 , _w_reg_N263 , _w_reg_N262 , _w_reg_N261 ,_w_reg_N260 , _w_reg_N259 , _w_reg_N258 , _w_reg_N257 , _w_reg_N256 ,_w_reg_N255 , _w_reg_N254 , _w_reg_N253 , _w_reg_N252 , _w_reg_N251 ,_w_reg_N250 , _w_reg_N249 , _w_reg_N248 , _w_reg_N247 , _w_reg_N246 ,_w_reg_N245 , _w_reg_N244 , _w_reg_N243 , _w_reg_N242 , _w_reg_N241 ,_w_reg_N240 , _w_reg_N239 , _w_reg_N238 , _w_reg_N237 , _w_reg_N236 ,_w_reg_N235 , _w_reg_N234 , _w_reg_N233 , _w_reg_N232 , _w_reg_N231 ,_w_reg_N230 , _w_reg_N229 , _w_reg_N228 , _w_reg_N227 , _w_reg_N226 ,_w_reg_N225 , _w_reg_N224 , _w_reg_N223 , _w_reg_N222 , _w_reg_N221 ,_w_reg_N220 , _w_reg_N219 , _w_reg_N218 , _w_reg_N217 , _w_reg_N216 ,_w_reg_N215 , _w_reg_N214 , _w_reg_N213 , _w_reg_N212 , _w_reg_N211 ,_w_reg_N210 , _w_reg_N209 , _w_reg_N208 , _w_reg_N207 , _w_reg_N206 ,_w_reg_N205 , _w_reg_N204 , _w_reg_N203 , _w_reg_N202 , _w_reg_N201 ,_w_reg_N200 , _w_reg_N199 , _w_reg_N198 , _w_reg_N197 , _w_reg_N196 ,_w_reg_N195 , _w_reg_N194 , _w_reg_N193 , _w_reg_N192 , _w_reg_N191 ,_w_reg_N190 , _w_reg_N189 , _w_reg_N188 , _w_reg_N187 , _w_reg_N186 ,_w_reg_N185 , _w_reg_N184 , _w_reg_N183 , _w_reg_N182 , _w_reg_N181 ,_w_reg_N180 , _w_reg_N179 , _w_reg_N178 , _w_reg_N177 , _w_reg_N176 ,_w_reg_N175 , _w_reg_N174 , _w_reg_N173 , _w_reg_N172 , _w_reg_N171 ,_w_reg_N170 , _w_reg_N169 , _w_reg_N168 , _w_reg_N167 , _w_reg_N166 ,_w_reg_N165 , _w_reg_N164 , _w_reg_N163 , _w_reg_N162 , _w_reg_N161 ,_w_reg_N160 , _w_reg_N159 , _w_reg_N158 , _w_reg_N157 , _w_reg_N156 ,_w_reg_N155 , _w_reg_N154 , _w_reg_N153 , _w_reg_N152 , _w_reg_N151 ,_w_reg_N150 , _w_reg_N149 , _w_reg_N148 , _w_reg_N147 , _w_reg_N146 ,_w_reg_N145 , _w_reg_N144 , _w_reg_N143 , _w_reg_N142 , _w_reg_N141 ,_w_reg_N140 , _w_reg_N139 , _w_reg_N138 , _w_reg_N137 , _w_reg_N136 ,_w_reg_N135 , _w_reg_N134 , _w_reg_N133 , _w_reg_N132 , _w_reg_N131 ,_w_reg_N130 , _w_reg_N129 , _w_reg_N128 , _w_reg_N127 , _w_reg_N126 ,_w_reg_N125 , _w_reg_N124 , _w_reg_N123 , _w_reg_N122 , _w_reg_N121 ,_w_reg_N120 , _w_reg_N119 , _w_reg_N118 , _w_reg_N117 , _w_reg_N116 ,_w_reg_N115 , _w_reg_N114 , _w_reg_N113 , _w_reg_N112 , _w_reg_N111 ,_w_reg_N110 , _w_reg_N109 , _w_reg_N108 , _w_reg_N107 , _w_reg_N106 ,_w_reg_N105 , _w_reg_N104 , _w_reg_N103 , _w_reg_N102 , _w_reg_N101 ,_w_reg_N100 , _w_reg_N99 , _w_reg_N98 , _w_reg_N97 , _w_reg_N96 ,_w_reg_N95 , _w_reg_N94 , _w_reg_N93 , _w_reg_N92 , _w_reg_N91 ,_w_reg_N90 , _w_reg_N89 , _w_reg_N88 , _w_reg_N87 , _w_reg_N86 ,_w_reg_N85 , _w_reg_N84 , _w_reg_N83 , _w_reg_N82 , _w_reg_N81 ,_w_reg_N80 , _w_reg_N79 , _w_reg_N78 , _w_reg_N77 , _w_reg_N76 ,_w_reg_N75 , _w_reg_N74 , _w_reg_N73 , _w_reg_N72 , _w_reg_N71 ,_w_reg_N70 , _w_reg_N69 , _w_reg_N68 , _w_reg_N67 , _w_reg_N66 ,_w_reg_N65 , _w_reg_N64 , _w_reg_N63 , _w_reg_N62 , _w_reg_N61 ,_w_reg_N60 , _w_reg_N59 , _w_reg_N58 , _w_reg_N57 , _w_reg_N56 ,_w_reg_N55 , _w_reg_N54 , _w_reg_N53 , _w_reg_N52 , _w_reg_N51 ,_w_reg_N50 , _w_reg_N49 , _w_reg_N48 , _w_reg_N47 , _w_reg_N46 ,_w_reg_N45 , _w_reg_N44 , _w_reg_N43 , _w_reg_N42 , _w_reg_N41 ,_w_reg_N40 , _w_reg_N39 , _w_reg_N38 , _w_reg_N37 , _w_reg_N36 ,_w_reg_N35 , _w_reg_N34 , _w_reg_N33 , _w_reg_N32 , _w_reg_N31 ,_w_reg_N30 , _w_reg_N29 , _w_reg_N28 , _w_reg_N27 , _w_reg_N26 ,_w_reg_N25 , _w_reg_N24 , _w_reg_N23 , _w_reg_N22 , _w_reg_N21 ,_w_reg_N20 , _w_reg_N19 , _w_reg_N18 , _w_reg_N17 , _w_reg_N16 ,_w_reg_N15 , _w_reg_N14 , _w_reg_N13 , _w_reg_N12 , _w_reg_N11 ,_w_reg_N10 , _w_reg_N9 , _w_reg_N8 , _w_reg_N7 , _w_reg_N6 ,_w_reg_N5 , _w_reg_N4 , _w_reg_N3 , _cv_reg_n330 , _cv_reg_n320 ,_cv_reg_n310 , _cv_reg_n300 , _cv_reg_n290 , _cv_reg_n280 ,_cv_reg_n270 , _cv_reg_n260 , _cv_reg_n250 , _cv_reg_n240 ,_cv_reg_n230 , _cv_reg_n220 , _cv_reg_n210 , _cv_reg_n200 ,_cv_reg_n190 , _cv_reg_n180 , _cv_reg_n170 , _cv_reg_N162 ,_cv_reg_N161 , _cv_reg_N160 , _cv_reg_N159 , _cv_reg_N158 ,_cv_reg_N157 , _cv_reg_N156 , _cv_reg_N155 , _cv_reg_N154 ,_cv_reg_N153 , _cv_reg_N152 , _cv_reg_N151 , _cv_reg_N150 ,_cv_reg_N149 , _cv_reg_N148 , _cv_reg_N147 , _cv_reg_N146 ,_cv_reg_N145 , _cv_reg_N144 , _cv_reg_N143 , _cv_reg_N142 ,_cv_reg_N141 , _cv_reg_N140 , _cv_reg_N139 , _cv_reg_N138 ,_cv_reg_N137 , _cv_reg_N136 , _cv_reg_N135 , _cv_reg_N134 ,_cv_reg_N133 , _cv_reg_N132 , _cv_reg_N131 , _cv_reg_N130 ,_cv_reg_N129 , _cv_reg_N128 , _cv_reg_N127 , _cv_reg_N126 ,_cv_reg_N125 , _cv_reg_N124 , _cv_reg_N123 , _cv_reg_N122 ,_cv_reg_N121 , _cv_reg_N120 , _cv_reg_N119 , _cv_reg_N118 ,_cv_reg_N117 , _cv_reg_N116 , _cv_reg_N115 , _cv_reg_N114 ,_cv_reg_N113 , _cv_reg_N112 , _cv_reg_N111 , _cv_reg_N110 ,_cv_reg_N109 , _cv_reg_N108 , _cv_reg_N107 , _cv_reg_N106 ,_cv_reg_N105 , _cv_reg_N104 , _cv_reg_N103 , _cv_reg_N102 ,_cv_reg_N101 , _cv_reg_N100 , _cv_reg_N99 , _cv_reg_N98 ,_cv_reg_N97 , _cv_reg_N96 , _cv_reg_N95 , _cv_reg_N94 , _cv_reg_N93 ,_cv_reg_N92 , _cv_reg_N91 , _cv_reg_N90 , _cv_reg_N89 , _cv_reg_N88 ,_cv_reg_N87 , _cv_reg_N86 , _cv_reg_N85 , _cv_reg_N84 , _cv_reg_N83 ,_cv_reg_N82 , _cv_reg_N81 , _cv_reg_N80 , _cv_reg_N79 , _cv_reg_N78 ,_cv_reg_N77 , _cv_reg_N76 , _cv_reg_N75 , _cv_reg_N74 , _cv_reg_N73 ,_cv_reg_N72 , _cv_reg_N71 , _cv_reg_N70 , _cv_reg_N69 , _cv_reg_N68 ,_cv_reg_N67 , _cv_reg_N66 , _cv_reg_N65 , _cv_reg_N64 , _cv_reg_N63 ,_cv_reg_N62 , _cv_reg_N61 , _cv_reg_N60 , _cv_reg_N59 , _cv_reg_N58 ,_cv_reg_N57 , _cv_reg_N56 , _cv_reg_N55 , _cv_reg_N54 , _cv_reg_N53 ,_cv_reg_N52 , _cv_reg_N51 , _cv_reg_N50 , _cv_reg_N49 , _cv_reg_N48 ,_cv_reg_N47 , _cv_reg_N46 , _cv_reg_N45 , _cv_reg_N44 , _cv_reg_N43 ,_cv_reg_N42 , _cv_reg_N41 , _cv_reg_N40 , _cv_reg_N39 , _cv_reg_N38 ,_cv_reg_N37 , _cv_reg_N36 , _cv_reg_N35 , _cv_reg_N34 , _cv_reg_N33 ,_cv_reg_N32 , _cv_reg_N31 , _cv_reg_N30 , _cv_reg_N29 , _cv_reg_N28 ,_cv_reg_N27 , _cv_reg_N26 , _cv_reg_N25 , _cv_reg_N24 , _cv_reg_N23 ,_cv_reg_N22 , _cv_reg_N21 , _cv_reg_N20 , _cv_reg_N19 , _cv_reg_N18 ,_cv_reg_N17 , _cv_reg_N16 , _cv_reg_N15 , _cv_reg_N14 , _cv_reg_N13 ,_cv_reg_N12 , _cv_reg_N11 , _cv_reg_N10 , _cv_reg_N9 , _cv_reg_N8 ,_cv_reg_N7 , _cv_reg_N6 , _cv_reg_N5 , _cv_reg_N4 , _cv_reg_N3 ,_rnd_reg_n320 , _rnd_reg_n310 , _rnd_reg_n300 , _rnd_reg_n290 ,_rnd_reg_n280 , _rnd_reg_n270 , _rnd_reg_n260 , _rnd_reg_n250 ,_rnd_reg_n240 , _rnd_reg_n230 , _rnd_reg_n220 , _rnd_reg_n210 ,_rnd_reg_n200 , _rnd_reg_n190 , _rnd_reg_n180 , _rnd_reg_n170 ,_rnd_reg_N162 , _rnd_reg_N161 , _rnd_reg_N160 , _rnd_reg_N159 ,_rnd_reg_N158 , _rnd_reg_N157 , _rnd_reg_N156 , _rnd_reg_N155 ,_rnd_reg_N154 , _rnd_reg_N153 , _rnd_reg_N152 , _rnd_reg_N151 ,_rnd_reg_N150 , _rnd_reg_N149 , _rnd_reg_N148 , _rnd_reg_N147 ,_rnd_reg_N146 , _rnd_reg_N145 , _rnd_reg_N144 , _rnd_reg_N143 ,_rnd_reg_N142 , _rnd_reg_N141 , _rnd_reg_N140 , _rnd_reg_N139 ,_rnd_reg_N138 , _rnd_reg_N137 , _rnd_reg_N136 , _rnd_reg_N135 ,_rnd_reg_N134 , _rnd_reg_N133 , _rnd_reg_N132 , _rnd_reg_N131 ,_rnd_reg_N130 , _rnd_reg_N129 , _rnd_reg_N128 , _rnd_reg_N127 ,_rnd_reg_N126 , _rnd_reg_N125 , _rnd_reg_N124 , _rnd_reg_N123 ,_rnd_reg_N122 , _rnd_reg_N121 , _rnd_reg_N120 , _rnd_reg_N119 ,_rnd_reg_N118 , _rnd_reg_N117 , _rnd_reg_N116 , _rnd_reg_N115 ,_rnd_reg_N114 , _rnd_reg_N113 , _rnd_reg_N112 , _rnd_reg_N111 ,_rnd_reg_N110 , _rnd_reg_N109 , _rnd_reg_N108 , _rnd_reg_N107 ,_rnd_reg_N106 , _rnd_reg_N105 , _rnd_reg_N104 , _rnd_reg_N103 ,_rnd_reg_N102 , _rnd_reg_N101 , _rnd_reg_N100 , _rnd_reg_N99 ,_rnd_reg_N98 , _rnd_reg_N97 , _rnd_reg_N96 , _rnd_reg_N95 ,_rnd_reg_N94 , _rnd_reg_N93 , _rnd_reg_N92 , _rnd_reg_N91 ,_rnd_reg_N90 , _rnd_reg_N89 , _rnd_reg_N88 , _rnd_reg_N87 ,_rnd_reg_N86 , _rnd_reg_N85 , _rnd_reg_N84 , _rnd_reg_N83 ,_rnd_reg_N82 , _rnd_reg_N81 , _rnd_reg_N80 , _rnd_reg_N79 ,_rnd_reg_N78 , _rnd_reg_N77 , _rnd_reg_N76 , _rnd_reg_N75 ,_rnd_reg_N74 , _rnd_reg_N73 , _rnd_reg_N72 , _rnd_reg_N71 ,_rnd_reg_N70 , _rnd_reg_N69 , _rnd_reg_N68 , _rnd_reg_N67 ,_rnd_reg_N66 , _rnd_reg_N65 , _rnd_reg_N64 , _rnd_reg_N63 ,_rnd_reg_N62 , _rnd_reg_N61 , _rnd_reg_N60 , _rnd_reg_N59 ,_rnd_reg_N58 , _rnd_reg_N57 , _rnd_reg_N56 , _rnd_reg_N55 ,_rnd_reg_N54 , _rnd_reg_N53 , _rnd_reg_N52 , _rnd_reg_N51 ,_rnd_reg_N50 , _rnd_reg_N49 , _rnd_reg_N48 , _rnd_reg_N47 ,_rnd_reg_N46 , _rnd_reg_N45 , _rnd_reg_N44 , _rnd_reg_N43 ,_rnd_reg_N42 , _rnd_reg_N41 , _rnd_reg_N40 , _rnd_reg_N39 ,_rnd_reg_N38 , _rnd_reg_N37 , _rnd_reg_N36 , _rnd_reg_N35 ,_rnd_reg_N34 , _rnd_reg_N33 , _rnd_reg_N32 , _rnd_reg_N31 ,_rnd_reg_N30 , _rnd_reg_N29 , _rnd_reg_N28 , _rnd_reg_N27 ,_rnd_reg_N26 , _rnd_reg_N25 , _rnd_reg_N24 , _rnd_reg_N23 ,_rnd_reg_N22 , _rnd_reg_N21 , _rnd_reg_N20 , _rnd_reg_N19 ,_rnd_reg_N18 , _rnd_reg_N17 , _rnd_reg_N16 , _rnd_reg_N15 ,_rnd_reg_N14 , _rnd_reg_N13 , _rnd_reg_N12 , _rnd_reg_N11 ,_rnd_reg_N10 , _rnd_reg_N9 , _rnd_reg_N8 , _rnd_reg_N7 , _rnd_reg_N6 ,_rnd_reg_N5 , _rnd_reg_N4 , _rnd_reg_N3 , _cv_next_reg_n320 ,_cv_next_reg_n310 , _cv_next_reg_n300 , _cv_next_reg_n290 ,_cv_next_reg_n280 , _cv_next_reg_n270 , _cv_next_reg_n260 ,_cv_next_reg_n250 , _cv_next_reg_n240 , _cv_next_reg_n230 ,_cv_next_reg_n220 , _cv_next_reg_n210 , _cv_next_reg_n200 ,_cv_next_reg_n190 , _cv_next_reg_n180 , _cv_next_reg_n170 ,_cv_next_reg_N162 , _cv_next_reg_N161 , _cv_next_reg_N160 ,_cv_next_reg_N159 , _cv_next_reg_N158 , _cv_next_reg_N157 ,_cv_next_reg_N156 , _cv_next_reg_N155 , _cv_next_reg_N154 ,_cv_next_reg_N153 , _cv_next_reg_N152 , _cv_next_reg_N151 ,_cv_next_reg_N150 , _cv_next_reg_N149 , _cv_next_reg_N148 ,_cv_next_reg_N147 , _cv_next_reg_N146 , _cv_next_reg_N145 ,_cv_next_reg_N144 , _cv_next_reg_N143 , _cv_next_reg_N142 ,_cv_next_reg_N141 , _cv_next_reg_N140 , _cv_next_reg_N139 ,_cv_next_reg_N138 , _cv_next_reg_N137 , _cv_next_reg_N136 ,_cv_next_reg_N135 , _cv_next_reg_N134 , _cv_next_reg_N133 ,_cv_next_reg_N132 , _cv_next_reg_N131 , _cv_next_reg_N130 ,_cv_next_reg_N129 , _cv_next_reg_N128 , _cv_next_reg_N127 ,_cv_next_reg_N126 , _cv_next_reg_N125 , _cv_next_reg_N124 ,_cv_next_reg_N123 , _cv_next_reg_N122 , _cv_next_reg_N121 ,_cv_next_reg_N120 , _cv_next_reg_N119 , _cv_next_reg_N118 ,_cv_next_reg_N117 , _cv_next_reg_N116 , _cv_next_reg_N115 ,_cv_next_reg_N114 , _cv_next_reg_N113 , _cv_next_reg_N112 ,_cv_next_reg_N111 , _cv_next_reg_N110 , _cv_next_reg_N109 ,_cv_next_reg_N108 , _cv_next_reg_N107 , _cv_next_reg_N106 ,_cv_next_reg_N105 , _cv_next_reg_N104 , _cv_next_reg_N103 ,_cv_next_reg_N102 , _cv_next_reg_N101 , _cv_next_reg_N100 ,_cv_next_reg_N99 , _cv_next_reg_N98 , _cv_next_reg_N97 ,_cv_next_reg_N96 , _cv_next_reg_N95 , _cv_next_reg_N94 ,_cv_next_reg_N93 , _cv_next_reg_N92 , _cv_next_reg_N91 ,_cv_next_reg_N90 , _cv_next_reg_N89 , _cv_next_reg_N88 ,_cv_next_reg_N87 , _cv_next_reg_N86 , _cv_next_reg_N85 ,_cv_next_reg_N84 , _cv_next_reg_N83 , _cv_next_reg_N82 ,_cv_next_reg_N81 , _cv_next_reg_N80 , _cv_next_reg_N79 ,_cv_next_reg_N78 , _cv_next_reg_N77 , _cv_next_reg_N76 ,_cv_next_reg_N75 , _cv_next_reg_N74 , _cv_next_reg_N73 ,_cv_next_reg_N72 , _cv_next_reg_N71 , _cv_next_reg_N70 ,_cv_next_reg_N69 , _cv_next_reg_N68 , _cv_next_reg_N67 ,_cv_next_reg_N66 , _cv_next_reg_N65 , _cv_next_reg_N64 ,_cv_next_reg_N63 , _cv_next_reg_N62 , _cv_next_reg_N61 ,_cv_next_reg_N60 , _cv_next_reg_N59 , _cv_next_reg_N58 ,_cv_next_reg_N57 , _cv_next_reg_N56 , _cv_next_reg_N55 ,_cv_next_reg_N54 , _cv_next_reg_N53 , _cv_next_reg_N52 ,_cv_next_reg_N51 , _cv_next_reg_N50 , _cv_next_reg_N49 ,_cv_next_reg_N48 , _cv_next_reg_N47 , _cv_next_reg_N46 ,_cv_next_reg_N45 , _cv_next_reg_N44 , _cv_next_reg_N43 ,_cv_next_reg_N42 , _cv_next_reg_N41 , _cv_next_reg_N40 ,_cv_next_reg_N39 , _cv_next_reg_N38 , _cv_next_reg_N37 ,_cv_next_reg_N36 , _cv_next_reg_N35 , _cv_next_reg_N34 ,_cv_next_reg_N33 , _cv_next_reg_N32 , _cv_next_reg_N31 ,_cv_next_reg_N30 , _cv_next_reg_N29 , _cv_next_reg_N28 ,_cv_next_reg_N27 , _cv_next_reg_N26 , _cv_next_reg_N25 ,_cv_next_reg_N24 , _cv_next_reg_N23 , _cv_next_reg_N22 ,_cv_next_reg_N21 , _cv_next_reg_N20 , _cv_next_reg_N19 ,_cv_next_reg_N18 , _cv_next_reg_N17 , _cv_next_reg_N16 ,_cv_next_reg_N15 , _cv_next_reg_N14 , _cv_next_reg_N13 ,_cv_next_reg_N12 , _cv_next_reg_N11 , _cv_next_reg_N10 ,_cv_next_reg_N9 , _cv_next_reg_N8 , _cv_next_reg_N7 ,_cv_next_reg_N6 , _cv_next_reg_N5 , _cv_next_reg_N4 ,_cv_next_reg_N3 , _add_98_2_n379 , _add_98_2_n378 , _add_98_2_n377 ,_add_98_2_n376 , _add_98_2_n375 , _add_98_2_n374 , _add_98_2_n373 ,_add_98_2_n372 , _add_98_2_n371 , _add_98_2_n370 , _add_98_2_n369 ,_add_98_2_n368 , _add_98_2_n367 , _add_98_2_n366 , _add_98_2_n365 ,_add_98_2_n364 , _add_98_2_n363 , _add_98_2_n362 , _add_98_2_n361 ,_add_98_2_n360 , _add_98_2_n359 , _add_98_2_n358 , _add_98_2_n357 ,_add_98_2_n356 , _add_98_2_n355 , _add_98_2_n354 , _add_98_2_n353 ,_add_98_2_n352 , _add_98_2_n351 , _add_98_2_n350 , _add_98_2_n349 ,_add_98_2_n348 , _add_98_2_n347 , _add_98_2_n346 , _add_98_2_n345 ,_add_98_2_n344 , _add_98_2_n343 , _add_98_2_n342 , _add_98_2_n341 ,_add_98_2_n340 , _add_98_2_n339 , _add_98_2_n338 , _add_98_2_n337 ,_add_98_2_n336 , _add_98_2_n335 , _add_98_2_n334 , _add_98_2_n333 ,_add_98_2_n332 , _add_98_2_n331 , _add_98_2_n330 , _add_98_2_n329 ,_add_98_2_n328 , _add_98_2_n327 , _add_98_2_n326 , _add_98_2_n325 ,_add_98_2_n324 , _add_98_2_n323 , _add_98_2_n322 , _add_98_2_n321 ,_add_98_2_n320 , _add_98_2_n319 , _add_98_2_n318 , _add_98_2_n317 ,_add_98_2_n316 , _add_98_2_n315 , _add_98_2_n314 , _add_98_2_n313 ,_add_98_2_n312 , _add_98_2_n311 , _add_98_2_n310 , _add_98_2_n309 ,_add_98_2_n308 , _add_98_2_n307 , _add_98_2_n306 , _add_98_2_n305 ,_add_98_2_n304 , _add_98_2_n303 , _add_98_2_n302 , _add_98_2_n301 ,_add_98_2_n300 , _add_98_2_n299 , _add_98_2_n298 , _add_98_2_n297 ,_add_98_2_n296 , _add_98_2_n295 , _add_98_2_n294 , _add_98_2_n293 ,_add_98_2_n292 , _add_98_2_n291 , _add_98_2_n290 , _add_98_2_n289 ,_add_98_2_n288 , _add_98_2_n287 , _add_98_2_n286 , _add_98_2_n285 ,_add_98_2_n284 , _add_98_2_n283 , _add_98_2_n282 , _add_98_2_n281 ,_add_98_2_n280 , _add_98_2_n279 , _add_98_2_n278 , _add_98_2_n277 ,_add_98_2_n276 , _add_98_2_n275 , _add_98_2_n274 , _add_98_2_n273 ,_add_98_2_n272 , _add_98_2_n271 , _add_98_2_n270 , _add_98_2_n269 ,_add_98_2_n268 , _add_98_2_n267 , _add_98_2_n266 , _add_98_2_n265 ,_add_98_2_n264 , _add_98_2_n263 , _add_98_2_n262 , _add_98_2_n261 ,_add_98_2_n260 , _add_98_2_n259 , _add_98_2_n258 , _add_98_2_n257 ,_add_98_2_n256 , _add_98_2_n255 , _add_98_2_n254 , _add_98_2_n253 ,_add_98_2_n252 , _add_98_2_n251 , _add_98_2_n250 , _add_98_2_n249 ,_add_98_2_n248 , _add_98_2_n247 , _add_98_2_n246 , _add_98_2_n245 ,_add_98_2_n244 , _add_98_2_n243 , _add_98_2_n242 , _add_98_2_n241 ,_add_98_2_n240 , _add_98_2_n239 , _add_98_2_n238 , _add_98_2_n237 ,_add_98_2_n236 , _add_98_2_n235 , _add_98_2_n234 , _add_98_2_n233 ,_add_98_2_n232 , _add_98_2_n231 , _add_98_2_n230 , _add_98_2_n229 ,_add_98_2_n228 , _add_98_2_n227 , _add_98_2_n226 , _add_98_2_n225 ,_add_98_2_n224 , _add_98_2_n223 , _add_98_2_n222 , _add_98_2_n221 ,_add_98_2_n220 , _add_98_2_n219 , _add_98_2_n218 , _add_98_2_n217 ,_add_98_2_n216 , _add_98_2_n215 , _add_98_2_n214 , _add_98_2_n213 ,_add_98_2_n212 , _add_98_2_n211 , _add_98_2_n210 , _add_98_2_n209 ,_add_98_2_n208 , _add_98_2_n207 , _add_98_2_n206 , _add_98_2_n205 ,_add_98_2_n204 , _add_98_2_n203 , _add_98_2_n202 , _add_98_2_n201 ,_add_98_2_n200 , _add_98_2_n199 , _add_98_2_n198 , _add_98_2_n197 ,_add_98_2_n196 , _add_98_2_n195 , _add_98_2_n194 , _add_98_2_n193 ,_add_98_2_n192 , _add_98_2_n191 , _add_98_2_n190 , _add_98_2_n189 ,_add_98_2_n188 , _add_98_2_n187 , _add_98_2_n186 , _add_98_2_n185 ,_add_98_2_n184 , _add_98_2_n183 , _add_98_2_n182 , _add_98_2_n181 ,_add_98_2_n180 , _add_98_2_n179 , _add_98_2_n178 , _add_98_2_n177 ,_add_98_2_n176 , _add_98_2_n175 , _add_98_2_n174 , _add_98_2_n173 ,_add_98_2_n172 , _add_98_2_n171 , _add_98_2_n170 , _add_98_2_n169 ,_add_98_2_n168 , _add_98_2_n167 , _add_98_2_n166 , _add_98_2_n165 ,_add_98_2_n164 , _add_98_2_n163 , _add_98_2_n162 , _add_98_2_n161 ,_add_98_2_n160 , _add_98_2_n159 , _add_98_2_n158 , _add_98_2_n157 ,_add_98_2_n156 , _add_98_2_n155 , _add_98_2_n154 , _add_98_2_n153 ,_add_98_2_n152 , _add_98_2_n151 , _add_98_2_n150 , _add_98_2_n149 ,_add_98_2_n148 , _add_98_2_n147 , _add_98_2_n146 , _add_98_2_n145 ,_add_98_2_n144 , _add_98_2_n143 , _add_98_2_n142 , _add_98_2_n141 ,_add_98_2_n140 , _add_98_2_n139 , _add_98_2_n138 , _add_98_2_n137 ,_add_98_2_n136 , _add_98_2_n135 , _add_98_2_n134 , _add_98_2_n133 ,_add_98_2_n132 , _add_98_2_n131 , _add_98_2_n130 , _add_98_2_n129 ,_add_98_2_n128 , _add_98_2_n127 , _add_98_2_n126 , _add_98_2_n125 ,_add_98_2_n124 , _add_98_2_n123 , _add_98_2_n122 , _add_98_2_n121 ,_add_98_2_n120 , _add_98_2_n119 , _add_98_2_n118 , _add_98_2_n117 ,_add_98_2_n116 , _add_98_2_n115 , _add_98_2_n114 , _add_98_2_n113 ,_add_98_2_n112 , _add_98_2_n111 , _add_98_2_n110 , _add_98_2_n109 ,_add_98_2_n108 , _add_98_2_n107 , _add_98_2_n106 , _add_98_2_n105 ,_add_98_2_n104 , _add_98_2_n103 , _add_98_2_n102 , _add_98_2_n101 ,_add_98_2_n100 , _add_98_2_n99 , _add_98_2_n98 , _add_98_2_n97 ,_add_98_2_n96 , _add_98_2_n95 , _add_98_2_n94 , _add_98_2_n93 ,_add_98_2_n92 , _add_98_2_n91 , _add_98_2_n90 , _add_98_2_n89 ,_add_98_2_n88 , _add_98_2_n87 , _add_98_2_n86 , _add_98_2_n85 ,_add_98_2_n84 , _add_98_2_n83 , _add_98_2_n82 , _add_98_2_n81 ,_add_98_2_n80 , _add_98_2_n79 , _add_98_2_n78 , _add_98_2_n77 ,_add_98_2_n76 , _add_98_2_n75 , _add_98_2_n74 , _add_98_2_n73 ,_add_98_2_n72 , _add_98_2_n71 , _add_98_2_n70 , _add_98_2_n69 ,_add_98_2_n68 , _add_98_2_n67 , _add_98_2_n66 , _add_98_2_n65 ,_add_98_2_n64 , _add_98_2_n63 , _add_98_2_n62 , _add_98_2_n61 ,_add_98_2_n60 , _add_98_2_n59 , _add_98_2_n58 , _add_98_2_n57 ,_add_98_2_n56 , _add_98_2_n55 , _add_98_2_n54 , _add_98_2_n53 ,_add_98_2_n52 , _add_98_2_n51 , _add_98_2_n50 , _add_98_2_n49 ,_add_98_2_n48 , _add_98_2_n47 , _add_98_2_n46 , _add_98_2_n45 ,_add_98_2_n44 , _add_98_2_n43 , _add_98_2_n42 , _add_98_2_n41 ,_add_98_2_n40 , _add_98_2_n39 , _add_98_2_n38 , _add_98_2_n37 ,_add_98_2_n36 , _add_98_2_n35 , _add_98_2_n34 , _add_98_2_n33 ,_add_98_2_n32 , _add_98_2_n31 , _add_98_2_n30 , _add_98_2_n29 ,_add_98_2_n28 , _add_98_2_n26 , _add_98_2_n25 , _add_98_2_n24 ,_add_98_2_n23 , _add_98_2_n22 , _add_98_2_n21 , _add_98_2_n20 ,_add_98_2_n19 , _add_98_2_n18 , _add_98_2_n17 , _add_98_2_n16 ,_add_98_2_n15 , _add_98_2_n14 , _add_98_2_n13 , _add_98_2_n12 ,_add_98_2_n11 , _add_98_2_n10 , _add_98_2_n9 , _add_98_2_n8 ,_add_98_2_n7 , _add_98_2_n6 , _add_98_2_n5 , _add_98_2_n4 ,_add_98_2_n3 , _add_98_2_n2 , _add_98_2_n1 , _add_98_3_n381 ,_add_98_3_n380 , _add_98_3_n379 , _add_98_3_n378 , _add_98_3_n377 ,_add_98_3_n376 , _add_98_3_n375 , _add_98_3_n374 , _add_98_3_n373 ,_add_98_3_n372 , _add_98_3_n371 , _add_98_3_n370 , _add_98_3_n369 ,_add_98_3_n368 , _add_98_3_n367 , _add_98_3_n366 , _add_98_3_n365 ,_add_98_3_n364 , _add_98_3_n363 , _add_98_3_n362 , _add_98_3_n361 ,_add_98_3_n360 , _add_98_3_n359 , _add_98_3_n358 , _add_98_3_n357 ,_add_98_3_n356 , _add_98_3_n355 , _add_98_3_n354 , _add_98_3_n353 ,_add_98_3_n352 , _add_98_3_n351 , _add_98_3_n350 , _add_98_3_n349 ,_add_98_3_n348 , _add_98_3_n347 , _add_98_3_n346 , _add_98_3_n345 ,_add_98_3_n344 , _add_98_3_n343 , _add_98_3_n342 , _add_98_3_n341 ,_add_98_3_n340 , _add_98_3_n339 , _add_98_3_n338 , _add_98_3_n337 ,_add_98_3_n336 , _add_98_3_n335 , _add_98_3_n334 , _add_98_3_n333 ,_add_98_3_n332 , _add_98_3_n331 , _add_98_3_n330 , _add_98_3_n329 ,_add_98_3_n328 , _add_98_3_n327 , _add_98_3_n326 , _add_98_3_n325 ,_add_98_3_n324 , _add_98_3_n323 , _add_98_3_n322 , _add_98_3_n321 ,_add_98_3_n320 , _add_98_3_n319 , _add_98_3_n318 , _add_98_3_n317 ,_add_98_3_n316 , _add_98_3_n315 , _add_98_3_n314 , _add_98_3_n313 ,_add_98_3_n312 , _add_98_3_n311 , _add_98_3_n310 , _add_98_3_n309 ,_add_98_3_n308 , _add_98_3_n307 , _add_98_3_n306 , _add_98_3_n305 ,_add_98_3_n304 , _add_98_3_n303 , _add_98_3_n302 , _add_98_3_n301 ,_add_98_3_n300 , _add_98_3_n299 , _add_98_3_n298 , _add_98_3_n297 ,_add_98_3_n296 , _add_98_3_n295 , _add_98_3_n294 , _add_98_3_n293 ,_add_98_3_n292 , _add_98_3_n291 , _add_98_3_n290 , _add_98_3_n289 ,_add_98_3_n288 , _add_98_3_n287 , _add_98_3_n286 , _add_98_3_n285 ,_add_98_3_n284 , _add_98_3_n283 , _add_98_3_n282 , _add_98_3_n281 ,_add_98_3_n280 , _add_98_3_n279 , _add_98_3_n278 , _add_98_3_n277 ,_add_98_3_n276 , _add_98_3_n275 , _add_98_3_n274 , _add_98_3_n273 ,_add_98_3_n272 , _add_98_3_n271 , _add_98_3_n270 , _add_98_3_n269 ,_add_98_3_n268 , _add_98_3_n267 , _add_98_3_n266 , _add_98_3_n265 ,_add_98_3_n264 , _add_98_3_n263 , _add_98_3_n262 , _add_98_3_n261 ,_add_98_3_n260 , _add_98_3_n259 , _add_98_3_n258 , _add_98_3_n257 ,_add_98_3_n256 , _add_98_3_n255 , _add_98_3_n254 , _add_98_3_n253 ,_add_98_3_n252 , _add_98_3_n251 , _add_98_3_n250 , _add_98_3_n249 ,_add_98_3_n248 , _add_98_3_n247 , _add_98_3_n246 , _add_98_3_n245 ,_add_98_3_n244 , _add_98_3_n243 , _add_98_3_n242 , _add_98_3_n241 ,_add_98_3_n240 , _add_98_3_n239 , _add_98_3_n238 , _add_98_3_n237 ,_add_98_3_n236 , _add_98_3_n235 , _add_98_3_n234 , _add_98_3_n233 ,_add_98_3_n232 , _add_98_3_n231 , _add_98_3_n230 , _add_98_3_n229 ,_add_98_3_n228 , _add_98_3_n227 , _add_98_3_n226 , _add_98_3_n225 ,_add_98_3_n224 , _add_98_3_n223 , _add_98_3_n222 , _add_98_3_n221 ,_add_98_3_n220 , _add_98_3_n219 , _add_98_3_n218 , _add_98_3_n217 ,_add_98_3_n216 , _add_98_3_n215 , _add_98_3_n214 , _add_98_3_n213 ,_add_98_3_n212 , _add_98_3_n211 , _add_98_3_n210 , _add_98_3_n209 ,_add_98_3_n208 , _add_98_3_n207 , _add_98_3_n206 , _add_98_3_n205 ,_add_98_3_n204 , _add_98_3_n203 , _add_98_3_n202 , _add_98_3_n201 ,_add_98_3_n200 , _add_98_3_n199 , _add_98_3_n198 , _add_98_3_n197 ,_add_98_3_n196 , _add_98_3_n195 , _add_98_3_n194 , _add_98_3_n193 ,_add_98_3_n192 , _add_98_3_n191 , _add_98_3_n190 , _add_98_3_n189 ,_add_98_3_n188 , _add_98_3_n187 , _add_98_3_n186 , _add_98_3_n185 ,_add_98_3_n184 , _add_98_3_n183 , _add_98_3_n182 , _add_98_3_n181 ,_add_98_3_n180 , _add_98_3_n179 , _add_98_3_n178 , _add_98_3_n177 ,_add_98_3_n176 , _add_98_3_n175 , _add_98_3_n174 , _add_98_3_n173 ,_add_98_3_n172 , _add_98_3_n171 , _add_98_3_n170 , _add_98_3_n169 ,_add_98_3_n168 , _add_98_3_n167 , _add_98_3_n166 , _add_98_3_n165 ,_add_98_3_n164 , _add_98_3_n163 , _add_98_3_n162 , _add_98_3_n161 ,_add_98_3_n160 , _add_98_3_n159 , _add_98_3_n158 , _add_98_3_n157 ,_add_98_3_n156 , _add_98_3_n155 , _add_98_3_n154 , _add_98_3_n153 ,_add_98_3_n152 , _add_98_3_n151 , _add_98_3_n150 , _add_98_3_n149 ,_add_98_3_n148 , _add_98_3_n147 , _add_98_3_n146 , _add_98_3_n145 ,_add_98_3_n144 , _add_98_3_n143 , _add_98_3_n142 , _add_98_3_n141 ,_add_98_3_n140 , _add_98_3_n139 , _add_98_3_n138 , _add_98_3_n137 ,_add_98_3_n136 , _add_98_3_n135 , _add_98_3_n134 , _add_98_3_n133 ,_add_98_3_n132 , _add_98_3_n131 , _add_98_3_n130 , _add_98_3_n129 ,_add_98_3_n128 , _add_98_3_n127 , _add_98_3_n126 , _add_98_3_n125 ,_add_98_3_n124 , _add_98_3_n123 , _add_98_3_n122 , _add_98_3_n121 ,_add_98_3_n120 , _add_98_3_n119 , _add_98_3_n118 , _add_98_3_n117 ,_add_98_3_n116 , _add_98_3_n115 , _add_98_3_n114 , _add_98_3_n113 ,_add_98_3_n112 , _add_98_3_n111 , _add_98_3_n110 , _add_98_3_n109 ,_add_98_3_n108 , _add_98_3_n107 , _add_98_3_n106 , _add_98_3_n105 ,_add_98_3_n104 , _add_98_3_n103 , _add_98_3_n102 , _add_98_3_n101 ,_add_98_3_n100 , _add_98_3_n99 , _add_98_3_n98 , _add_98_3_n97 ,_add_98_3_n96 , _add_98_3_n95 , _add_98_3_n94 , _add_98_3_n93 ,_add_98_3_n92 , _add_98_3_n91 , _add_98_3_n90 , _add_98_3_n89 ,_add_98_3_n88 , _add_98_3_n87 , _add_98_3_n86 , _add_98_3_n85 ,_add_98_3_n84 , _add_98_3_n83 , _add_98_3_n82 , _add_98_3_n81 ,_add_98_3_n80 , _add_98_3_n79 , _add_98_3_n78 , _add_98_3_n77 ,_add_98_3_n76 , _add_98_3_n75 , _add_98_3_n74 , _add_98_3_n73 ,_add_98_3_n72 , _add_98_3_n71 , _add_98_3_n70 , _add_98_3_n69 ,_add_98_3_n68 , _add_98_3_n67 , _add_98_3_n66 , _add_98_3_n65 ,_add_98_3_n64 , _add_98_3_n63 , _add_98_3_n62 , _add_98_3_n61 ,_add_98_3_n60 , _add_98_3_n59 , _add_98_3_n58 , _add_98_3_n57 ,_add_98_3_n56 , _add_98_3_n55 , _add_98_3_n54 , _add_98_3_n53 ,_add_98_3_n52 , _add_98_3_n51 , _add_98_3_n50 , _add_98_3_n49 ,_add_98_3_n48 , _add_98_3_n47 , _add_98_3_n46 , _add_98_3_n45 ,_add_98_3_n44 , _add_98_3_n43 , _add_98_3_n42 , _add_98_3_n41 ,_add_98_3_n40 , _add_98_3_n39 , _add_98_3_n38 , _add_98_3_n37 ,_add_98_3_n36 , _add_98_3_n35 , _add_98_3_n34 , _add_98_3_n33 ,_add_98_3_n32 , _add_98_3_n31 , _add_98_3_n30 , _add_98_3_n29 ,_add_98_3_n28 , _add_98_3_n26 , _add_98_3_n25 , _add_98_3_n24 ,_add_98_3_n23 , _add_98_3_n22 , _add_98_3_n21 , _add_98_3_n20 ,_add_98_3_n19 , _add_98_3_n18 , _add_98_3_n17 , _add_98_3_n16 ,_add_98_3_n15 , _add_98_3_n14 , _add_98_3_n13 , _add_98_3_n12 ,_add_98_3_n11 , _add_98_3_n10 , _add_98_3_n9 , _add_98_3_n8 ,_add_98_3_n7 , _add_98_3_n6 , _add_98_3_n5 , _add_98_3_n4 ,_add_98_3_n3 , _add_98_3_n2 , _add_98_3_n1 , _add_98_5_n392 ,_add_98_5_n391 , _add_98_5_n390 , _add_98_5_n389 , _add_98_5_n388 ,_add_98_5_n387 , _add_98_5_n386 , _add_98_5_n385 , _add_98_5_n384 ,_add_98_5_n383 , _add_98_5_n382 , _add_98_5_n381 , _add_98_5_n380 ,_add_98_5_n379 , _add_98_5_n378 , _add_98_5_n377 , _add_98_5_n376 ,_add_98_5_n375 , _add_98_5_n374 , _add_98_5_n373 , _add_98_5_n372 ,_add_98_5_n371 , _add_98_5_n370 , _add_98_5_n369 , _add_98_5_n368 ,_add_98_5_n367 , _add_98_5_n366 , _add_98_5_n365 , _add_98_5_n364 ,_add_98_5_n363 , _add_98_5_n362 , _add_98_5_n361 , _add_98_5_n360 ,_add_98_5_n359 , _add_98_5_n358 , _add_98_5_n357 , _add_98_5_n356 ,_add_98_5_n355 , _add_98_5_n354 , _add_98_5_n353 , _add_98_5_n352 ,_add_98_5_n351 , _add_98_5_n350 , _add_98_5_n349 , _add_98_5_n348 ,_add_98_5_n347 , _add_98_5_n346 , _add_98_5_n345 , _add_98_5_n344 ,_add_98_5_n343 , _add_98_5_n342 , _add_98_5_n341 , _add_98_5_n340 ,_add_98_5_n339 , _add_98_5_n338 , _add_98_5_n337 , _add_98_5_n336 ,_add_98_5_n335 , _add_98_5_n334 , _add_98_5_n333 , _add_98_5_n332 ,_add_98_5_n331 , _add_98_5_n330 , _add_98_5_n329 , _add_98_5_n328 ,_add_98_5_n327 , _add_98_5_n326 , _add_98_5_n325 , _add_98_5_n324 ,_add_98_5_n323 , _add_98_5_n322 , _add_98_5_n321 , _add_98_5_n320 ,_add_98_5_n319 , _add_98_5_n318 , _add_98_5_n317 , _add_98_5_n316 ,_add_98_5_n315 , _add_98_5_n314 , _add_98_5_n313 , _add_98_5_n312 ,_add_98_5_n311 , _add_98_5_n310 , _add_98_5_n309 , _add_98_5_n308 ,_add_98_5_n307 , _add_98_5_n306 , _add_98_5_n305 , _add_98_5_n304 ,_add_98_5_n303 , _add_98_5_n302 , _add_98_5_n301 , _add_98_5_n300 ,_add_98_5_n299 , _add_98_5_n298 , _add_98_5_n297 , _add_98_5_n296 ,_add_98_5_n295 , _add_98_5_n294 , _add_98_5_n293 , _add_98_5_n292 ,_add_98_5_n291 , _add_98_5_n290 , _add_98_5_n289 , _add_98_5_n288 ,_add_98_5_n287 , _add_98_5_n286 , _add_98_5_n285 , _add_98_5_n284 ,_add_98_5_n283 , _add_98_5_n282 , _add_98_5_n281 , _add_98_5_n280 ,_add_98_5_n279 , _add_98_5_n278 , _add_98_5_n277 , _add_98_5_n276 ,_add_98_5_n275 , _add_98_5_n274 , _add_98_5_n273 , _add_98_5_n272 ,_add_98_5_n271 , _add_98_5_n270 , _add_98_5_n269 , _add_98_5_n268 ,_add_98_5_n267 , _add_98_5_n266 , _add_98_5_n265 , _add_98_5_n264 ,_add_98_5_n263 , _add_98_5_n262 , _add_98_5_n261 , _add_98_5_n260 ,_add_98_5_n259 , _add_98_5_n258 , _add_98_5_n257 , _add_98_5_n256 ,_add_98_5_n255 , _add_98_5_n254 , _add_98_5_n253 , _add_98_5_n252 ,_add_98_5_n251 , _add_98_5_n250 , _add_98_5_n249 , _add_98_5_n248 ,_add_98_5_n247 , _add_98_5_n246 , _add_98_5_n245 , _add_98_5_n244 ,_add_98_5_n243 , _add_98_5_n242 , _add_98_5_n241 , _add_98_5_n240 ,_add_98_5_n239 , _add_98_5_n238 , _add_98_5_n237 , _add_98_5_n236 ,_add_98_5_n235 , _add_98_5_n234 , _add_98_5_n233 , _add_98_5_n232 ,_add_98_5_n231 , _add_98_5_n230 , _add_98_5_n229 , _add_98_5_n228 ,_add_98_5_n227 , _add_98_5_n226 , _add_98_5_n225 , _add_98_5_n224 ,_add_98_5_n223 , _add_98_5_n222 , _add_98_5_n221 , _add_98_5_n220 ,_add_98_5_n219 , _add_98_5_n218 , _add_98_5_n217 , _add_98_5_n216 ,_add_98_5_n215 , _add_98_5_n214 , _add_98_5_n213 , _add_98_5_n212 ,_add_98_5_n211 , _add_98_5_n210 , _add_98_5_n209 , _add_98_5_n208 ,_add_98_5_n207 , _add_98_5_n206 , _add_98_5_n205 , _add_98_5_n204 ,_add_98_5_n203 , _add_98_5_n202 , _add_98_5_n201 , _add_98_5_n200 ,_add_98_5_n199 , _add_98_5_n198 , _add_98_5_n197 , _add_98_5_n196 ,_add_98_5_n195 , _add_98_5_n194 , _add_98_5_n193 , _add_98_5_n192 ,_add_98_5_n191 , _add_98_5_n190 , _add_98_5_n189 , _add_98_5_n188 ,_add_98_5_n187 , _add_98_5_n186 , _add_98_5_n185 , _add_98_5_n184 ,_add_98_5_n183 , _add_98_5_n182 , _add_98_5_n181 , _add_98_5_n180 ,_add_98_5_n179 , _add_98_5_n178 , _add_98_5_n177 , _add_98_5_n176 ,_add_98_5_n175 , _add_98_5_n174 , _add_98_5_n173 , _add_98_5_n172 ,_add_98_5_n171 , _add_98_5_n170 , _add_98_5_n169 , _add_98_5_n168 ,_add_98_5_n167 , _add_98_5_n166 , _add_98_5_n165 , _add_98_5_n164 ,_add_98_5_n163 , _add_98_5_n162 , _add_98_5_n161 , _add_98_5_n160 ,_add_98_5_n159 , _add_98_5_n158 , _add_98_5_n157 , _add_98_5_n156 ,_add_98_5_n155 , _add_98_5_n154 , _add_98_5_n153 , _add_98_5_n152 ,_add_98_5_n151 , _add_98_5_n150 , _add_98_5_n149 , _add_98_5_n148 ,_add_98_5_n147 , _add_98_5_n146 , _add_98_5_n145 , _add_98_5_n144 ,_add_98_5_n143 , _add_98_5_n142 , _add_98_5_n141 , _add_98_5_n140 ,_add_98_5_n139 , _add_98_5_n138 , _add_98_5_n137 , _add_98_5_n136 ,_add_98_5_n135 , _add_98_5_n134 , _add_98_5_n133 , _add_98_5_n132 ,_add_98_5_n131 , _add_98_5_n130 , _add_98_5_n129 , _add_98_5_n128 ,_add_98_5_n127 , _add_98_5_n126 , _add_98_5_n125 , _add_98_5_n124 ,_add_98_5_n123 , _add_98_5_n122 , _add_98_5_n121 , _add_98_5_n120 ,_add_98_5_n119 , _add_98_5_n118 , _add_98_5_n117 , _add_98_5_n116 ,_add_98_5_n115 , _add_98_5_n114 , _add_98_5_n113 , _add_98_5_n112 ,_add_98_5_n111 , _add_98_5_n110 , _add_98_5_n109 , _add_98_5_n108 ,_add_98_5_n107 , _add_98_5_n106 , _add_98_5_n105 , _add_98_5_n104 ,_add_98_5_n103 , _add_98_5_n102 , _add_98_5_n101 , _add_98_5_n100 ,_add_98_5_n99 , _add_98_5_n98 , _add_98_5_n97 , _add_98_5_n96 ,_add_98_5_n95 , _add_98_5_n94 , _add_98_5_n93 , _add_98_5_n92 ,_add_98_5_n91 , _add_98_5_n90 , _add_98_5_n89 , _add_98_5_n88 ,_add_98_5_n87 , _add_98_5_n86 , _add_98_5_n85 , _add_98_5_n84 ,_add_98_5_n83 , _add_98_5_n82 , _add_98_5_n81 , _add_98_5_n80 ,_add_98_5_n79 , _add_98_5_n78 , _add_98_5_n77 , _add_98_5_n76 ,_add_98_5_n75 , _add_98_5_n74 , _add_98_5_n73 , _add_98_5_n72 ,_add_98_5_n71 , _add_98_5_n70 , _add_98_5_n69 , _add_98_5_n68 ,_add_98_5_n67 , _add_98_5_n66 , _add_98_5_n65 , _add_98_5_n64 ,_add_98_5_n63 , _add_98_5_n62 , _add_98_5_n61 , _add_98_5_n60 ,_add_98_5_n59 , _add_98_5_n58 , _add_98_5_n57 , _add_98_5_n56 ,_add_98_5_n55 , _add_98_5_n54 , _add_98_5_n53 , _add_98_5_n52 ,_add_98_5_n51 , _add_98_5_n50 , _add_98_5_n49 , _add_98_5_n48 ,_add_98_5_n47 , _add_98_5_n46 , _add_98_5_n45 , _add_98_5_n44 ,_add_98_5_n43 , _add_98_5_n42 , _add_98_5_n41 , _add_98_5_n40 ,_add_98_5_n39 , _add_98_5_n38 , _add_98_5_n37 , _add_98_5_n36 ,_add_98_5_n35 , _add_98_5_n34 , _add_98_5_n33 , _add_98_5_n32 ,_add_98_5_n31 , _add_98_5_n29 , _add_98_5_n28 , _add_98_5_n27 ,_add_98_5_n26 , _add_98_5_n25 , _add_98_5_n24 , _add_98_5_n23 ,_add_98_5_n22 , _add_98_5_n21 , _add_98_5_n20 , _add_98_5_n19 ,_add_98_5_n18 , _add_98_5_n17 , _add_98_5_n16 , _add_98_5_n15 ,_add_98_5_n14 , _add_98_5_n13 , _add_98_5_n12 , _add_98_5_n11 ,_add_98_5_n10 , _add_98_5_n9 , _add_98_5_n8 , _add_98_5_n7 ,_add_98_5_n6 , _add_98_5_n5 , _add_98_5_n4 , _add_98_5_n3 ,_add_98_5_n2 , _add_98_5_n1 , _add_98_n394 , _add_98_n393 ,_add_98_n392 , _add_98_n391 , _add_98_n390 , _add_98_n389 ,_add_98_n388 , _add_98_n387 , _add_98_n386 , _add_98_n385 ,_add_98_n384 , _add_98_n383 , _add_98_n382 , _add_98_n381 ,_add_98_n380 , _add_98_n379 , _add_98_n378 , _add_98_n377 ,_add_98_n376 , _add_98_n375 , _add_98_n374 , _add_98_n373 ,_add_98_n372 , _add_98_n371 , _add_98_n370 , _add_98_n369 ,_add_98_n368 , _add_98_n367 , _add_98_n366 , _add_98_n365 ,_add_98_n364 , _add_98_n363 , _add_98_n362 , _add_98_n361 ,_add_98_n360 , _add_98_n359 , _add_98_n358 , _add_98_n357 ,_add_98_n356 , _add_98_n355 , _add_98_n354 , _add_98_n353 ,_add_98_n352 , _add_98_n351 , _add_98_n350 , _add_98_n349 ,_add_98_n348 , _add_98_n347 , _add_98_n346 , _add_98_n345 ,_add_98_n344 , _add_98_n343 , _add_98_n342 , _add_98_n341 ,_add_98_n340 , _add_98_n339 , _add_98_n338 , _add_98_n337 ,_add_98_n336 , _add_98_n335 , _add_98_n334 , _add_98_n333 ,_add_98_n332 , _add_98_n331 , _add_98_n330 , _add_98_n329 ,_add_98_n328 , _add_98_n327 , _add_98_n326 , _add_98_n325 ,_add_98_n324 , _add_98_n323 , _add_98_n322 , _add_98_n321 ,_add_98_n320 , _add_98_n319 , _add_98_n318 , _add_98_n317 ,_add_98_n316 , _add_98_n315 , _add_98_n314 , _add_98_n313 ,_add_98_n312 , _add_98_n311 , _add_98_n310 , _add_98_n309 ,_add_98_n308 , _add_98_n307 , _add_98_n306 , _add_98_n305 ,_add_98_n304 , _add_98_n303 , _add_98_n302 , _add_98_n301 ,_add_98_n300 , _add_98_n299 , _add_98_n298 , _add_98_n297 ,_add_98_n296 , _add_98_n295 , _add_98_n294 , _add_98_n293 ,_add_98_n292 , _add_98_n291 , _add_98_n290 , _add_98_n289 ,_add_98_n288 , _add_98_n287 , _add_98_n286 , _add_98_n285 ,_add_98_n284 , _add_98_n283 , _add_98_n282 , _add_98_n281 ,_add_98_n280 , _add_98_n279 , _add_98_n278 , _add_98_n277 ,_add_98_n276 , _add_98_n275 , _add_98_n274 , _add_98_n273 ,_add_98_n272 , _add_98_n271 , _add_98_n270 , _add_98_n269 ,_add_98_n268 , _add_98_n267 , _add_98_n266 , _add_98_n265 ,_add_98_n264 , _add_98_n263 , _add_98_n262 , _add_98_n261 ,_add_98_n260 , _add_98_n259 , _add_98_n258 , _add_98_n257 ,_add_98_n256 , _add_98_n255 , _add_98_n254 , _add_98_n253 ,_add_98_n252 , _add_98_n251 , _add_98_n250 , _add_98_n249 ,_add_98_n248 , _add_98_n247 , _add_98_n246 , _add_98_n245 ,_add_98_n244 , _add_98_n243 , _add_98_n242 , _add_98_n241 ,_add_98_n240 , _add_98_n239 , _add_98_n238 , _add_98_n237 ,_add_98_n236 , _add_98_n235 , _add_98_n234 , _add_98_n233 ,_add_98_n232 , _add_98_n231 , _add_98_n230 , _add_98_n229 ,_add_98_n228 , _add_98_n227 , _add_98_n226 , _add_98_n225 ,_add_98_n224 , _add_98_n223 , _add_98_n222 , _add_98_n221 ,_add_98_n220 , _add_98_n219 , _add_98_n218 , _add_98_n217 ,_add_98_n216 , _add_98_n215 , _add_98_n214 , _add_98_n213 ,_add_98_n212 , _add_98_n211 , _add_98_n210 , _add_98_n209 ,_add_98_n208 , _add_98_n207 , _add_98_n206 , _add_98_n205 ,_add_98_n204 , _add_98_n203 , _add_98_n202 , _add_98_n201 ,_add_98_n200 , _add_98_n199 , _add_98_n198 , _add_98_n197 ,_add_98_n196 , _add_98_n195 , _add_98_n194 , _add_98_n193 ,_add_98_n192 , _add_98_n191 , _add_98_n190 , _add_98_n189 ,_add_98_n188 , _add_98_n187 , _add_98_n186 , _add_98_n185 ,_add_98_n184 , _add_98_n183 , _add_98_n182 , _add_98_n181 ,_add_98_n180 , _add_98_n179 , _add_98_n178 , _add_98_n177 ,_add_98_n176 , _add_98_n175 , _add_98_n174 , _add_98_n173 ,_add_98_n172 , _add_98_n171 , _add_98_n170 , _add_98_n169 ,_add_98_n168 , _add_98_n167 , _add_98_n166 , _add_98_n165 ,_add_98_n164 , _add_98_n163 , _add_98_n162 , _add_98_n161 ,_add_98_n160 , _add_98_n159 , _add_98_n158 , _add_98_n157 ,_add_98_n156 , _add_98_n155 , _add_98_n154 , _add_98_n153 ,_add_98_n152 , _add_98_n151 , _add_98_n150 , _add_98_n149 ,_add_98_n148 , _add_98_n147 , _add_98_n146 , _add_98_n145 ,_add_98_n144 , _add_98_n143 , _add_98_n142 , _add_98_n141 ,_add_98_n140 , _add_98_n139 , _add_98_n138 , _add_98_n137 ,_add_98_n136 , _add_98_n135 , _add_98_n134 , _add_98_n133 ,_add_98_n132 , _add_98_n131 , _add_98_n130 , _add_98_n129 ,_add_98_n128 , _add_98_n127 , _add_98_n126 , _add_98_n125 ,_add_98_n124 , _add_98_n123 , _add_98_n122 , _add_98_n121 ,_add_98_n120 , _add_98_n119 , _add_98_n118 , _add_98_n117 ,_add_98_n116 , _add_98_n115 , _add_98_n114 , _add_98_n113 ,_add_98_n112 , _add_98_n111 , _add_98_n110 , _add_98_n109 ,_add_98_n108 , _add_98_n107 , _add_98_n106 , _add_98_n105 ,_add_98_n104 , _add_98_n103 , _add_98_n102 , _add_98_n101 ,_add_98_n100 , _add_98_n99 , _add_98_n98 , _add_98_n97 , _add_98_n96 ,_add_98_n95 , _add_98_n94 , _add_98_n93 , _add_98_n92 , _add_98_n91 ,_add_98_n90 , _add_98_n89 , _add_98_n88 , _add_98_n87 , _add_98_n86 ,_add_98_n85 , _add_98_n84 , _add_98_n83 , _add_98_n82 , _add_98_n81 ,_add_98_n80 , _add_98_n79 , _add_98_n78 , _add_98_n77 , _add_98_n76 ,_add_98_n75 , _add_98_n74 , _add_98_n73 , _add_98_n72 , _add_98_n71 ,_add_98_n70 , _add_98_n69 , _add_98_n68 , _add_98_n67 , _add_98_n66 ,_add_98_n65 , _add_98_n64 , _add_98_n63 , _add_98_n62 , _add_98_n61 ,_add_98_n60 , _add_98_n59 , _add_98_n58 , _add_98_n57 , _add_98_n56 ,_add_98_n55 , _add_98_n54 , _add_98_n53 , _add_98_n52 , _add_98_n51 ,_add_98_n50 , _add_98_n49 , _add_98_n48 , _add_98_n47 , _add_98_n46 ,_add_98_n45 , _add_98_n44 , _add_98_n43 , _add_98_n42 , _add_98_n41 ,_add_98_n40 , _add_98_n39 , _add_98_n38 , _add_98_n37 , _add_98_n36 ,_add_98_n35 , _add_98_n34 , _add_98_n32 , _add_98_n31 , _add_98_n30 ,_add_98_n29 , _add_98_n28 , _add_98_n27 , _add_98_n26 , _add_98_n25 ,_add_98_n24 , _add_98_n23 , _add_98_n22 , _add_98_n21 , _add_98_n20 ,_add_98_n19 , _add_98_n18 , _add_98_n17 , _add_98_n16 , _add_98_n15 ,_add_98_n14 , _add_98_n13 , _add_98_n12 , _add_98_n11 , _add_98_n10 ,_add_98_n9 , _add_98_n8 , _add_98_n7 , _add_98_n6 , _add_98_n5 ,_add_98_n4 , _add_98_n3 , _add_98_n2 , _add_98_n1 , _add_98_4_n389 ,_add_98_4_n388 , _add_98_4_n387 , _add_98_4_n386 , _add_98_4_n385 ,_add_98_4_n384 , _add_98_4_n383 , _add_98_4_n382 , _add_98_4_n381 ,_add_98_4_n380 , _add_98_4_n379 , _add_98_4_n378 , _add_98_4_n377 ,_add_98_4_n376 , _add_98_4_n375 , _add_98_4_n374 , _add_98_4_n373 ,_add_98_4_n372 , _add_98_4_n371 , _add_98_4_n370 , _add_98_4_n369 ,_add_98_4_n368 , _add_98_4_n367 , _add_98_4_n366 , _add_98_4_n365 ,_add_98_4_n364 , _add_98_4_n363 , _add_98_4_n362 , _add_98_4_n361 ,_add_98_4_n360 , _add_98_4_n359 , _add_98_4_n358 , _add_98_4_n357 ,_add_98_4_n356 , _add_98_4_n355 , _add_98_4_n354 , _add_98_4_n353 ,_add_98_4_n352 , _add_98_4_n351 , _add_98_4_n350 , _add_98_4_n349 ,_add_98_4_n348 , _add_98_4_n347 , _add_98_4_n346 , _add_98_4_n345 ,_add_98_4_n344 , _add_98_4_n343 , _add_98_4_n342 , _add_98_4_n341 ,_add_98_4_n340 , _add_98_4_n339 , _add_98_4_n338 , _add_98_4_n337 ,_add_98_4_n336 , _add_98_4_n335 , _add_98_4_n334 , _add_98_4_n333 ,_add_98_4_n332 , _add_98_4_n331 , _add_98_4_n330 , _add_98_4_n329 ,_add_98_4_n328 , _add_98_4_n327 , _add_98_4_n326 , _add_98_4_n325 ,_add_98_4_n324 , _add_98_4_n323 , _add_98_4_n322 , _add_98_4_n321 ,_add_98_4_n320 , _add_98_4_n319 , _add_98_4_n318 , _add_98_4_n317 ,_add_98_4_n316 , _add_98_4_n315 , _add_98_4_n314 , _add_98_4_n313 ,_add_98_4_n312 , _add_98_4_n311 , _add_98_4_n310 , _add_98_4_n309 ,_add_98_4_n308 , _add_98_4_n307 , _add_98_4_n306 , _add_98_4_n305 ,_add_98_4_n304 , _add_98_4_n303 , _add_98_4_n302 , _add_98_4_n301 ,_add_98_4_n300 , _add_98_4_n299 , _add_98_4_n298 , _add_98_4_n297 ,_add_98_4_n296 , _add_98_4_n295 , _add_98_4_n294 , _add_98_4_n293 ,_add_98_4_n292 , _add_98_4_n291 , _add_98_4_n290 , _add_98_4_n289 ,_add_98_4_n288 , _add_98_4_n287 , _add_98_4_n286 , _add_98_4_n285 ,_add_98_4_n284 , _add_98_4_n283 , _add_98_4_n282 , _add_98_4_n281 ,_add_98_4_n280 , _add_98_4_n279 , _add_98_4_n278 , _add_98_4_n277 ,_add_98_4_n276 , _add_98_4_n275 , _add_98_4_n274 , _add_98_4_n273 ,_add_98_4_n272 , _add_98_4_n271 , _add_98_4_n270 , _add_98_4_n269 ,_add_98_4_n268 , _add_98_4_n267 , _add_98_4_n266 , _add_98_4_n265 ,_add_98_4_n264 , _add_98_4_n263 , _add_98_4_n262 , _add_98_4_n261 ,_add_98_4_n260 , _add_98_4_n259 , _add_98_4_n258 , _add_98_4_n257 ,_add_98_4_n256 , _add_98_4_n255 , _add_98_4_n254 , _add_98_4_n253 ,_add_98_4_n252 , _add_98_4_n251 , _add_98_4_n250 , _add_98_4_n249 ,_add_98_4_n248 , _add_98_4_n247 , _add_98_4_n246 , _add_98_4_n245 ,_add_98_4_n244 , _add_98_4_n243 , _add_98_4_n242 , _add_98_4_n241 ,_add_98_4_n240 , _add_98_4_n239 , _add_98_4_n238 , _add_98_4_n237 ,_add_98_4_n236 , _add_98_4_n235 , _add_98_4_n234 , _add_98_4_n233 ,_add_98_4_n232 , _add_98_4_n231 , _add_98_4_n230 , _add_98_4_n229 ,_add_98_4_n228 , _add_98_4_n227 , _add_98_4_n226 , _add_98_4_n225 ,_add_98_4_n224 , _add_98_4_n223 , _add_98_4_n222 , _add_98_4_n221 ,_add_98_4_n220 , _add_98_4_n219 , _add_98_4_n218 , _add_98_4_n217 ,_add_98_4_n216 , _add_98_4_n215 , _add_98_4_n214 , _add_98_4_n213 ,_add_98_4_n212 , _add_98_4_n211 , _add_98_4_n210 , _add_98_4_n209 ,_add_98_4_n208 , _add_98_4_n207 , _add_98_4_n206 , _add_98_4_n205 ,_add_98_4_n204 , _add_98_4_n203 , _add_98_4_n202 , _add_98_4_n201 ,_add_98_4_n200 , _add_98_4_n199 , _add_98_4_n198 , _add_98_4_n197 ,_add_98_4_n196 , _add_98_4_n195 , _add_98_4_n194 , _add_98_4_n193 ,_add_98_4_n192 , _add_98_4_n191 , _add_98_4_n190 , _add_98_4_n189 ,_add_98_4_n188 , _add_98_4_n187 , _add_98_4_n186 , _add_98_4_n185 ,_add_98_4_n184 , _add_98_4_n183 , _add_98_4_n182 , _add_98_4_n181 ,_add_98_4_n180 , _add_98_4_n179 , _add_98_4_n178 , _add_98_4_n177 ,_add_98_4_n176 , _add_98_4_n175 , _add_98_4_n174 , _add_98_4_n173 ,_add_98_4_n172 , _add_98_4_n171 , _add_98_4_n170 , _add_98_4_n169 ,_add_98_4_n168 , _add_98_4_n167 , _add_98_4_n166 , _add_98_4_n165 ,_add_98_4_n164 , _add_98_4_n163 , _add_98_4_n162 , _add_98_4_n161 ,_add_98_4_n160 , _add_98_4_n159 , _add_98_4_n158 , _add_98_4_n157 ,_add_98_4_n156 , _add_98_4_n155 , _add_98_4_n154 , _add_98_4_n153 ,_add_98_4_n152 , _add_98_4_n151 , _add_98_4_n150 , _add_98_4_n149 ,_add_98_4_n148 , _add_98_4_n147 , _add_98_4_n146 , _add_98_4_n145 ,_add_98_4_n144 , _add_98_4_n143 , _add_98_4_n142 , _add_98_4_n141 ,_add_98_4_n140 , _add_98_4_n139 , _add_98_4_n138 , _add_98_4_n137 ,_add_98_4_n136 , _add_98_4_n135 , _add_98_4_n134 , _add_98_4_n133 ,_add_98_4_n132 , _add_98_4_n131 , _add_98_4_n130 , _add_98_4_n129 ,_add_98_4_n128 , _add_98_4_n127 , _add_98_4_n126 , _add_98_4_n125 ,_add_98_4_n124 , _add_98_4_n123 , _add_98_4_n122 , _add_98_4_n121 ,_add_98_4_n120 , _add_98_4_n119 , _add_98_4_n118 , _add_98_4_n117 ,_add_98_4_n116 , _add_98_4_n115 , _add_98_4_n114 , _add_98_4_n113 ,_add_98_4_n112 , _add_98_4_n111 , _add_98_4_n110 , _add_98_4_n109 ,_add_98_4_n108 , _add_98_4_n107 , _add_98_4_n106 , _add_98_4_n105 ,_add_98_4_n104 , _add_98_4_n103 , _add_98_4_n102 , _add_98_4_n101 ,_add_98_4_n100 , _add_98_4_n99 , _add_98_4_n98 , _add_98_4_n97 ,_add_98_4_n96 , _add_98_4_n95 , _add_98_4_n94 , _add_98_4_n93 ,_add_98_4_n92 , _add_98_4_n91 , _add_98_4_n90 , _add_98_4_n89 ,_add_98_4_n88 , _add_98_4_n87 , _add_98_4_n86 , _add_98_4_n85 ,_add_98_4_n84 , _add_98_4_n83 , _add_98_4_n82 , _add_98_4_n81 ,_add_98_4_n80 , _add_98_4_n79 , _add_98_4_n78 , _add_98_4_n77 ,_add_98_4_n76 , _add_98_4_n75 , _add_98_4_n74 , _add_98_4_n73 ,_add_98_4_n72 , _add_98_4_n71 , _add_98_4_n70 , _add_98_4_n69 ,_add_98_4_n68 , _add_98_4_n67 , _add_98_4_n66 , _add_98_4_n65 ,_add_98_4_n64 , _add_98_4_n63 , _add_98_4_n62 , _add_98_4_n61 ,_add_98_4_n60 , _add_98_4_n59 , _add_98_4_n58 , _add_98_4_n57 ,_add_98_4_n56 , _add_98_4_n55 , _add_98_4_n54 , _add_98_4_n53 ,_add_98_4_n52 , _add_98_4_n51 , _add_98_4_n50 , _add_98_4_n49 ,_add_98_4_n48 , _add_98_4_n47 , _add_98_4_n46 , _add_98_4_n45 ,_add_98_4_n44 , _add_98_4_n43 , _add_98_4_n42 , _add_98_4_n41 ,_add_98_4_n40 , _add_98_4_n39 , _add_98_4_n38 , _add_98_4_n37 ,_add_98_4_n36 , _add_98_4_n35 , _add_98_4_n34 , _add_98_4_n33 ,_add_98_4_n32 , _add_98_4_n31 , _add_98_4_n30 , _add_98_4_n29 ,_add_98_4_n27 , _add_98_4_n26 , _add_98_4_n25 , _add_98_4_n24 ,_add_98_4_n23 , _add_98_4_n22 , _add_98_4_n21 , _add_98_4_n20 ,_add_98_4_n19 , _add_98_4_n18 , _add_98_4_n17 , _add_98_4_n16 ,_add_98_4_n15 , _add_98_4_n14 , _add_98_4_n13 , _add_98_4_n12 ,_add_98_4_n11 , _add_98_4_n10 , _add_98_4_n9 , _add_98_4_n8 ,_add_98_4_n7 , _add_98_4_n6 , _add_98_4_n5 , _add_98_4_n4 ,_add_98_4_n3 , _add_98_4_n2 , _add_98_4_n1 ;
wire   [6:0] rnd_cnt_q;
wire   [511:0] w_d;
wire   [479:0] w_q;
wire   [1:0] state;
wire   [31:0] w;
wire   [159:0] rnd_q;
wire   [159:0] sha1_round_wire;
wire   [159:0] rnd_d;
wire   [159:0] cv_d;
wire   [159:0] cv_q;
wire   [159:0] cv_next_d;
wire   [6:0] rnd_cnt_d;
wire   [1:0] next_state;
wire   [31:0] _sha1_round_f ;
NAND2_X2 U3406 ( .A1(w[9]), .A2(n7159), .ZN(n4656) );
NAND2_X2 U3407 ( .A1(w_q[9]), .A2(n7279), .ZN(n4655) );
NAND2_X2 U3409 ( .A1(n4660), .A2(n4661), .ZN(w_d[99]) );
NAND2_X2 U3410 ( .A1(w_q[67]), .A2(n7216), .ZN(n4661) );
NAND2_X2 U3411 ( .A1(w_q[99]), .A2(n7279), .ZN(n4660) );
NAND2_X2 U3412 ( .A1(n4663), .A2(n4664), .ZN(w_d[98]) );
NAND2_X2 U3413 ( .A1(w_q[66]), .A2(n7216), .ZN(n4664) );
NAND2_X2 U3414 ( .A1(w_q[98]), .A2(n7279), .ZN(n4663) );
NAND2_X2 U3415 ( .A1(n4665), .A2(n4666), .ZN(w_d[97]) );
NAND2_X2 U3416 ( .A1(w_q[65]), .A2(n7216), .ZN(n4666) );
NAND2_X2 U3417 ( .A1(w_q[97]), .A2(n7279), .ZN(n4665) );
NAND2_X2 U3418 ( .A1(n4667), .A2(n4668), .ZN(w_d[96]) );
NAND2_X2 U3419 ( .A1(w_q[64]), .A2(n7216), .ZN(n4668) );
NAND2_X2 U3420 ( .A1(w_q[96]), .A2(n7279), .ZN(n4667) );
NAND2_X2 U3422 ( .A1(w[8]), .A2(n7159), .ZN(n4671) );
NAND2_X2 U3423 ( .A1(w_q[8]), .A2(n7279), .ZN(n4670) );
NAND2_X2 U3426 ( .A1(w[7]), .A2(n7159), .ZN(n4674) );
NAND2_X2 U3427 ( .A1(w_q[7]), .A2(n7278), .ZN(n4673) );
NAND2_X2 U3430 ( .A1(w[6]), .A2(n7159), .ZN(n4677) );
NAND2_X2 U3431 ( .A1(w_q[6]), .A2(n7278), .ZN(n4676) );
NAND2_X2 U3433 ( .A1(n4678), .A2(n4679), .ZN(w_d[63]) );
NAND2_X2 U3434 ( .A1(w_q[31]), .A2(n7216), .ZN(n4679) );
NAND2_X2 U3435 ( .A1(w_q[63]), .A2(n7278), .ZN(n4678) );
NAND2_X2 U3436 ( .A1(n4680), .A2(n4681), .ZN(w_d[62]) );
NAND2_X2 U3437 ( .A1(w_q[30]), .A2(n7216), .ZN(n4681) );
NAND2_X2 U3438 ( .A1(w_q[62]), .A2(n7278), .ZN(n4680) );
NAND2_X2 U3439 ( .A1(n4682), .A2(n4683), .ZN(w_d[61]) );
NAND2_X2 U3440 ( .A1(w_q[29]), .A2(n7216), .ZN(n4683) );
NAND2_X2 U3441 ( .A1(w_q[61]), .A2(n7278), .ZN(n4682) );
NAND2_X2 U3442 ( .A1(n4684), .A2(n4685), .ZN(w_d[60]) );
NAND2_X2 U3443 ( .A1(w_q[28]), .A2(n7215), .ZN(n4685) );
NAND2_X2 U3444 ( .A1(w_q[60]), .A2(n7278), .ZN(n4684) );
NAND2_X2 U3446 ( .A1(w[5]), .A2(n7159), .ZN(n4688) );
NAND2_X2 U3447 ( .A1(w_q[5]), .A2(n7278), .ZN(n4687) );
NAND2_X2 U3449 ( .A1(n4689), .A2(n4690), .ZN(w_d[59]) );
NAND2_X2 U3450 ( .A1(w_q[27]), .A2(n7215), .ZN(n4690) );
NAND2_X2 U3451 ( .A1(w_q[59]), .A2(n7278), .ZN(n4689) );
NAND2_X2 U3452 ( .A1(n4691), .A2(n4692), .ZN(w_d[58]) );
NAND2_X2 U3453 ( .A1(w_q[26]), .A2(n7215), .ZN(n4692) );
NAND2_X2 U3454 ( .A1(w_q[58]), .A2(n7278), .ZN(n4691) );
NAND2_X2 U3455 ( .A1(n4693), .A2(n4694), .ZN(w_d[57]) );
NAND2_X2 U3456 ( .A1(w_q[25]), .A2(n7215), .ZN(n4694) );
NAND2_X2 U3457 ( .A1(w_q[57]), .A2(n7278), .ZN(n4693) );
NAND2_X2 U3458 ( .A1(n4695), .A2(n4696), .ZN(w_d[56]) );
NAND2_X2 U3459 ( .A1(w_q[24]), .A2(n7215), .ZN(n4696) );
NAND2_X2 U3460 ( .A1(w_q[56]), .A2(n7278), .ZN(n4695) );
NAND2_X2 U3461 ( .A1(n4697), .A2(n4698), .ZN(w_d[55]) );
NAND2_X2 U3462 ( .A1(w_q[23]), .A2(n7215), .ZN(n4698) );
NAND2_X2 U3463 ( .A1(w_q[55]), .A2(n7277), .ZN(n4697) );
NAND2_X2 U3464 ( .A1(n4699), .A2(n4700), .ZN(w_d[54]) );
NAND2_X2 U3465 ( .A1(w_q[22]), .A2(n7215), .ZN(n4700) );
NAND2_X2 U3466 ( .A1(w_q[54]), .A2(n7277), .ZN(n4699) );
NAND2_X2 U3467 ( .A1(n4701), .A2(n4702), .ZN(w_d[53]) );
NAND2_X2 U3468 ( .A1(w_q[21]), .A2(n7215), .ZN(n4702) );
NAND2_X2 U3469 ( .A1(w_q[53]), .A2(n7277), .ZN(n4701) );
NAND2_X2 U3470 ( .A1(n4703), .A2(n4704), .ZN(w_d[52]) );
NAND2_X2 U3471 ( .A1(w_q[20]), .A2(n7215), .ZN(n4704) );
NAND2_X2 U3472 ( .A1(w_q[52]), .A2(n7277), .ZN(n4703) );
NAND2_X2 U3473 ( .A1(n4705), .A2(n4706), .ZN(w_d[51]) );
NAND2_X2 U3474 ( .A1(w_q[19]), .A2(n7215), .ZN(n4706) );
NAND2_X2 U3475 ( .A1(w_q[51]), .A2(n7277), .ZN(n4705) );
NAND2_X2 U3476 ( .A1(n4707), .A2(n4708), .ZN(w_d[511]) );
NAND2_X2 U3477 ( .A1(n7179), .A2(n4709), .ZN(n4708) );
XOR2_X2 U3478 ( .A(n4710), .B(n4711), .Z(n4709) );
XOR2_X2 U3479 ( .A(w_d[254]), .B(n4712), .Z(n4711) );
XOR2_X2 U3480 ( .A(w_d[94]), .B(w_d[446]), .Z(n4710) );
NAND2_X2 U3481 ( .A1(n4713), .A2(n4714), .ZN(w_d[94]) );
NAND2_X2 U3482 ( .A1(w_q[62]), .A2(n7215), .ZN(n4714) );
NAND2_X2 U3483 ( .A1(w_q[94]), .A2(n7277), .ZN(n4713) );
NAND2_X2 U3484 ( .A1(n4715), .A2(n7181), .ZN(n4707) );
NAND2_X2 U3485 ( .A1(n4717), .A2(n4718), .ZN(w_d[510]) );
NAND2_X2 U3486 ( .A1(n7179), .A2(n4719), .ZN(n4718) );
XOR2_X2 U3487 ( .A(n4720), .B(n4721), .Z(n4719) );
XOR2_X2 U3488 ( .A(w_d[253]), .B(n4722), .Z(n4721) );
XOR2_X2 U3489 ( .A(w_d[93]), .B(w_d[445]), .Z(n4720) );
NAND2_X2 U3490 ( .A1(n4723), .A2(n4724), .ZN(w_d[93]) );
NAND2_X2 U3491 ( .A1(w_q[61]), .A2(n7220), .ZN(n4724) );
NAND2_X2 U3492 ( .A1(w_q[93]), .A2(n7277), .ZN(n4723) );
NAND2_X2 U3493 ( .A1(n4712), .A2(n7181), .ZN(n4717) );
NAND2_X2 U3494 ( .A1(n4725), .A2(n4726), .ZN(n4712) );
NAND2_X2 U3495 ( .A1(w_q[478]), .A2(n7225), .ZN(n4726) );
NAND2_X2 U3496 ( .A1(w[30]), .A2(n7277), .ZN(n4725) );
NAND2_X2 U3497 ( .A1(n4727), .A2(n4728), .ZN(w_d[50]) );
NAND2_X2 U3498 ( .A1(w_q[18]), .A2(n7196), .ZN(n4728) );
NAND2_X2 U3499 ( .A1(w_q[50]), .A2(n7277), .ZN(n4727) );
NAND2_X2 U3500 ( .A1(n4729), .A2(n4730), .ZN(w_d[509]) );
NAND2_X2 U3501 ( .A1(n7179), .A2(n4731), .ZN(n4730) );
XOR2_X2 U3502 ( .A(n4732), .B(n4733), .Z(n4731) );
XOR2_X2 U3503 ( .A(w_d[252]), .B(n4734), .Z(n4733) );
XOR2_X2 U3504 ( .A(w_d[92]), .B(w_d[444]), .Z(n4732) );
NAND2_X2 U3505 ( .A1(n4735), .A2(n4736), .ZN(w_d[92]) );
NAND2_X2 U3506 ( .A1(w_q[60]), .A2(n7219), .ZN(n4736) );
NAND2_X2 U3507 ( .A1(w_q[92]), .A2(n7277), .ZN(n4735) );
NAND2_X2 U3508 ( .A1(n4722), .A2(n7181), .ZN(n4729) );
NAND2_X2 U3509 ( .A1(n4737), .A2(n4738), .ZN(n4722) );
NAND2_X2 U3510 ( .A1(w_q[477]), .A2(n7224), .ZN(n4738) );
NAND2_X2 U3511 ( .A1(w[29]), .A2(n7277), .ZN(n4737) );
NAND2_X2 U3512 ( .A1(n4739), .A2(n4740), .ZN(w_d[508]) );
NAND2_X2 U3513 ( .A1(n7179), .A2(n4741), .ZN(n4740) );
XOR2_X2 U3514 ( .A(n4742), .B(n4743), .Z(n4741) );
XOR2_X2 U3515 ( .A(w_d[251]), .B(n4744), .Z(n4743) );
XOR2_X2 U3516 ( .A(w_d[91]), .B(w_d[443]), .Z(n4742) );
NAND2_X2 U3517 ( .A1(n4745), .A2(n4746), .ZN(w_d[91]) );
NAND2_X2 U3518 ( .A1(w_q[59]), .A2(n7226), .ZN(n4746) );
NAND2_X2 U3519 ( .A1(w_q[91]), .A2(n7236), .ZN(n4745) );
NAND2_X2 U3520 ( .A1(n4734), .A2(n7181), .ZN(n4739) );
NAND2_X2 U3521 ( .A1(n4747), .A2(n4748), .ZN(n4734) );
NAND2_X2 U3522 ( .A1(w_q[476]), .A2(n7223), .ZN(n4748) );
NAND2_X2 U3523 ( .A1(w[28]), .A2(n7231), .ZN(n4747) );
NAND2_X2 U3524 ( .A1(n4749), .A2(n4750), .ZN(w_d[507]) );
NAND2_X2 U3525 ( .A1(n7179), .A2(n4751), .ZN(n4750) );
XOR2_X2 U3526 ( .A(n4752), .B(n4753), .Z(n4751) );
XOR2_X2 U3527 ( .A(w_d[250]), .B(n4754), .Z(n4753) );
XOR2_X2 U3528 ( .A(w_d[90]), .B(w_d[442]), .Z(n4752) );
NAND2_X2 U3529 ( .A1(n4755), .A2(n4756), .ZN(w_d[90]) );
NAND2_X2 U3530 ( .A1(w_q[58]), .A2(n7220), .ZN(n4756) );
NAND2_X2 U3531 ( .A1(w_q[90]), .A2(n7232), .ZN(n4755) );
NAND2_X2 U3532 ( .A1(n4744), .A2(n7181), .ZN(n4749) );
NAND2_X2 U3533 ( .A1(n4757), .A2(n4758), .ZN(n4744) );
NAND2_X2 U3534 ( .A1(w_q[475]), .A2(n7222), .ZN(n4758) );
NAND2_X2 U3535 ( .A1(w[27]), .A2(n7233), .ZN(n4757) );
NAND2_X2 U3536 ( .A1(n4759), .A2(n4760), .ZN(w_d[506]) );
NAND2_X2 U3537 ( .A1(n7179), .A2(n4761), .ZN(n4760) );
XOR2_X2 U3538 ( .A(n4762), .B(n4763), .Z(n4761) );
XOR2_X2 U3539 ( .A(w_d[249]), .B(n4764), .Z(n4763) );
XOR2_X2 U3540 ( .A(w_d[89]), .B(w_d[441]), .Z(n4762) );
NAND2_X2 U3541 ( .A1(n4765), .A2(n4766), .ZN(w_d[89]) );
NAND2_X2 U3542 ( .A1(w_q[57]), .A2(n7219), .ZN(n4766) );
NAND2_X2 U3543 ( .A1(w_q[89]), .A2(n7236), .ZN(n4765) );
NAND2_X2 U3544 ( .A1(n4754), .A2(n7181), .ZN(n4759) );
NAND2_X2 U3545 ( .A1(n4767), .A2(n4768), .ZN(n4754) );
NAND2_X2 U3546 ( .A1(w_q[474]), .A2(n7221), .ZN(n4768) );
NAND2_X2 U3547 ( .A1(w[26]), .A2(n7234), .ZN(n4767) );
NAND2_X2 U3548 ( .A1(n4769), .A2(n4770), .ZN(w_d[505]) );
NAND2_X2 U3549 ( .A1(n7179), .A2(n4771), .ZN(n4770) );
XOR2_X2 U3550 ( .A(n4772), .B(n4773), .Z(n4771) );
XOR2_X2 U3551 ( .A(w_d[248]), .B(n4774), .Z(n4773) );
XOR2_X2 U3552 ( .A(w_d[88]), .B(w_d[440]), .Z(n4772) );
NAND2_X2 U3553 ( .A1(n4775), .A2(n4776), .ZN(w_d[88]) );
NAND2_X2 U3554 ( .A1(w_q[56]), .A2(n7219), .ZN(n4776) );
NAND2_X2 U3555 ( .A1(w_q[88]), .A2(n7235), .ZN(n4775) );
NAND2_X2 U3556 ( .A1(n4764), .A2(n7181), .ZN(n4769) );
NAND2_X2 U3557 ( .A1(n4777), .A2(n4778), .ZN(n4764) );
NAND2_X2 U3558 ( .A1(w_q[473]), .A2(n7225), .ZN(n4778) );
NAND2_X2 U3559 ( .A1(w[25]), .A2(n7238), .ZN(n4777) );
NAND2_X2 U3560 ( .A1(n4779), .A2(n4780), .ZN(w_d[504]) );
NAND2_X2 U3561 ( .A1(n7179), .A2(n4781), .ZN(n4780) );
XOR2_X2 U3562 ( .A(n4782), .B(n4783), .Z(n4781) );
XOR2_X2 U3563 ( .A(w_d[247]), .B(n4784), .Z(n4783) );
XOR2_X2 U3564 ( .A(w_d[87]), .B(w_d[439]), .Z(n4782) );
NAND2_X2 U3565 ( .A1(n4785), .A2(n4786), .ZN(w_d[87]) );
NAND2_X2 U3566 ( .A1(w_q[55]), .A2(n7226), .ZN(n4786) );
NAND2_X2 U3567 ( .A1(w_q[87]), .A2(n7238), .ZN(n4785) );
NAND2_X2 U3568 ( .A1(n4774), .A2(n7181), .ZN(n4779) );
NAND2_X2 U3569 ( .A1(n4787), .A2(n4788), .ZN(n4774) );
NAND2_X2 U3570 ( .A1(w_q[472]), .A2(n7224), .ZN(n4788) );
NAND2_X2 U3571 ( .A1(w[24]), .A2(n7230), .ZN(n4787) );
NAND2_X2 U3572 ( .A1(n4789), .A2(n4790), .ZN(w_d[503]) );
NAND2_X2 U3573 ( .A1(n7179), .A2(n4791), .ZN(n4790) );
XOR2_X2 U3574 ( .A(n4792), .B(n4793), .Z(n4791) );
XOR2_X2 U3575 ( .A(w_d[246]), .B(n4794), .Z(n4793) );
XOR2_X2 U3576 ( .A(w_d[86]), .B(w_d[438]), .Z(n4792) );
NAND2_X2 U3577 ( .A1(n4795), .A2(n4796), .ZN(w_d[86]) );
NAND2_X2 U3578 ( .A1(w_q[54]), .A2(n7219), .ZN(n4796) );
NAND2_X2 U3579 ( .A1(w_q[86]), .A2(n7236), .ZN(n4795) );
NAND2_X2 U3580 ( .A1(n4784), .A2(n7181), .ZN(n4789) );
NAND2_X2 U3581 ( .A1(n4797), .A2(n4798), .ZN(n4784) );
NAND2_X2 U3582 ( .A1(w_q[471]), .A2(n7223), .ZN(n4798) );
NAND2_X2 U3583 ( .A1(w[23]), .A2(n7276), .ZN(n4797) );
NAND2_X2 U3584 ( .A1(n4799), .A2(n4800), .ZN(w_d[502]) );
NAND2_X2 U3585 ( .A1(n7179), .A2(n4801), .ZN(n4800) );
XOR2_X2 U3586 ( .A(n4802), .B(n4803), .Z(n4801) );
XOR2_X2 U3587 ( .A(w_d[245]), .B(n4804), .Z(n4803) );
XOR2_X2 U3588 ( .A(w_d[85]), .B(w_d[437]), .Z(n4802) );
NAND2_X2 U3589 ( .A1(n4805), .A2(n4806), .ZN(w_d[85]) );
NAND2_X2 U3590 ( .A1(w_q[53]), .A2(n7220), .ZN(n4806) );
NAND2_X2 U3591 ( .A1(w_q[85]), .A2(n7276), .ZN(n4805) );
NAND2_X2 U3592 ( .A1(n4794), .A2(n7181), .ZN(n4799) );
NAND2_X2 U3593 ( .A1(n4807), .A2(n4808), .ZN(n4794) );
NAND2_X2 U3594 ( .A1(w_q[470]), .A2(n7222), .ZN(n4808) );
NAND2_X2 U3595 ( .A1(w[22]), .A2(n7276), .ZN(n4807) );
NAND2_X2 U3596 ( .A1(n4809), .A2(n4810), .ZN(w_d[501]) );
NAND2_X2 U3597 ( .A1(n7178), .A2(n4811), .ZN(n4810) );
XOR2_X2 U3598 ( .A(n4812), .B(n4813), .Z(n4811) );
XOR2_X2 U3599 ( .A(w_d[244]), .B(n4814), .Z(n4813) );
XOR2_X2 U3600 ( .A(w_d[84]), .B(w_d[436]), .Z(n4812) );
NAND2_X2 U3601 ( .A1(n4815), .A2(n4816), .ZN(w_d[84]) );
NAND2_X2 U3602 ( .A1(w_q[52]), .A2(n7226), .ZN(n4816) );
NAND2_X2 U3603 ( .A1(w_q[84]), .A2(n7276), .ZN(n4815) );
NAND2_X2 U3604 ( .A1(n4804), .A2(n7181), .ZN(n4809) );
NAND2_X2 U3605 ( .A1(n4817), .A2(n4818), .ZN(n4804) );
NAND2_X2 U3606 ( .A1(w_q[469]), .A2(n7221), .ZN(n4818) );
NAND2_X2 U3607 ( .A1(w[21]), .A2(n7276), .ZN(n4817) );
NAND2_X2 U3608 ( .A1(n4819), .A2(n4820), .ZN(w_d[500]) );
NAND2_X2 U3609 ( .A1(n7178), .A2(n4821), .ZN(n4820) );
XOR2_X2 U3610 ( .A(n4822), .B(n4823), .Z(n4821) );
XOR2_X2 U3611 ( .A(w_d[243]), .B(n4824), .Z(n4823) );
XOR2_X2 U3612 ( .A(w_d[83]), .B(w_d[435]), .Z(n4822) );
NAND2_X2 U3613 ( .A1(n4825), .A2(n4826), .ZN(w_d[83]) );
NAND2_X2 U3614 ( .A1(w_q[51]), .A2(n7220), .ZN(n4826) );
NAND2_X2 U3615 ( .A1(w_q[83]), .A2(n7276), .ZN(n4825) );
NAND2_X2 U3616 ( .A1(n4814), .A2(n7180), .ZN(n4819) );
NAND2_X2 U3617 ( .A1(n4827), .A2(n4828), .ZN(n4814) );
NAND2_X2 U3618 ( .A1(w_q[468]), .A2(n7225), .ZN(n4828) );
NAND2_X2 U3619 ( .A1(w[20]), .A2(n7276), .ZN(n4827) );
NAND2_X2 U3621 ( .A1(w[4]), .A2(n7159), .ZN(n4831) );
NAND2_X2 U3622 ( .A1(w_q[4]), .A2(n7276), .ZN(n4830) );
NAND2_X2 U3624 ( .A1(n4832), .A2(n4833), .ZN(w_d[49]) );
NAND2_X2 U3625 ( .A1(w_q[17]), .A2(n7197), .ZN(n4833) );
NAND2_X2 U3626 ( .A1(w_q[49]), .A2(n7276), .ZN(n4832) );
NAND2_X2 U3627 ( .A1(n4834), .A2(n4835), .ZN(w_d[499]) );
NAND2_X2 U3628 ( .A1(n7178), .A2(n4836), .ZN(n4835) );
XOR2_X2 U3629 ( .A(n4837), .B(n4838), .Z(n4836) );
XOR2_X2 U3630 ( .A(w_d[242]), .B(n4839), .Z(n4838) );
XOR2_X2 U3631 ( .A(w_d[82]), .B(w_d[434]), .Z(n4837) );
NAND2_X2 U3632 ( .A1(n4840), .A2(n4841), .ZN(w_d[82]) );
NAND2_X2 U3633 ( .A1(w_q[50]), .A2(n7226), .ZN(n4841) );
NAND2_X2 U3634 ( .A1(w_q[82]), .A2(n7276), .ZN(n4840) );
NAND2_X2 U3635 ( .A1(n4824), .A2(n7180), .ZN(n4834) );
NAND2_X2 U3636 ( .A1(n4842), .A2(n4843), .ZN(n4824) );
NAND2_X2 U3637 ( .A1(w_q[467]), .A2(n7224), .ZN(n4843) );
NAND2_X2 U3638 ( .A1(w[19]), .A2(n7276), .ZN(n4842) );
NAND2_X2 U3639 ( .A1(n4844), .A2(n4845), .ZN(w_d[498]) );
NAND2_X2 U3640 ( .A1(n7178), .A2(n4846), .ZN(n4845) );
XOR2_X2 U3641 ( .A(n4847), .B(n4848), .Z(n4846) );
XOR2_X2 U3642 ( .A(w_d[241]), .B(n4849), .Z(n4848) );
XOR2_X2 U3643 ( .A(w_d[81]), .B(w_d[433]), .Z(n4847) );
NAND2_X2 U3644 ( .A1(n4850), .A2(n4851), .ZN(w_d[81]) );
NAND2_X2 U3645 ( .A1(w_q[49]), .A2(n7220), .ZN(n4851) );
NAND2_X2 U3646 ( .A1(w_q[81]), .A2(n7235), .ZN(n4850) );
NAND2_X2 U3647 ( .A1(n4839), .A2(n7180), .ZN(n4844) );
NAND2_X2 U3648 ( .A1(n4852), .A2(n4853), .ZN(n4839) );
NAND2_X2 U3649 ( .A1(w_q[466]), .A2(n7221), .ZN(n4853) );
NAND2_X2 U3650 ( .A1(w[18]), .A2(n7230), .ZN(n4852) );
NAND2_X2 U3651 ( .A1(n4854), .A2(n4855), .ZN(w_d[497]) );
NAND2_X2 U3652 ( .A1(n7178), .A2(n4856), .ZN(n4855) );
XOR2_X2 U3653 ( .A(n4857), .B(n4858), .Z(n4856) );
XOR2_X2 U3654 ( .A(w_d[240]), .B(n4859), .Z(n4858) );
XOR2_X2 U3655 ( .A(w_d[80]), .B(w_d[432]), .Z(n4857) );
NAND2_X2 U3656 ( .A1(n4860), .A2(n4861), .ZN(w_d[80]) );
NAND2_X2 U3657 ( .A1(w_q[48]), .A2(n7219), .ZN(n4861) );
NAND2_X2 U3658 ( .A1(w_q[80]), .A2(n7236), .ZN(n4860) );
NAND2_X2 U3659 ( .A1(n4849), .A2(n7180), .ZN(n4854) );
NAND2_X2 U3660 ( .A1(n4862), .A2(n4863), .ZN(n4849) );
NAND2_X2 U3661 ( .A1(w_q[465]), .A2(n7223), .ZN(n4863) );
NAND2_X2 U3662 ( .A1(w[17]), .A2(n7233), .ZN(n4862) );
NAND2_X2 U3663 ( .A1(n4864), .A2(n4865), .ZN(w_d[496]) );
NAND2_X2 U3664 ( .A1(n7178), .A2(n4866), .ZN(n4865) );
XOR2_X2 U3665 ( .A(n4867), .B(n4868), .Z(n4866) );
XOR2_X2 U3666 ( .A(w_d[239]), .B(n4869), .Z(n4868) );
XOR2_X2 U3667 ( .A(w_d[79]), .B(w_d[431]), .Z(n4867) );
NAND2_X2 U3668 ( .A1(n4870), .A2(n4871), .ZN(w_d[79]) );
NAND2_X2 U3669 ( .A1(w_q[47]), .A2(n7226), .ZN(n4871) );
NAND2_X2 U3670 ( .A1(w_q[79]), .A2(n7231), .ZN(n4870) );
NAND2_X2 U3671 ( .A1(n4859), .A2(n7180), .ZN(n4864) );
NAND2_X2 U3672 ( .A1(n4872), .A2(n4873), .ZN(n4859) );
NAND2_X2 U3673 ( .A1(w_q[464]), .A2(n7222), .ZN(n4873) );
NAND2_X2 U3674 ( .A1(w[16]), .A2(n7234), .ZN(n4872) );
NAND2_X2 U3675 ( .A1(n4874), .A2(n4875), .ZN(w_d[495]) );
NAND2_X2 U3676 ( .A1(n7178), .A2(n4876), .ZN(n4875) );
XOR2_X2 U3677 ( .A(n4877), .B(n4878), .Z(n4876) );
XOR2_X2 U3678 ( .A(w_d[238]), .B(n4879), .Z(n4878) );
XOR2_X2 U3679 ( .A(w_d[78]), .B(w_d[430]), .Z(n4877) );
NAND2_X2 U3680 ( .A1(n4880), .A2(n4881), .ZN(w_d[78]) );
NAND2_X2 U3681 ( .A1(w_q[46]), .A2(n7220), .ZN(n4881) );
NAND2_X2 U3682 ( .A1(w_q[78]), .A2(n7235), .ZN(n4880) );
NAND2_X2 U3683 ( .A1(n4869), .A2(n7180), .ZN(n4874) );
NAND2_X2 U3684 ( .A1(n4882), .A2(n4883), .ZN(n4869) );
NAND2_X2 U3685 ( .A1(w_q[463]), .A2(n7224), .ZN(n4883) );
NAND2_X2 U3686 ( .A1(w[15]), .A2(n7234), .ZN(n4882) );
NAND2_X2 U3687 ( .A1(n4884), .A2(n4885), .ZN(w_d[494]) );
NAND2_X2 U3688 ( .A1(n7178), .A2(n4886), .ZN(n4885) );
XOR2_X2 U3689 ( .A(n4887), .B(n4888), .Z(n4886) );
XOR2_X2 U3690 ( .A(w_d[237]), .B(n4889), .Z(n4888) );
XOR2_X2 U3691 ( .A(w_d[77]), .B(w_d[429]), .Z(n4887) );
NAND2_X2 U3692 ( .A1(n4890), .A2(n4891), .ZN(w_d[77]) );
NAND2_X2 U3693 ( .A1(w_q[45]), .A2(n7221), .ZN(n4891) );
NAND2_X2 U3694 ( .A1(w_q[77]), .A2(n7236), .ZN(n4890) );
NAND2_X2 U3695 ( .A1(n4879), .A2(n7180), .ZN(n4884) );
NAND2_X2 U3696 ( .A1(n4892), .A2(n4893), .ZN(n4879) );
NAND2_X2 U3697 ( .A1(w_q[462]), .A2(n7223), .ZN(n4893) );
NAND2_X2 U3698 ( .A1(w[14]), .A2(n7232), .ZN(n4892) );
NAND2_X2 U3699 ( .A1(n4894), .A2(n4895), .ZN(w_d[493]) );
NAND2_X2 U3700 ( .A1(n7178), .A2(n4896), .ZN(n4895) );
XOR2_X2 U3701 ( .A(n4897), .B(n4898), .Z(n4896) );
XOR2_X2 U3702 ( .A(w_d[236]), .B(n4899), .Z(n4898) );
XOR2_X2 U3703 ( .A(w_d[76]), .B(w_d[428]), .Z(n4897) );
NAND2_X2 U3704 ( .A1(n4900), .A2(n4901), .ZN(w_d[76]) );
NAND2_X2 U3705 ( .A1(w_q[44]), .A2(n7223), .ZN(n4901) );
NAND2_X2 U3706 ( .A1(w_q[76]), .A2(n7238), .ZN(n4900) );
NAND2_X2 U3707 ( .A1(n4889), .A2(n7180), .ZN(n4894) );
NAND2_X2 U3708 ( .A1(n4902), .A2(n4903), .ZN(n4889) );
NAND2_X2 U3709 ( .A1(w_q[461]), .A2(n7222), .ZN(n4903) );
NAND2_X2 U3710 ( .A1(w[13]), .A2(n7235), .ZN(n4902) );
NAND2_X2 U3711 ( .A1(n4904), .A2(n4905), .ZN(w_d[492]) );
NAND2_X2 U3712 ( .A1(n7178), .A2(n4906), .ZN(n4905) );
XOR2_X2 U3713 ( .A(n4907), .B(n4908), .Z(n4906) );
XOR2_X2 U3714 ( .A(w_d[235]), .B(n4909), .Z(n4908) );
XOR2_X2 U3715 ( .A(w_d[75]), .B(w_d[427]), .Z(n4907) );
NAND2_X2 U3716 ( .A1(n4910), .A2(n4911), .ZN(w_d[75]) );
NAND2_X2 U3717 ( .A1(w_q[43]), .A2(n7222), .ZN(n4911) );
NAND2_X2 U3718 ( .A1(w_q[75]), .A2(n7231), .ZN(n4910) );
NAND2_X2 U3719 ( .A1(n4899), .A2(n7180), .ZN(n4904) );
NAND2_X2 U3720 ( .A1(n4912), .A2(n4913), .ZN(n4899) );
NAND2_X2 U3721 ( .A1(w_q[460]), .A2(n7225), .ZN(n4913) );
NAND2_X2 U3722 ( .A1(w[12]), .A2(n7230), .ZN(n4912) );
NAND2_X2 U3723 ( .A1(n4914), .A2(n4915), .ZN(w_d[491]) );
NAND2_X2 U3724 ( .A1(n7178), .A2(n4916), .ZN(n4915) );
XOR2_X2 U3725 ( .A(n4917), .B(n4918), .Z(n4916) );
XOR2_X2 U3726 ( .A(w_d[234]), .B(n4919), .Z(n4918) );
XOR2_X2 U3727 ( .A(w_d[74]), .B(w_d[426]), .Z(n4917) );
NAND2_X2 U3728 ( .A1(n4920), .A2(n4921), .ZN(w_d[74]) );
NAND2_X2 U3729 ( .A1(w_q[42]), .A2(n7225), .ZN(n4921) );
NAND2_X2 U3730 ( .A1(w_q[74]), .A2(n7232), .ZN(n4920) );
NAND2_X2 U3731 ( .A1(n4909), .A2(n7180), .ZN(n4914) );
NAND2_X2 U3732 ( .A1(n4922), .A2(n4923), .ZN(n4909) );
NAND2_X2 U3733 ( .A1(w_q[459]), .A2(n7221), .ZN(n4923) );
NAND2_X2 U3735 ( .A1(n4924), .A2(n4925), .ZN(w_d[490]) );
NAND2_X2 U3736 ( .A1(n7177), .A2(n4926), .ZN(n4925) );
XOR2_X2 U3737 ( .A(n4927), .B(n4928), .Z(n4926) );
XOR2_X2 U3738 ( .A(w_d[233]), .B(n4929), .Z(n4928) );
XOR2_X2 U3739 ( .A(w_d[73]), .B(w_d[425]), .Z(n4927) );
NAND2_X2 U3740 ( .A1(n4930), .A2(n4931), .ZN(w_d[73]) );
NAND2_X2 U3741 ( .A1(w_q[41]), .A2(n7219), .ZN(n4931) );
NAND2_X2 U3742 ( .A1(w_q[73]), .A2(n7235), .ZN(n4930) );
NAND2_X2 U3743 ( .A1(n4919), .A2(n7180), .ZN(n4924) );
NAND2_X2 U3744 ( .A1(n4932), .A2(n4933), .ZN(n4919) );
NAND2_X2 U3745 ( .A1(w_q[458]), .A2(n7224), .ZN(n4933) );
NAND2_X2 U3746 ( .A1(w[10]), .A2(n7234), .ZN(n4932) );
NAND2_X2 U3747 ( .A1(n4934), .A2(n4935), .ZN(w_d[48]) );
NAND2_X2 U3748 ( .A1(w_q[16]), .A2(n7212), .ZN(n4935) );
NAND2_X2 U3749 ( .A1(w_q[48]), .A2(n7273), .ZN(n4934) );
NAND2_X2 U3750 ( .A1(n4936), .A2(n4937), .ZN(w_d[489]) );
NAND2_X2 U3751 ( .A1(n7177), .A2(n4938), .ZN(n4937) );
XOR2_X2 U3752 ( .A(n4939), .B(n4940), .Z(n4938) );
XOR2_X2 U3753 ( .A(w_d[232]), .B(n4941), .Z(n4940) );
XOR2_X2 U3754 ( .A(w_d[72]), .B(w_d[424]), .Z(n4939) );
NAND2_X2 U3755 ( .A1(n4942), .A2(n4943), .ZN(w_d[72]) );
NAND2_X2 U3756 ( .A1(w_q[40]), .A2(n7226), .ZN(n4943) );
NAND2_X2 U3757 ( .A1(w_q[72]), .A2(n7236), .ZN(n4942) );
NAND2_X2 U3758 ( .A1(n4929), .A2(n7180), .ZN(n4936) );
NAND2_X2 U3759 ( .A1(n4944), .A2(n4945), .ZN(n4929) );
NAND2_X2 U3760 ( .A1(w_q[457]), .A2(n7221), .ZN(n4945) );
NAND2_X2 U3761 ( .A1(w[9]), .A2(n7233), .ZN(n4944) );
NAND2_X2 U3762 ( .A1(n4946), .A2(n4947), .ZN(w_d[488]) );
NAND2_X2 U3763 ( .A1(n7177), .A2(n4948), .ZN(n4947) );
XOR2_X2 U3764 ( .A(n4949), .B(n4950), .Z(n4948) );
XOR2_X2 U3765 ( .A(w_d[231]), .B(n4951), .Z(n4950) );
XOR2_X2 U3766 ( .A(w_d[71]), .B(w_d[423]), .Z(n4949) );
NAND2_X2 U3767 ( .A1(n4952), .A2(n4953), .ZN(w_d[71]) );
NAND2_X2 U3768 ( .A1(w_q[39]), .A2(n7220), .ZN(n4953) );
NAND2_X2 U3769 ( .A1(w_q[71]), .A2(n7231), .ZN(n4952) );
NAND2_X2 U3770 ( .A1(n4941), .A2(n7180), .ZN(n4946) );
NAND2_X2 U3771 ( .A1(n4954), .A2(n4955), .ZN(n4941) );
NAND2_X2 U3772 ( .A1(w_q[456]), .A2(n7224), .ZN(n4955) );
NAND2_X2 U3773 ( .A1(w[8]), .A2(n7230), .ZN(n4954) );
NAND2_X2 U3774 ( .A1(n4956), .A2(n4957), .ZN(w_d[487]) );
NAND2_X2 U3775 ( .A1(n7177), .A2(n4958), .ZN(n4957) );
XOR2_X2 U3776 ( .A(n4959), .B(n4960), .Z(n4958) );
XOR2_X2 U3777 ( .A(w_d[230]), .B(n4961), .Z(n4960) );
XOR2_X2 U3778 ( .A(w_d[70]), .B(w_d[422]), .Z(n4959) );
NAND2_X2 U3779 ( .A1(n4962), .A2(n4963), .ZN(w_d[70]) );
NAND2_X2 U3780 ( .A1(w_q[38]), .A2(n7219), .ZN(n4963) );
NAND2_X2 U3781 ( .A1(w_q[70]), .A2(n7236), .ZN(n4962) );
NAND2_X2 U3782 ( .A1(n4951), .A2(n7180), .ZN(n4956) );
NAND2_X2 U3783 ( .A1(n4964), .A2(n4965), .ZN(n4951) );
NAND2_X2 U3784 ( .A1(w_q[455]), .A2(n7225), .ZN(n4965) );
NAND2_X2 U3785 ( .A1(w[7]), .A2(n7233), .ZN(n4964) );
NAND2_X2 U3786 ( .A1(n4966), .A2(n4967), .ZN(w_d[486]) );
NAND2_X2 U3787 ( .A1(n7177), .A2(n4968), .ZN(n4967) );
XOR2_X2 U3788 ( .A(n4969), .B(n4970), .Z(n4968) );
XOR2_X2 U3789 ( .A(w_d[229]), .B(n4971), .Z(n4970) );
XOR2_X2 U3790 ( .A(w_d[69]), .B(w_d[421]), .Z(n4969) );
NAND2_X2 U3791 ( .A1(n4972), .A2(n4973), .ZN(w_d[69]) );
NAND2_X2 U3792 ( .A1(w_q[37]), .A2(n7221), .ZN(n4973) );
NAND2_X2 U3793 ( .A1(w_q[69]), .A2(n7238), .ZN(n4972) );
NAND2_X2 U3794 ( .A1(n4961), .A2(n7180), .ZN(n4966) );
NAND2_X2 U3795 ( .A1(n4974), .A2(n4975), .ZN(n4961) );
NAND2_X2 U3796 ( .A1(w_q[454]), .A2(n7223), .ZN(n4975) );
NAND2_X2 U3797 ( .A1(w[6]), .A2(n7234), .ZN(n4974) );
NAND2_X2 U3798 ( .A1(n4976), .A2(n4977), .ZN(w_d[485]) );
NAND2_X2 U3799 ( .A1(n7177), .A2(n4978), .ZN(n4977) );
XOR2_X2 U3800 ( .A(n4979), .B(n4980), .Z(n4978) );
XOR2_X2 U3801 ( .A(w_d[228]), .B(n4981), .Z(n4980) );
XOR2_X2 U3802 ( .A(w_d[68]), .B(w_d[420]), .Z(n4979) );
NAND2_X2 U3803 ( .A1(n4982), .A2(n4983), .ZN(w_d[68]) );
NAND2_X2 U3804 ( .A1(w_q[36]), .A2(n7224), .ZN(n4983) );
NAND2_X2 U3805 ( .A1(w_q[68]), .A2(n7230), .ZN(n4982) );
NAND2_X2 U3806 ( .A1(n4971), .A2(n7180), .ZN(n4976) );
NAND2_X2 U3807 ( .A1(n4984), .A2(n4985), .ZN(n4971) );
NAND2_X2 U3808 ( .A1(w_q[453]), .A2(n7222), .ZN(n4985) );
NAND2_X2 U3809 ( .A1(w[5]), .A2(n7232), .ZN(n4984) );
NAND2_X2 U3810 ( .A1(n4986), .A2(n4987), .ZN(w_d[484]) );
NAND2_X2 U3811 ( .A1(n7177), .A2(n4988), .ZN(n4987) );
XOR2_X2 U3812 ( .A(n4989), .B(n4990), .Z(n4988) );
XOR2_X2 U3813 ( .A(w_d[227]), .B(n4991), .Z(n4990) );
XOR2_X2 U3814 ( .A(w_d[67]), .B(w_d[419]), .Z(n4989) );
NAND2_X2 U3815 ( .A1(n4992), .A2(n4993), .ZN(w_d[67]) );
NAND2_X2 U3816 ( .A1(w_q[35]), .A2(n7217), .ZN(n4993) );
NAND2_X2 U3817 ( .A1(w_q[67]), .A2(n7232), .ZN(n4992) );
NAND2_X2 U3818 ( .A1(n4981), .A2(n7180), .ZN(n4986) );
NAND2_X2 U3819 ( .A1(n4994), .A2(n4995), .ZN(n4981) );
NAND2_X2 U3820 ( .A1(w_q[452]), .A2(n7217), .ZN(n4995) );
NAND2_X2 U3821 ( .A1(w[4]), .A2(n7233), .ZN(n4994) );
NAND2_X2 U3822 ( .A1(n4996), .A2(n4997), .ZN(w_d[483]) );
NAND2_X2 U3823 ( .A1(n7177), .A2(n4998), .ZN(n4997) );
XOR2_X2 U3824 ( .A(n4999), .B(n5000), .Z(n4998) );
XOR2_X2 U3825 ( .A(w_d[226]), .B(n5001), .Z(n5000) );
XOR2_X2 U3826 ( .A(w_d[66]), .B(w_d[418]), .Z(n4999) );
NAND2_X2 U3827 ( .A1(n5002), .A2(n5003), .ZN(w_d[66]) );
NAND2_X2 U3828 ( .A1(w_q[34]), .A2(n7217), .ZN(n5003) );
NAND2_X2 U3829 ( .A1(w_q[66]), .A2(n7235), .ZN(n5002) );
NAND2_X2 U3830 ( .A1(n4991), .A2(n7180), .ZN(n4996) );
NAND2_X2 U3831 ( .A1(n5004), .A2(n5005), .ZN(n4991) );
NAND2_X2 U3832 ( .A1(w_q[451]), .A2(n7217), .ZN(n5005) );
NAND2_X2 U3833 ( .A1(w[3]), .A2(n7231), .ZN(n5004) );
NAND2_X2 U3834 ( .A1(n5006), .A2(n5007), .ZN(w_d[482]) );
NAND2_X2 U3835 ( .A1(n7177), .A2(n5008), .ZN(n5007) );
XOR2_X2 U3836 ( .A(n5009), .B(n5010), .Z(n5008) );
XOR2_X2 U3837 ( .A(w_d[225]), .B(n5011), .Z(n5010) );
XOR2_X2 U3838 ( .A(w_d[65]), .B(w_d[417]), .Z(n5009) );
NAND2_X2 U3839 ( .A1(n5012), .A2(n5013), .ZN(w_d[65]) );
NAND2_X2 U3840 ( .A1(w_q[33]), .A2(n7217), .ZN(n5013) );
NAND2_X2 U3841 ( .A1(w_q[65]), .A2(n7275), .ZN(n5012) );
NAND2_X2 U3842 ( .A1(n5001), .A2(n7180), .ZN(n5006) );
NAND2_X2 U3843 ( .A1(n5014), .A2(n5015), .ZN(n5001) );
NAND2_X2 U3844 ( .A1(w_q[450]), .A2(n7217), .ZN(n5015) );
NAND2_X2 U3845 ( .A1(w[2]), .A2(n7275), .ZN(n5014) );
NAND2_X2 U3846 ( .A1(n5016), .A2(n5017), .ZN(w_d[481]) );
NAND2_X2 U3847 ( .A1(n7177), .A2(n5018), .ZN(n5017) );
XOR2_X2 U3848 ( .A(n5019), .B(n5020), .Z(n5018) );
XOR2_X2 U3849 ( .A(w_d[224]), .B(n5021), .Z(n5020) );
XOR2_X2 U3850 ( .A(w_d[64]), .B(w_d[416]), .Z(n5019) );
NAND2_X2 U3851 ( .A1(n5022), .A2(n5023), .ZN(w_d[64]) );
NAND2_X2 U3852 ( .A1(w_q[32]), .A2(n7225), .ZN(n5023) );
NAND2_X2 U3853 ( .A1(w_q[64]), .A2(n7275), .ZN(n5022) );
NAND2_X2 U3854 ( .A1(n5011), .A2(n7180), .ZN(n5016) );
NAND2_X2 U3855 ( .A1(n5024), .A2(n5025), .ZN(n5011) );
NAND2_X2 U3856 ( .A1(w_q[449]), .A2(n7217), .ZN(n5025) );
NAND2_X2 U3857 ( .A1(w[1]), .A2(n7275), .ZN(n5024) );
NAND2_X2 U3858 ( .A1(n5026), .A2(n5027), .ZN(w_d[480]) );
NAND2_X2 U3859 ( .A1(n5021), .A2(n7180), .ZN(n5027) );
NAND2_X2 U3860 ( .A1(n5028), .A2(n5029), .ZN(n5021) );
NAND2_X2 U3861 ( .A1(w_q[448]), .A2(n7217), .ZN(n5029) );
NAND2_X2 U3862 ( .A1(w[0]), .A2(n7275), .ZN(n5028) );
NAND2_X2 U3863 ( .A1(n7177), .A2(n5030), .ZN(n5026) );
XOR2_X2 U3864 ( .A(n5031), .B(n5032), .Z(n5030) );
XOR2_X2 U3865 ( .A(w_d[447]), .B(w_d[255]), .Z(n5032) );
XOR2_X2 U3866 ( .A(w_d[95]), .B(n4715), .Z(n5031) );
NAND2_X2 U3867 ( .A1(n5033), .A2(n5034), .ZN(n4715) );
NAND2_X2 U3868 ( .A1(w_q[479]), .A2(n7223), .ZN(n5034) );
NAND2_X2 U3869 ( .A1(w[31]), .A2(n7275), .ZN(n5033) );
NAND2_X2 U3870 ( .A1(n5035), .A2(n5036), .ZN(w_d[95]) );
NAND2_X2 U3871 ( .A1(w_q[63]), .A2(n7222), .ZN(n5036) );
NAND2_X2 U3872 ( .A1(w_q[95]), .A2(n7275), .ZN(n5035) );
NAND2_X2 U3875 ( .A1(n5039), .A2(n5040), .ZN(w_d[47]) );
NAND2_X2 U3876 ( .A1(w_q[15]), .A2(n7214), .ZN(n5040) );
NAND2_X2 U3877 ( .A1(w_q[47]), .A2(n7275), .ZN(n5039) );
NAND2_X2 U3878 ( .A1(n5041), .A2(n5042), .ZN(w_d[479]) );
NAND2_X2 U3879 ( .A1(w_q[447]), .A2(n7214), .ZN(n5042) );
NAND2_X2 U3880 ( .A1(w_q[479]), .A2(n7275), .ZN(n5041) );
NAND2_X2 U3881 ( .A1(n5043), .A2(n5044), .ZN(w_d[478]) );
NAND2_X2 U3882 ( .A1(w_q[446]), .A2(n7214), .ZN(n5044) );
NAND2_X2 U3883 ( .A1(w_q[478]), .A2(n7275), .ZN(n5043) );
NAND2_X2 U3884 ( .A1(n5045), .A2(n5046), .ZN(w_d[477]) );
NAND2_X2 U3885 ( .A1(w_q[445]), .A2(n7214), .ZN(n5046) );
NAND2_X2 U3886 ( .A1(w_q[477]), .A2(n7275), .ZN(n5045) );
NAND2_X2 U3887 ( .A1(n5047), .A2(n5048), .ZN(w_d[476]) );
NAND2_X2 U3888 ( .A1(w_q[444]), .A2(n7214), .ZN(n5048) );
NAND2_X2 U3889 ( .A1(w_q[476]), .A2(n7274), .ZN(n5047) );
NAND2_X2 U3890 ( .A1(n5049), .A2(n5050), .ZN(w_d[475]) );
NAND2_X2 U3891 ( .A1(w_q[443]), .A2(n7214), .ZN(n5050) );
NAND2_X2 U3892 ( .A1(w_q[475]), .A2(n7274), .ZN(n5049) );
NAND2_X2 U3893 ( .A1(n5051), .A2(n5052), .ZN(w_d[474]) );
NAND2_X2 U3894 ( .A1(w_q[442]), .A2(n7214), .ZN(n5052) );
NAND2_X2 U3895 ( .A1(w_q[474]), .A2(n7274), .ZN(n5051) );
NAND2_X2 U3896 ( .A1(n5053), .A2(n5054), .ZN(w_d[473]) );
NAND2_X2 U3897 ( .A1(w_q[441]), .A2(n7214), .ZN(n5054) );
NAND2_X2 U3898 ( .A1(w_q[473]), .A2(n7274), .ZN(n5053) );
NAND2_X2 U3899 ( .A1(n5055), .A2(n5056), .ZN(w_d[472]) );
NAND2_X2 U3900 ( .A1(w_q[440]), .A2(n7214), .ZN(n5056) );
NAND2_X2 U3901 ( .A1(w_q[472]), .A2(n7274), .ZN(n5055) );
NAND2_X2 U3902 ( .A1(n5057), .A2(n5058), .ZN(w_d[471]) );
NAND2_X2 U3903 ( .A1(w_q[439]), .A2(n7214), .ZN(n5058) );
NAND2_X2 U3904 ( .A1(w_q[471]), .A2(n7274), .ZN(n5057) );
NAND2_X2 U3905 ( .A1(n5059), .A2(n5060), .ZN(w_d[470]) );
NAND2_X2 U3906 ( .A1(w_q[438]), .A2(n7214), .ZN(n5060) );
NAND2_X2 U3907 ( .A1(w_q[470]), .A2(n7274), .ZN(n5059) );
NAND2_X2 U3908 ( .A1(n5061), .A2(n5062), .ZN(w_d[46]) );
NAND2_X2 U3909 ( .A1(w_q[14]), .A2(n7213), .ZN(n5062) );
NAND2_X2 U3910 ( .A1(w_q[46]), .A2(n7274), .ZN(n5061) );
NAND2_X2 U3911 ( .A1(n5063), .A2(n5064), .ZN(w_d[469]) );
NAND2_X2 U3912 ( .A1(w_q[437]), .A2(n7213), .ZN(n5064) );
NAND2_X2 U3913 ( .A1(w_q[469]), .A2(n7274), .ZN(n5063) );
NAND2_X2 U3914 ( .A1(n5065), .A2(n5066), .ZN(w_d[468]) );
NAND2_X2 U3915 ( .A1(w_q[436]), .A2(n7213), .ZN(n5066) );
NAND2_X2 U3916 ( .A1(w_q[468]), .A2(n7274), .ZN(n5065) );
NAND2_X2 U3917 ( .A1(n5067), .A2(n5068), .ZN(w_d[467]) );
NAND2_X2 U3918 ( .A1(w_q[435]), .A2(n7213), .ZN(n5068) );
NAND2_X2 U3919 ( .A1(w_q[467]), .A2(n7274), .ZN(n5067) );
NAND2_X2 U3920 ( .A1(n5069), .A2(n5070), .ZN(w_d[466]) );
NAND2_X2 U3921 ( .A1(w_q[434]), .A2(n7213), .ZN(n5070) );
NAND2_X2 U3922 ( .A1(w_q[466]), .A2(n7273), .ZN(n5069) );
NAND2_X2 U3923 ( .A1(n5071), .A2(n5072), .ZN(w_d[465]) );
NAND2_X2 U3924 ( .A1(w_q[433]), .A2(n7213), .ZN(n5072) );
NAND2_X2 U3925 ( .A1(w_q[465]), .A2(n7273), .ZN(n5071) );
NAND2_X2 U3926 ( .A1(n5073), .A2(n5074), .ZN(w_d[464]) );
NAND2_X2 U3927 ( .A1(w_q[432]), .A2(n7213), .ZN(n5074) );
NAND2_X2 U3928 ( .A1(w_q[464]), .A2(n7273), .ZN(n5073) );
NAND2_X2 U3929 ( .A1(n5075), .A2(n5076), .ZN(w_d[463]) );
NAND2_X2 U3930 ( .A1(w_q[431]), .A2(n7213), .ZN(n5076) );
NAND2_X2 U3931 ( .A1(w_q[463]), .A2(n7273), .ZN(n5075) );
NAND2_X2 U3932 ( .A1(n5077), .A2(n5078), .ZN(w_d[462]) );
NAND2_X2 U3933 ( .A1(w_q[430]), .A2(n7213), .ZN(n5078) );
NAND2_X2 U3934 ( .A1(w_q[462]), .A2(n7273), .ZN(n5077) );
NAND2_X2 U3935 ( .A1(n5079), .A2(n5080), .ZN(w_d[461]) );
NAND2_X2 U3936 ( .A1(w_q[429]), .A2(n7213), .ZN(n5080) );
NAND2_X2 U3937 ( .A1(w_q[461]), .A2(n7273), .ZN(n5079) );
NAND2_X2 U3938 ( .A1(n5081), .A2(n5082), .ZN(w_d[460]) );
NAND2_X2 U3939 ( .A1(w_q[428]), .A2(n7213), .ZN(n5082) );
NAND2_X2 U3940 ( .A1(w_q[460]), .A2(n7273), .ZN(n5081) );
NAND2_X2 U3941 ( .A1(n5083), .A2(n5084), .ZN(w_d[45]) );
NAND2_X2 U3942 ( .A1(w_q[13]), .A2(n7212), .ZN(n5084) );
NAND2_X2 U3943 ( .A1(w_q[45]), .A2(n7273), .ZN(n5083) );
NAND2_X2 U3944 ( .A1(n5085), .A2(n5086), .ZN(w_d[459]) );
NAND2_X2 U3945 ( .A1(w_q[427]), .A2(n7212), .ZN(n5086) );
NAND2_X2 U3946 ( .A1(w_q[459]), .A2(n7273), .ZN(n5085) );
NAND2_X2 U3947 ( .A1(n5087), .A2(n5088), .ZN(w_d[458]) );
NAND2_X2 U3948 ( .A1(w_q[426]), .A2(n7212), .ZN(n5088) );
NAND2_X2 U3949 ( .A1(w_q[458]), .A2(n7273), .ZN(n5087) );
NAND2_X2 U3950 ( .A1(n5089), .A2(n5090), .ZN(w_d[457]) );
NAND2_X2 U3951 ( .A1(w_q[425]), .A2(n7212), .ZN(n5090) );
NAND2_X2 U3952 ( .A1(w_q[457]), .A2(n7273), .ZN(n5089) );
NAND2_X2 U3953 ( .A1(n5091), .A2(n5092), .ZN(w_d[456]) );
NAND2_X2 U3954 ( .A1(w_q[424]), .A2(n7212), .ZN(n5092) );
NAND2_X2 U3955 ( .A1(w_q[456]), .A2(n7272), .ZN(n5091) );
NAND2_X2 U3956 ( .A1(n5093), .A2(n5094), .ZN(w_d[455]) );
NAND2_X2 U3957 ( .A1(w_q[423]), .A2(n7212), .ZN(n5094) );
NAND2_X2 U3958 ( .A1(w_q[455]), .A2(n7272), .ZN(n5093) );
NAND2_X2 U3959 ( .A1(n5095), .A2(n5096), .ZN(w_d[454]) );
NAND2_X2 U3960 ( .A1(w_q[422]), .A2(n7212), .ZN(n5096) );
NAND2_X2 U3961 ( .A1(w_q[454]), .A2(n7272), .ZN(n5095) );
NAND2_X2 U3962 ( .A1(n5097), .A2(n5098), .ZN(w_d[453]) );
NAND2_X2 U3963 ( .A1(w_q[421]), .A2(n7212), .ZN(n5098) );
NAND2_X2 U3964 ( .A1(w_q[453]), .A2(n7272), .ZN(n5097) );
NAND2_X2 U3965 ( .A1(n5099), .A2(n5100), .ZN(w_d[452]) );
NAND2_X2 U3966 ( .A1(w_q[420]), .A2(n7212), .ZN(n5100) );
NAND2_X2 U3967 ( .A1(w_q[452]), .A2(n7272), .ZN(n5099) );
NAND2_X2 U3968 ( .A1(n5101), .A2(n5102), .ZN(w_d[451]) );
NAND2_X2 U3969 ( .A1(w_q[419]), .A2(n7212), .ZN(n5102) );
NAND2_X2 U3970 ( .A1(w_q[451]), .A2(n7272), .ZN(n5101) );
NAND2_X2 U3971 ( .A1(n5103), .A2(n5104), .ZN(w_d[450]) );
NAND2_X2 U3972 ( .A1(w_q[418]), .A2(n7212), .ZN(n5104) );
NAND2_X2 U3973 ( .A1(w_q[450]), .A2(n7272), .ZN(n5103) );
NAND2_X2 U3974 ( .A1(n5105), .A2(n5106), .ZN(w_d[44]) );
NAND2_X2 U3975 ( .A1(w_q[12]), .A2(n7216), .ZN(n5106) );
NAND2_X2 U3976 ( .A1(w_q[44]), .A2(n7272), .ZN(n5105) );
NAND2_X2 U3977 ( .A1(n5107), .A2(n5108), .ZN(w_d[449]) );
NAND2_X2 U3978 ( .A1(w_q[417]), .A2(n7196), .ZN(n5108) );
NAND2_X2 U3979 ( .A1(w_q[449]), .A2(n7272), .ZN(n5107) );
NAND2_X2 U3980 ( .A1(n5109), .A2(n5110), .ZN(w_d[448]) );
NAND2_X2 U3981 ( .A1(w_q[416]), .A2(n7197), .ZN(n5110) );
NAND2_X2 U3982 ( .A1(w_q[448]), .A2(n7272), .ZN(n5109) );
NAND2_X2 U3983 ( .A1(n5111), .A2(n5112), .ZN(w_d[447]) );
NAND2_X2 U3984 ( .A1(w_q[415]), .A2(n7218), .ZN(n5112) );
NAND2_X2 U3985 ( .A1(w_q[447]), .A2(n7272), .ZN(n5111) );
NAND2_X2 U3986 ( .A1(n5113), .A2(n5114), .ZN(w_d[446]) );
NAND2_X2 U3987 ( .A1(w_q[414]), .A2(n7218), .ZN(n5114) );
NAND2_X2 U3988 ( .A1(w_q[446]), .A2(n7271), .ZN(n5113) );
NAND2_X2 U3989 ( .A1(n5115), .A2(n5116), .ZN(w_d[445]) );
NAND2_X2 U3990 ( .A1(w_q[413]), .A2(n7218), .ZN(n5116) );
NAND2_X2 U3991 ( .A1(w_q[445]), .A2(n7271), .ZN(n5115) );
NAND2_X2 U3992 ( .A1(n5117), .A2(n5118), .ZN(w_d[444]) );
NAND2_X2 U3993 ( .A1(w_q[412]), .A2(n7218), .ZN(n5118) );
NAND2_X2 U3994 ( .A1(w_q[444]), .A2(n7271), .ZN(n5117) );
NAND2_X2 U3995 ( .A1(n5119), .A2(n5120), .ZN(w_d[443]) );
NAND2_X2 U3996 ( .A1(w_q[411]), .A2(n7218), .ZN(n5120) );
NAND2_X2 U3997 ( .A1(w_q[443]), .A2(n7271), .ZN(n5119) );
NAND2_X2 U3998 ( .A1(n5121), .A2(n5122), .ZN(w_d[442]) );
NAND2_X2 U3999 ( .A1(w_q[410]), .A2(n7218), .ZN(n5122) );
NAND2_X2 U4000 ( .A1(w_q[442]), .A2(n7271), .ZN(n5121) );
NAND2_X2 U4001 ( .A1(n5123), .A2(n5124), .ZN(w_d[441]) );
NAND2_X2 U4002 ( .A1(w_q[409]), .A2(n7218), .ZN(n5124) );
NAND2_X2 U4003 ( .A1(w_q[441]), .A2(n7271), .ZN(n5123) );
NAND2_X2 U4004 ( .A1(n5125), .A2(n5126), .ZN(w_d[440]) );
NAND2_X2 U4005 ( .A1(w_q[408]), .A2(n7218), .ZN(n5126) );
NAND2_X2 U4006 ( .A1(w_q[440]), .A2(n7271), .ZN(n5125) );
NAND2_X2 U4007 ( .A1(n5127), .A2(n5128), .ZN(w_d[43]) );
NAND2_X2 U4008 ( .A1(w_q[11]), .A2(n7216), .ZN(n5128) );
NAND2_X2 U4009 ( .A1(w_q[43]), .A2(n7271), .ZN(n5127) );
NAND2_X2 U4010 ( .A1(n5129), .A2(n5130), .ZN(w_d[439]) );
NAND2_X2 U4011 ( .A1(w_q[407]), .A2(n7225), .ZN(n5130) );
NAND2_X2 U4012 ( .A1(w_q[439]), .A2(n7271), .ZN(n5129) );
NAND2_X2 U4013 ( .A1(n5131), .A2(n5132), .ZN(w_d[438]) );
NAND2_X2 U4014 ( .A1(w_q[406]), .A2(n7223), .ZN(n5132) );
NAND2_X2 U4015 ( .A1(w_q[438]), .A2(n7271), .ZN(n5131) );
NAND2_X2 U4016 ( .A1(n5133), .A2(n5134), .ZN(w_d[437]) );
NAND2_X2 U4017 ( .A1(w_q[405]), .A2(n7222), .ZN(n5134) );
NAND2_X2 U4018 ( .A1(w_q[437]), .A2(n7271), .ZN(n5133) );
NAND2_X2 U4019 ( .A1(n5135), .A2(n5136), .ZN(w_d[436]) );
NAND2_X2 U4020 ( .A1(w_q[404]), .A2(n7226), .ZN(n5136) );
NAND2_X2 U4021 ( .A1(w_q[436]), .A2(n7270), .ZN(n5135) );
NAND2_X2 U4022 ( .A1(n5137), .A2(n5138), .ZN(w_d[435]) );
NAND2_X2 U4023 ( .A1(w_q[403]), .A2(n7220), .ZN(n5138) );
NAND2_X2 U4024 ( .A1(w_q[435]), .A2(n7270), .ZN(n5137) );
NAND2_X2 U4025 ( .A1(n5139), .A2(n5140), .ZN(w_d[434]) );
NAND2_X2 U4026 ( .A1(w_q[402]), .A2(n7219), .ZN(n5140) );
NAND2_X2 U4027 ( .A1(w_q[434]), .A2(n7270), .ZN(n5139) );
NAND2_X2 U4028 ( .A1(n5141), .A2(n5142), .ZN(w_d[433]) );
NAND2_X2 U4029 ( .A1(w_q[401]), .A2(n7218), .ZN(n5142) );
NAND2_X2 U4030 ( .A1(w_q[433]), .A2(n7270), .ZN(n5141) );
NAND2_X2 U4031 ( .A1(n5143), .A2(n5144), .ZN(w_d[432]) );
NAND2_X2 U4032 ( .A1(w_q[400]), .A2(n7217), .ZN(n5144) );
NAND2_X2 U4033 ( .A1(w_q[432]), .A2(n7270), .ZN(n5143) );
NAND2_X2 U4034 ( .A1(n5145), .A2(n5146), .ZN(w_d[431]) );
NAND2_X2 U4035 ( .A1(w_q[399]), .A2(n7221), .ZN(n5146) );
NAND2_X2 U4036 ( .A1(w_q[431]), .A2(n7270), .ZN(n5145) );
NAND2_X2 U4037 ( .A1(n5147), .A2(n5148), .ZN(w_d[430]) );
NAND2_X2 U4038 ( .A1(w_q[398]), .A2(n7224), .ZN(n5148) );
NAND2_X2 U4039 ( .A1(w_q[430]), .A2(n7270), .ZN(n5147) );
NAND2_X2 U4040 ( .A1(n5149), .A2(n5150), .ZN(w_d[42]) );
NAND2_X2 U4041 ( .A1(w_q[10]), .A2(n7211), .ZN(n5150) );
NAND2_X2 U4042 ( .A1(w_q[42]), .A2(n7270), .ZN(n5149) );
NAND2_X2 U4043 ( .A1(n5151), .A2(n5152), .ZN(w_d[429]) );
NAND2_X2 U4044 ( .A1(w_q[397]), .A2(n7211), .ZN(n5152) );
NAND2_X2 U4045 ( .A1(w_q[429]), .A2(n7270), .ZN(n5151) );
NAND2_X2 U4046 ( .A1(n5153), .A2(n5154), .ZN(w_d[428]) );
NAND2_X2 U4047 ( .A1(w_q[396]), .A2(n7211), .ZN(n5154) );
NAND2_X2 U4048 ( .A1(w_q[428]), .A2(n7270), .ZN(n5153) );
NAND2_X2 U4049 ( .A1(n5155), .A2(n5156), .ZN(w_d[427]) );
NAND2_X2 U4050 ( .A1(w_q[395]), .A2(n7211), .ZN(n5156) );
NAND2_X2 U4051 ( .A1(w_q[427]), .A2(n7270), .ZN(n5155) );
NAND2_X2 U4052 ( .A1(n5157), .A2(n5158), .ZN(w_d[426]) );
NAND2_X2 U4053 ( .A1(w_q[394]), .A2(n7211), .ZN(n5158) );
NAND2_X2 U4054 ( .A1(w_q[426]), .A2(n7269), .ZN(n5157) );
NAND2_X2 U4055 ( .A1(n5159), .A2(n5160), .ZN(w_d[425]) );
NAND2_X2 U4056 ( .A1(w_q[393]), .A2(n7211), .ZN(n5160) );
NAND2_X2 U4057 ( .A1(w_q[425]), .A2(n7269), .ZN(n5159) );
NAND2_X2 U4058 ( .A1(n5161), .A2(n5162), .ZN(w_d[424]) );
NAND2_X2 U4059 ( .A1(w_q[392]), .A2(n7211), .ZN(n5162) );
NAND2_X2 U4060 ( .A1(w_q[424]), .A2(n7269), .ZN(n5161) );
NAND2_X2 U4061 ( .A1(n5163), .A2(n5164), .ZN(w_d[423]) );
NAND2_X2 U4062 ( .A1(w_q[391]), .A2(n7211), .ZN(n5164) );
NAND2_X2 U4063 ( .A1(w_q[423]), .A2(n7269), .ZN(n5163) );
NAND2_X2 U4064 ( .A1(n5165), .A2(n5166), .ZN(w_d[422]) );
NAND2_X2 U4065 ( .A1(w_q[390]), .A2(n7211), .ZN(n5166) );
NAND2_X2 U4066 ( .A1(w_q[422]), .A2(n7269), .ZN(n5165) );
NAND2_X2 U4067 ( .A1(n5167), .A2(n5168), .ZN(w_d[421]) );
NAND2_X2 U4068 ( .A1(w_q[389]), .A2(n7211), .ZN(n5168) );
NAND2_X2 U4069 ( .A1(w_q[421]), .A2(n7269), .ZN(n5167) );
NAND2_X2 U4070 ( .A1(n5169), .A2(n5170), .ZN(w_d[420]) );
NAND2_X2 U4071 ( .A1(w_q[388]), .A2(n7211), .ZN(n5170) );
NAND2_X2 U4072 ( .A1(w_q[420]), .A2(n7269), .ZN(n5169) );
NAND2_X2 U4073 ( .A1(n5171), .A2(n5172), .ZN(w_d[41]) );
NAND2_X2 U4074 ( .A1(w_q[9]), .A2(n7210), .ZN(n5172) );
NAND2_X2 U4075 ( .A1(w_q[41]), .A2(n7269), .ZN(n5171) );
NAND2_X2 U4076 ( .A1(n5173), .A2(n5174), .ZN(w_d[419]) );
NAND2_X2 U4077 ( .A1(w_q[387]), .A2(n7210), .ZN(n5174) );
NAND2_X2 U4078 ( .A1(w_q[419]), .A2(n7269), .ZN(n5173) );
NAND2_X2 U4079 ( .A1(n5175), .A2(n5176), .ZN(w_d[418]) );
NAND2_X2 U4080 ( .A1(w_q[386]), .A2(n7210), .ZN(n5176) );
NAND2_X2 U4081 ( .A1(w_q[418]), .A2(n7269), .ZN(n5175) );
NAND2_X2 U4082 ( .A1(n5177), .A2(n5178), .ZN(w_d[417]) );
NAND2_X2 U4083 ( .A1(w_q[385]), .A2(n7210), .ZN(n5178) );
NAND2_X2 U4084 ( .A1(w_q[417]), .A2(n7269), .ZN(n5177) );
NAND2_X2 U4085 ( .A1(n5179), .A2(n5180), .ZN(w_d[416]) );
NAND2_X2 U4086 ( .A1(w_q[384]), .A2(n7210), .ZN(n5180) );
NAND2_X2 U4087 ( .A1(w_q[416]), .A2(n7268), .ZN(n5179) );
NAND2_X2 U4088 ( .A1(n5181), .A2(n5182), .ZN(w_d[415]) );
NAND2_X2 U4089 ( .A1(w_q[383]), .A2(n7210), .ZN(n5182) );
NAND2_X2 U4090 ( .A1(w_q[415]), .A2(n7268), .ZN(n5181) );
NAND2_X2 U4091 ( .A1(n5183), .A2(n5184), .ZN(w_d[414]) );
NAND2_X2 U4092 ( .A1(w_q[382]), .A2(n7210), .ZN(n5184) );
NAND2_X2 U4093 ( .A1(w_q[414]), .A2(n7268), .ZN(n5183) );
NAND2_X2 U4094 ( .A1(n5185), .A2(n5186), .ZN(w_d[413]) );
NAND2_X2 U4095 ( .A1(w_q[381]), .A2(n7210), .ZN(n5186) );
NAND2_X2 U4096 ( .A1(w_q[413]), .A2(n7268), .ZN(n5185) );
NAND2_X2 U4097 ( .A1(n5187), .A2(n5188), .ZN(w_d[412]) );
NAND2_X2 U4098 ( .A1(w_q[380]), .A2(n7210), .ZN(n5188) );
NAND2_X2 U4099 ( .A1(w_q[412]), .A2(n7268), .ZN(n5187) );
NAND2_X2 U4100 ( .A1(n5189), .A2(n5190), .ZN(w_d[411]) );
NAND2_X2 U4101 ( .A1(w_q[379]), .A2(n7210), .ZN(n5190) );
NAND2_X2 U4102 ( .A1(w_q[411]), .A2(n7268), .ZN(n5189) );
NAND2_X2 U4103 ( .A1(n5191), .A2(n5192), .ZN(w_d[410]) );
NAND2_X2 U4104 ( .A1(w_q[378]), .A2(n7210), .ZN(n5192) );
NAND2_X2 U4105 ( .A1(w_q[410]), .A2(n7268), .ZN(n5191) );
NAND2_X2 U4106 ( .A1(n5193), .A2(n5194), .ZN(w_d[40]) );
NAND2_X2 U4107 ( .A1(w_q[8]), .A2(n7209), .ZN(n5194) );
NAND2_X2 U4108 ( .A1(w_q[40]), .A2(n7268), .ZN(n5193) );
NAND2_X2 U4109 ( .A1(n5195), .A2(n5196), .ZN(w_d[409]) );
NAND2_X2 U4110 ( .A1(w_q[377]), .A2(n7209), .ZN(n5196) );
NAND2_X2 U4111 ( .A1(w_q[409]), .A2(n7268), .ZN(n5195) );
NAND2_X2 U4112 ( .A1(n5197), .A2(n5198), .ZN(w_d[408]) );
NAND2_X2 U4113 ( .A1(w_q[376]), .A2(n7209), .ZN(n5198) );
NAND2_X2 U4114 ( .A1(w_q[408]), .A2(n7268), .ZN(n5197) );
NAND2_X2 U4115 ( .A1(n5199), .A2(n5200), .ZN(w_d[407]) );
NAND2_X2 U4116 ( .A1(w_q[375]), .A2(n7209), .ZN(n5200) );
NAND2_X2 U4117 ( .A1(w_q[407]), .A2(n7268), .ZN(n5199) );
NAND2_X2 U4118 ( .A1(n5201), .A2(n5202), .ZN(w_d[406]) );
NAND2_X2 U4119 ( .A1(w_q[374]), .A2(n7209), .ZN(n5202) );
NAND2_X2 U4120 ( .A1(w_q[406]), .A2(n7267), .ZN(n5201) );
NAND2_X2 U4121 ( .A1(n5203), .A2(n5204), .ZN(w_d[405]) );
NAND2_X2 U4122 ( .A1(w_q[373]), .A2(n7209), .ZN(n5204) );
NAND2_X2 U4123 ( .A1(w_q[405]), .A2(n7267), .ZN(n5203) );
NAND2_X2 U4124 ( .A1(n5205), .A2(n5206), .ZN(w_d[404]) );
NAND2_X2 U4125 ( .A1(w_q[372]), .A2(n7209), .ZN(n5206) );
NAND2_X2 U4126 ( .A1(w_q[404]), .A2(n7267), .ZN(n5205) );
NAND2_X2 U4127 ( .A1(n5207), .A2(n5208), .ZN(w_d[403]) );
NAND2_X2 U4128 ( .A1(w_q[371]), .A2(n7209), .ZN(n5208) );
NAND2_X2 U4129 ( .A1(w_q[403]), .A2(n7267), .ZN(n5207) );
NAND2_X2 U4130 ( .A1(n5209), .A2(n5210), .ZN(w_d[402]) );
NAND2_X2 U4131 ( .A1(w_q[370]), .A2(n7209), .ZN(n5210) );
NAND2_X2 U4132 ( .A1(w_q[402]), .A2(n7267), .ZN(n5209) );
NAND2_X2 U4133 ( .A1(n5211), .A2(n5212), .ZN(w_d[401]) );
NAND2_X2 U4134 ( .A1(w_q[369]), .A2(n7209), .ZN(n5212) );
NAND2_X2 U4135 ( .A1(w_q[401]), .A2(n7267), .ZN(n5211) );
NAND2_X2 U4136 ( .A1(n5213), .A2(n5214), .ZN(w_d[400]) );
NAND2_X2 U4137 ( .A1(w_q[368]), .A2(n7209), .ZN(n5214) );
NAND2_X2 U4138 ( .A1(w_q[400]), .A2(n7267), .ZN(n5213) );
NAND2_X2 U4140 ( .A1(w[3]), .A2(n7159), .ZN(n5217) );
NAND2_X2 U4141 ( .A1(w_q[3]), .A2(n7267), .ZN(n5216) );
NAND2_X2 U4143 ( .A1(n5218), .A2(n5219), .ZN(w_d[39]) );
NAND2_X2 U4144 ( .A1(w_q[7]), .A2(n7208), .ZN(n5219) );
NAND2_X2 U4145 ( .A1(w_q[39]), .A2(n7267), .ZN(n5218) );
NAND2_X2 U4146 ( .A1(n5220), .A2(n5221), .ZN(w_d[399]) );
NAND2_X2 U4147 ( .A1(w_q[367]), .A2(n7208), .ZN(n5221) );
NAND2_X2 U4148 ( .A1(w_q[399]), .A2(n7267), .ZN(n5220) );
NAND2_X2 U4149 ( .A1(n5222), .A2(n5223), .ZN(w_d[398]) );
NAND2_X2 U4150 ( .A1(w_q[366]), .A2(n7208), .ZN(n5223) );
NAND2_X2 U4151 ( .A1(w_q[398]), .A2(n7267), .ZN(n5222) );
NAND2_X2 U4152 ( .A1(n5224), .A2(n5225), .ZN(w_d[397]) );
NAND2_X2 U4153 ( .A1(w_q[365]), .A2(n7208), .ZN(n5225) );
NAND2_X2 U4154 ( .A1(w_q[397]), .A2(n7266), .ZN(n5224) );
NAND2_X2 U4155 ( .A1(n5226), .A2(n5227), .ZN(w_d[396]) );
NAND2_X2 U4156 ( .A1(w_q[364]), .A2(n7208), .ZN(n5227) );
NAND2_X2 U4157 ( .A1(w_q[396]), .A2(n7266), .ZN(n5226) );
NAND2_X2 U4158 ( .A1(n5228), .A2(n5229), .ZN(w_d[395]) );
NAND2_X2 U4159 ( .A1(w_q[363]), .A2(n7208), .ZN(n5229) );
NAND2_X2 U4160 ( .A1(w_q[395]), .A2(n7266), .ZN(n5228) );
NAND2_X2 U4161 ( .A1(n5230), .A2(n5231), .ZN(w_d[394]) );
NAND2_X2 U4162 ( .A1(w_q[362]), .A2(n7208), .ZN(n5231) );
NAND2_X2 U4163 ( .A1(w_q[394]), .A2(n7266), .ZN(n5230) );
NAND2_X2 U4164 ( .A1(n5232), .A2(n5233), .ZN(w_d[393]) );
NAND2_X2 U4165 ( .A1(w_q[361]), .A2(n7208), .ZN(n5233) );
NAND2_X2 U4166 ( .A1(w_q[393]), .A2(n7266), .ZN(n5232) );
NAND2_X2 U4167 ( .A1(n5234), .A2(n5235), .ZN(w_d[392]) );
NAND2_X2 U4168 ( .A1(w_q[360]), .A2(n7208), .ZN(n5235) );
NAND2_X2 U4169 ( .A1(w_q[392]), .A2(n7266), .ZN(n5234) );
NAND2_X2 U4170 ( .A1(n5236), .A2(n5237), .ZN(w_d[391]) );
NAND2_X2 U4171 ( .A1(w_q[359]), .A2(n7208), .ZN(n5237) );
NAND2_X2 U4172 ( .A1(w_q[391]), .A2(n7266), .ZN(n5236) );
NAND2_X2 U4173 ( .A1(n5238), .A2(n5239), .ZN(w_d[390]) );
NAND2_X2 U4174 ( .A1(w_q[358]), .A2(n7208), .ZN(n5239) );
NAND2_X2 U4175 ( .A1(w_q[390]), .A2(n7266), .ZN(n5238) );
NAND2_X2 U4176 ( .A1(n5240), .A2(n5241), .ZN(w_d[38]) );
NAND2_X2 U4177 ( .A1(w_q[6]), .A2(n7207), .ZN(n5241) );
NAND2_X2 U4178 ( .A1(w_q[38]), .A2(n7266), .ZN(n5240) );
NAND2_X2 U4179 ( .A1(n5242), .A2(n5243), .ZN(w_d[389]) );
NAND2_X2 U4180 ( .A1(w_q[357]), .A2(n7207), .ZN(n5243) );
NAND2_X2 U4181 ( .A1(w_q[389]), .A2(n7266), .ZN(n5242) );
NAND2_X2 U4182 ( .A1(n5244), .A2(n5245), .ZN(w_d[388]) );
NAND2_X2 U4183 ( .A1(w_q[356]), .A2(n7207), .ZN(n5245) );
NAND2_X2 U4184 ( .A1(w_q[388]), .A2(n7266), .ZN(n5244) );
NAND2_X2 U4185 ( .A1(n5246), .A2(n5247), .ZN(w_d[387]) );
NAND2_X2 U4186 ( .A1(w_q[355]), .A2(n7207), .ZN(n5247) );
NAND2_X2 U4187 ( .A1(w_q[387]), .A2(n7265), .ZN(n5246) );
NAND2_X2 U4188 ( .A1(n5248), .A2(n5249), .ZN(w_d[386]) );
NAND2_X2 U4189 ( .A1(w_q[354]), .A2(n7207), .ZN(n5249) );
NAND2_X2 U4190 ( .A1(w_q[386]), .A2(n7265), .ZN(n5248) );
NAND2_X2 U4191 ( .A1(n5250), .A2(n5251), .ZN(w_d[385]) );
NAND2_X2 U4192 ( .A1(w_q[353]), .A2(n7207), .ZN(n5251) );
NAND2_X2 U4193 ( .A1(w_q[385]), .A2(n7265), .ZN(n5250) );
NAND2_X2 U4194 ( .A1(n5252), .A2(n5253), .ZN(w_d[384]) );
NAND2_X2 U4195 ( .A1(w_q[352]), .A2(n7207), .ZN(n5253) );
NAND2_X2 U4196 ( .A1(w_q[384]), .A2(n7265), .ZN(n5252) );
NAND2_X2 U4197 ( .A1(n5254), .A2(n5255), .ZN(w_d[383]) );
NAND2_X2 U4198 ( .A1(w_q[351]), .A2(n7207), .ZN(n5255) );
NAND2_X2 U4199 ( .A1(w_q[383]), .A2(n7265), .ZN(n5254) );
NAND2_X2 U4200 ( .A1(n5256), .A2(n5257), .ZN(w_d[382]) );
NAND2_X2 U4201 ( .A1(w_q[350]), .A2(n7207), .ZN(n5257) );
NAND2_X2 U4202 ( .A1(w_q[382]), .A2(n7265), .ZN(n5256) );
NAND2_X2 U4203 ( .A1(n5258), .A2(n5259), .ZN(w_d[381]) );
NAND2_X2 U4204 ( .A1(w_q[349]), .A2(n7207), .ZN(n5259) );
NAND2_X2 U4205 ( .A1(w_q[381]), .A2(n7265), .ZN(n5258) );
NAND2_X2 U4206 ( .A1(n5260), .A2(n5261), .ZN(w_d[380]) );
NAND2_X2 U4207 ( .A1(w_q[348]), .A2(n7207), .ZN(n5261) );
NAND2_X2 U4208 ( .A1(w_q[380]), .A2(n7265), .ZN(n5260) );
NAND2_X2 U4209 ( .A1(n5262), .A2(n5263), .ZN(w_d[37]) );
NAND2_X2 U4210 ( .A1(w_q[5]), .A2(n7206), .ZN(n5263) );
NAND2_X2 U4211 ( .A1(w_q[37]), .A2(n7265), .ZN(n5262) );
NAND2_X2 U4212 ( .A1(n5264), .A2(n5265), .ZN(w_d[379]) );
NAND2_X2 U4213 ( .A1(w_q[347]), .A2(n7206), .ZN(n5265) );
NAND2_X2 U4214 ( .A1(w_q[379]), .A2(n7265), .ZN(n5264) );
NAND2_X2 U4215 ( .A1(n5266), .A2(n5267), .ZN(w_d[378]) );
NAND2_X2 U4216 ( .A1(w_q[346]), .A2(n7206), .ZN(n5267) );
NAND2_X2 U4217 ( .A1(w_q[378]), .A2(n7265), .ZN(n5266) );
NAND2_X2 U4218 ( .A1(n5268), .A2(n5269), .ZN(w_d[377]) );
NAND2_X2 U4219 ( .A1(w_q[345]), .A2(n7206), .ZN(n5269) );
NAND2_X2 U4220 ( .A1(w_q[377]), .A2(n7264), .ZN(n5268) );
NAND2_X2 U4221 ( .A1(n5270), .A2(n5271), .ZN(w_d[376]) );
NAND2_X2 U4222 ( .A1(w_q[344]), .A2(n7206), .ZN(n5271) );
NAND2_X2 U4223 ( .A1(w_q[376]), .A2(n7264), .ZN(n5270) );
NAND2_X2 U4224 ( .A1(n5272), .A2(n5273), .ZN(w_d[375]) );
NAND2_X2 U4225 ( .A1(w_q[343]), .A2(n7206), .ZN(n5273) );
NAND2_X2 U4226 ( .A1(w_q[375]), .A2(n7264), .ZN(n5272) );
NAND2_X2 U4227 ( .A1(n5274), .A2(n5275), .ZN(w_d[374]) );
NAND2_X2 U4228 ( .A1(w_q[342]), .A2(n7206), .ZN(n5275) );
NAND2_X2 U4229 ( .A1(w_q[374]), .A2(n7264), .ZN(n5274) );
NAND2_X2 U4230 ( .A1(n5276), .A2(n5277), .ZN(w_d[373]) );
NAND2_X2 U4231 ( .A1(w_q[341]), .A2(n7206), .ZN(n5277) );
NAND2_X2 U4232 ( .A1(w_q[373]), .A2(n7264), .ZN(n5276) );
NAND2_X2 U4233 ( .A1(n5278), .A2(n5279), .ZN(w_d[372]) );
NAND2_X2 U4234 ( .A1(w_q[340]), .A2(n7206), .ZN(n5279) );
NAND2_X2 U4235 ( .A1(w_q[372]), .A2(n7264), .ZN(n5278) );
NAND2_X2 U4236 ( .A1(n5280), .A2(n5281), .ZN(w_d[371]) );
NAND2_X2 U4237 ( .A1(w_q[339]), .A2(n7206), .ZN(n5281) );
NAND2_X2 U4238 ( .A1(w_q[371]), .A2(n7264), .ZN(n5280) );
NAND2_X2 U4239 ( .A1(n5282), .A2(n5283), .ZN(w_d[370]) );
NAND2_X2 U4240 ( .A1(w_q[338]), .A2(n7206), .ZN(n5283) );
NAND2_X2 U4241 ( .A1(w_q[370]), .A2(n7264), .ZN(n5282) );
NAND2_X2 U4242 ( .A1(n5284), .A2(n5285), .ZN(w_d[36]) );
NAND2_X2 U4243 ( .A1(w_q[4]), .A2(n7205), .ZN(n5285) );
NAND2_X2 U4244 ( .A1(w_q[36]), .A2(n7264), .ZN(n5284) );
NAND2_X2 U4245 ( .A1(n5286), .A2(n5287), .ZN(w_d[369]) );
NAND2_X2 U4246 ( .A1(w_q[337]), .A2(n7205), .ZN(n5287) );
NAND2_X2 U4247 ( .A1(w_q[369]), .A2(n7264), .ZN(n5286) );
NAND2_X2 U4248 ( .A1(n5288), .A2(n5289), .ZN(w_d[368]) );
NAND2_X2 U4249 ( .A1(w_q[336]), .A2(n7205), .ZN(n5289) );
NAND2_X2 U4250 ( .A1(w_q[368]), .A2(n7264), .ZN(n5288) );
NAND2_X2 U4251 ( .A1(n5290), .A2(n5291), .ZN(w_d[367]) );
NAND2_X2 U4252 ( .A1(w_q[335]), .A2(n7205), .ZN(n5291) );
NAND2_X2 U4253 ( .A1(w_q[367]), .A2(n7263), .ZN(n5290) );
NAND2_X2 U4254 ( .A1(n5292), .A2(n5293), .ZN(w_d[366]) );
NAND2_X2 U4255 ( .A1(w_q[334]), .A2(n7205), .ZN(n5293) );
NAND2_X2 U4256 ( .A1(w_q[366]), .A2(n7263), .ZN(n5292) );
NAND2_X2 U4257 ( .A1(n5294), .A2(n5295), .ZN(w_d[365]) );
NAND2_X2 U4258 ( .A1(w_q[333]), .A2(n7205), .ZN(n5295) );
NAND2_X2 U4259 ( .A1(w_q[365]), .A2(n7263), .ZN(n5294) );
NAND2_X2 U4260 ( .A1(n5296), .A2(n5297), .ZN(w_d[364]) );
NAND2_X2 U4261 ( .A1(w_q[332]), .A2(n7205), .ZN(n5297) );
NAND2_X2 U4262 ( .A1(w_q[364]), .A2(n7263), .ZN(n5296) );
NAND2_X2 U4263 ( .A1(n5298), .A2(n5299), .ZN(w_d[363]) );
NAND2_X2 U4264 ( .A1(w_q[331]), .A2(n7205), .ZN(n5299) );
NAND2_X2 U4265 ( .A1(w_q[363]), .A2(n7263), .ZN(n5298) );
NAND2_X2 U4266 ( .A1(n5300), .A2(n5301), .ZN(w_d[362]) );
NAND2_X2 U4267 ( .A1(w_q[330]), .A2(n7205), .ZN(n5301) );
NAND2_X2 U4268 ( .A1(w_q[362]), .A2(n7263), .ZN(n5300) );
NAND2_X2 U4269 ( .A1(n5302), .A2(n5303), .ZN(w_d[361]) );
NAND2_X2 U4270 ( .A1(w_q[329]), .A2(n7205), .ZN(n5303) );
NAND2_X2 U4271 ( .A1(w_q[361]), .A2(n7263), .ZN(n5302) );
NAND2_X2 U4272 ( .A1(n5304), .A2(n5305), .ZN(w_d[360]) );
NAND2_X2 U4273 ( .A1(w_q[328]), .A2(n7205), .ZN(n5305) );
NAND2_X2 U4274 ( .A1(w_q[360]), .A2(n7263), .ZN(n5304) );
NAND2_X2 U4275 ( .A1(n5306), .A2(n5307), .ZN(w_d[35]) );
NAND2_X2 U4276 ( .A1(w_q[3]), .A2(n7204), .ZN(n5307) );
NAND2_X2 U4277 ( .A1(w_q[35]), .A2(n7263), .ZN(n5306) );
NAND2_X2 U4278 ( .A1(n5308), .A2(n5309), .ZN(w_d[359]) );
NAND2_X2 U4279 ( .A1(w_q[327]), .A2(n7204), .ZN(n5309) );
NAND2_X2 U4280 ( .A1(w_q[359]), .A2(n7263), .ZN(n5308) );
NAND2_X2 U4281 ( .A1(n5310), .A2(n5311), .ZN(w_d[358]) );
NAND2_X2 U4282 ( .A1(w_q[326]), .A2(n7204), .ZN(n5311) );
NAND2_X2 U4283 ( .A1(w_q[358]), .A2(n7263), .ZN(n5310) );
NAND2_X2 U4284 ( .A1(n5312), .A2(n5313), .ZN(w_d[357]) );
NAND2_X2 U4285 ( .A1(w_q[325]), .A2(n7204), .ZN(n5313) );
NAND2_X2 U4286 ( .A1(w_q[357]), .A2(n7262), .ZN(n5312) );
NAND2_X2 U4287 ( .A1(n5314), .A2(n5315), .ZN(w_d[356]) );
NAND2_X2 U4288 ( .A1(w_q[324]), .A2(n7204), .ZN(n5315) );
NAND2_X2 U4289 ( .A1(w_q[356]), .A2(n7262), .ZN(n5314) );
NAND2_X2 U4290 ( .A1(n5316), .A2(n5317), .ZN(w_d[355]) );
NAND2_X2 U4291 ( .A1(w_q[323]), .A2(n7204), .ZN(n5317) );
NAND2_X2 U4292 ( .A1(w_q[355]), .A2(n7262), .ZN(n5316) );
NAND2_X2 U4293 ( .A1(n5318), .A2(n5319), .ZN(w_d[354]) );
NAND2_X2 U4294 ( .A1(w_q[322]), .A2(n7204), .ZN(n5319) );
NAND2_X2 U4295 ( .A1(w_q[354]), .A2(n7262), .ZN(n5318) );
NAND2_X2 U4296 ( .A1(n5320), .A2(n5321), .ZN(w_d[353]) );
NAND2_X2 U4297 ( .A1(w_q[321]), .A2(n7204), .ZN(n5321) );
NAND2_X2 U4298 ( .A1(w_q[353]), .A2(n7262), .ZN(n5320) );
NAND2_X2 U4299 ( .A1(n5322), .A2(n5323), .ZN(w_d[352]) );
NAND2_X2 U4300 ( .A1(w_q[320]), .A2(n7204), .ZN(n5323) );
NAND2_X2 U4301 ( .A1(w_q[352]), .A2(n7262), .ZN(n5322) );
NAND2_X2 U4302 ( .A1(n5324), .A2(n5325), .ZN(w_d[351]) );
NAND2_X2 U4303 ( .A1(w_q[319]), .A2(n7204), .ZN(n5325) );
NAND2_X2 U4304 ( .A1(w_q[351]), .A2(n7262), .ZN(n5324) );
NAND2_X2 U4305 ( .A1(n5326), .A2(n5327), .ZN(w_d[350]) );
NAND2_X2 U4306 ( .A1(w_q[318]), .A2(n7204), .ZN(n5327) );
NAND2_X2 U4307 ( .A1(w_q[350]), .A2(n7262), .ZN(n5326) );
NAND2_X2 U4308 ( .A1(n5328), .A2(n5329), .ZN(w_d[34]) );
NAND2_X2 U4309 ( .A1(w_q[2]), .A2(n7203), .ZN(n5329) );
NAND2_X2 U4310 ( .A1(w_q[34]), .A2(n7262), .ZN(n5328) );
NAND2_X2 U4311 ( .A1(n5330), .A2(n5331), .ZN(w_d[349]) );
NAND2_X2 U4312 ( .A1(w_q[317]), .A2(n7203), .ZN(n5331) );
NAND2_X2 U4313 ( .A1(w_q[349]), .A2(n7262), .ZN(n5330) );
NAND2_X2 U4314 ( .A1(n5332), .A2(n5333), .ZN(w_d[348]) );
NAND2_X2 U4315 ( .A1(w_q[316]), .A2(n7203), .ZN(n5333) );
NAND2_X2 U4316 ( .A1(w_q[348]), .A2(n7262), .ZN(n5332) );
NAND2_X2 U4317 ( .A1(n5334), .A2(n5335), .ZN(w_d[347]) );
NAND2_X2 U4318 ( .A1(w_q[315]), .A2(n7203), .ZN(n5335) );
NAND2_X2 U4319 ( .A1(w_q[347]), .A2(n7261), .ZN(n5334) );
NAND2_X2 U4320 ( .A1(n5336), .A2(n5337), .ZN(w_d[346]) );
NAND2_X2 U4321 ( .A1(w_q[314]), .A2(n7203), .ZN(n5337) );
NAND2_X2 U4322 ( .A1(w_q[346]), .A2(n7261), .ZN(n5336) );
NAND2_X2 U4323 ( .A1(n5338), .A2(n5339), .ZN(w_d[345]) );
NAND2_X2 U4324 ( .A1(w_q[313]), .A2(n7203), .ZN(n5339) );
NAND2_X2 U4325 ( .A1(w_q[345]), .A2(n7261), .ZN(n5338) );
NAND2_X2 U4326 ( .A1(n5340), .A2(n5341), .ZN(w_d[344]) );
NAND2_X2 U4327 ( .A1(w_q[312]), .A2(n7203), .ZN(n5341) );
NAND2_X2 U4328 ( .A1(w_q[344]), .A2(n7261), .ZN(n5340) );
NAND2_X2 U4329 ( .A1(n5342), .A2(n5343), .ZN(w_d[343]) );
NAND2_X2 U4330 ( .A1(w_q[311]), .A2(n7203), .ZN(n5343) );
NAND2_X2 U4331 ( .A1(w_q[343]), .A2(n7261), .ZN(n5342) );
NAND2_X2 U4332 ( .A1(n5344), .A2(n5345), .ZN(w_d[342]) );
NAND2_X2 U4333 ( .A1(w_q[310]), .A2(n7203), .ZN(n5345) );
NAND2_X2 U4334 ( .A1(w_q[342]), .A2(n7261), .ZN(n5344) );
NAND2_X2 U4335 ( .A1(n5346), .A2(n5347), .ZN(w_d[341]) );
NAND2_X2 U4336 ( .A1(w_q[309]), .A2(n7203), .ZN(n5347) );
NAND2_X2 U4337 ( .A1(w_q[341]), .A2(n7261), .ZN(n5346) );
NAND2_X2 U4338 ( .A1(n5348), .A2(n5349), .ZN(w_d[340]) );
NAND2_X2 U4339 ( .A1(w_q[308]), .A2(n7203), .ZN(n5349) );
NAND2_X2 U4340 ( .A1(w_q[340]), .A2(n7261), .ZN(n5348) );
NAND2_X2 U4341 ( .A1(n5350), .A2(n5351), .ZN(w_d[33]) );
NAND2_X2 U4342 ( .A1(w_q[1]), .A2(n7202), .ZN(n5351) );
NAND2_X2 U4343 ( .A1(w_q[33]), .A2(n7261), .ZN(n5350) );
NAND2_X2 U4344 ( .A1(n5352), .A2(n5353), .ZN(w_d[339]) );
NAND2_X2 U4345 ( .A1(w_q[307]), .A2(n7202), .ZN(n5353) );
NAND2_X2 U4346 ( .A1(w_q[339]), .A2(n7261), .ZN(n5352) );
NAND2_X2 U4347 ( .A1(n5354), .A2(n5355), .ZN(w_d[338]) );
NAND2_X2 U4348 ( .A1(w_q[306]), .A2(n7202), .ZN(n5355) );
NAND2_X2 U4349 ( .A1(w_q[338]), .A2(n7261), .ZN(n5354) );
NAND2_X2 U4350 ( .A1(n5356), .A2(n5357), .ZN(w_d[337]) );
NAND2_X2 U4351 ( .A1(w_q[305]), .A2(n7202), .ZN(n5357) );
NAND2_X2 U4352 ( .A1(w_q[337]), .A2(n7260), .ZN(n5356) );
NAND2_X2 U4353 ( .A1(n5358), .A2(n5359), .ZN(w_d[336]) );
NAND2_X2 U4354 ( .A1(w_q[304]), .A2(n7202), .ZN(n5359) );
NAND2_X2 U4355 ( .A1(w_q[336]), .A2(n7260), .ZN(n5358) );
NAND2_X2 U4356 ( .A1(n5360), .A2(n5361), .ZN(w_d[335]) );
NAND2_X2 U4357 ( .A1(w_q[303]), .A2(n7202), .ZN(n5361) );
NAND2_X2 U4358 ( .A1(w_q[335]), .A2(n7260), .ZN(n5360) );
NAND2_X2 U4359 ( .A1(n5362), .A2(n5363), .ZN(w_d[334]) );
NAND2_X2 U4360 ( .A1(w_q[302]), .A2(n7202), .ZN(n5363) );
NAND2_X2 U4361 ( .A1(w_q[334]), .A2(n7260), .ZN(n5362) );
NAND2_X2 U4362 ( .A1(n5364), .A2(n5365), .ZN(w_d[333]) );
NAND2_X2 U4363 ( .A1(w_q[301]), .A2(n7202), .ZN(n5365) );
NAND2_X2 U4364 ( .A1(w_q[333]), .A2(n7260), .ZN(n5364) );
NAND2_X2 U4365 ( .A1(n5366), .A2(n5367), .ZN(w_d[332]) );
NAND2_X2 U4366 ( .A1(w_q[300]), .A2(n7202), .ZN(n5367) );
NAND2_X2 U4367 ( .A1(w_q[332]), .A2(n7260), .ZN(n5366) );
NAND2_X2 U4368 ( .A1(n5368), .A2(n5369), .ZN(w_d[331]) );
NAND2_X2 U4369 ( .A1(w_q[299]), .A2(n7202), .ZN(n5369) );
NAND2_X2 U4370 ( .A1(w_q[331]), .A2(n7260), .ZN(n5368) );
NAND2_X2 U4371 ( .A1(n5370), .A2(n5371), .ZN(w_d[330]) );
NAND2_X2 U4372 ( .A1(w_q[298]), .A2(n7202), .ZN(n5371) );
NAND2_X2 U4373 ( .A1(w_q[330]), .A2(n7260), .ZN(n5370) );
NAND2_X2 U4374 ( .A1(n5372), .A2(n5373), .ZN(w_d[32]) );
NAND2_X2 U4375 ( .A1(w_q[0]), .A2(n7201), .ZN(n5373) );
NAND2_X2 U4376 ( .A1(w_q[32]), .A2(n7260), .ZN(n5372) );
NAND2_X2 U4377 ( .A1(n5374), .A2(n5375), .ZN(w_d[329]) );
NAND2_X2 U4378 ( .A1(w_q[297]), .A2(n7201), .ZN(n5375) );
NAND2_X2 U4379 ( .A1(w_q[329]), .A2(n7260), .ZN(n5374) );
NAND2_X2 U4380 ( .A1(n5376), .A2(n5377), .ZN(w_d[328]) );
NAND2_X2 U4381 ( .A1(w_q[296]), .A2(n7201), .ZN(n5377) );
NAND2_X2 U4382 ( .A1(w_q[328]), .A2(n7260), .ZN(n5376) );
NAND2_X2 U4383 ( .A1(n5378), .A2(n5379), .ZN(w_d[327]) );
NAND2_X2 U4384 ( .A1(w_q[295]), .A2(n7201), .ZN(n5379) );
NAND2_X2 U4385 ( .A1(w_q[327]), .A2(n7259), .ZN(n5378) );
NAND2_X2 U4386 ( .A1(n5380), .A2(n5381), .ZN(w_d[326]) );
NAND2_X2 U4387 ( .A1(w_q[294]), .A2(n7201), .ZN(n5381) );
NAND2_X2 U4388 ( .A1(w_q[326]), .A2(n7259), .ZN(n5380) );
NAND2_X2 U4389 ( .A1(n5382), .A2(n5383), .ZN(w_d[325]) );
NAND2_X2 U4390 ( .A1(w_q[293]), .A2(n7201), .ZN(n5383) );
NAND2_X2 U4391 ( .A1(w_q[325]), .A2(n7259), .ZN(n5382) );
NAND2_X2 U4392 ( .A1(n5384), .A2(n5385), .ZN(w_d[324]) );
NAND2_X2 U4393 ( .A1(w_q[292]), .A2(n7201), .ZN(n5385) );
NAND2_X2 U4394 ( .A1(w_q[324]), .A2(n7259), .ZN(n5384) );
NAND2_X2 U4395 ( .A1(n5386), .A2(n5387), .ZN(w_d[323]) );
NAND2_X2 U4396 ( .A1(w_q[291]), .A2(n7201), .ZN(n5387) );
NAND2_X2 U4397 ( .A1(w_q[323]), .A2(n7259), .ZN(n5386) );
NAND2_X2 U4398 ( .A1(n5388), .A2(n5389), .ZN(w_d[322]) );
NAND2_X2 U4399 ( .A1(w_q[290]), .A2(n7201), .ZN(n5389) );
NAND2_X2 U4400 ( .A1(w_q[322]), .A2(n7259), .ZN(n5388) );
NAND2_X2 U4401 ( .A1(n5390), .A2(n5391), .ZN(w_d[321]) );
NAND2_X2 U4402 ( .A1(w_q[289]), .A2(n7201), .ZN(n5391) );
NAND2_X2 U4403 ( .A1(w_q[321]), .A2(n7259), .ZN(n5390) );
NAND2_X2 U4404 ( .A1(n5392), .A2(n5393), .ZN(w_d[320]) );
NAND2_X2 U4405 ( .A1(w_q[288]), .A2(n7201), .ZN(n5393) );
NAND2_X2 U4406 ( .A1(w_q[320]), .A2(n7259), .ZN(n5392) );
NAND2_X2 U4408 ( .A1(w[31]), .A2(n7159), .ZN(n5396) );
NAND2_X2 U4409 ( .A1(w_q[31]), .A2(n7259), .ZN(n5395) );
NAND2_X2 U4411 ( .A1(n5397), .A2(n5398), .ZN(w_d[319]) );
NAND2_X2 U4412 ( .A1(w_q[287]), .A2(n7200), .ZN(n5398) );
NAND2_X2 U4413 ( .A1(w_q[319]), .A2(n7259), .ZN(n5397) );
NAND2_X2 U4414 ( .A1(n5399), .A2(n5400), .ZN(w_d[318]) );
NAND2_X2 U4415 ( .A1(w_q[286]), .A2(n7200), .ZN(n5400) );
NAND2_X2 U4416 ( .A1(w_q[318]), .A2(n7259), .ZN(n5399) );
NAND2_X2 U4417 ( .A1(n5401), .A2(n5402), .ZN(w_d[317]) );
NAND2_X2 U4418 ( .A1(w_q[285]), .A2(n7200), .ZN(n5402) );
NAND2_X2 U4419 ( .A1(w_q[317]), .A2(n7258), .ZN(n5401) );
NAND2_X2 U4420 ( .A1(n5403), .A2(n5404), .ZN(w_d[316]) );
NAND2_X2 U4421 ( .A1(w_q[284]), .A2(n7200), .ZN(n5404) );
NAND2_X2 U4422 ( .A1(w_q[316]), .A2(n7258), .ZN(n5403) );
NAND2_X2 U4423 ( .A1(n5405), .A2(n5406), .ZN(w_d[315]) );
NAND2_X2 U4424 ( .A1(w_q[283]), .A2(n7200), .ZN(n5406) );
NAND2_X2 U4425 ( .A1(w_q[315]), .A2(n7258), .ZN(n5405) );
NAND2_X2 U4426 ( .A1(n5407), .A2(n5408), .ZN(w_d[314]) );
NAND2_X2 U4427 ( .A1(w_q[282]), .A2(n7200), .ZN(n5408) );
NAND2_X2 U4428 ( .A1(w_q[314]), .A2(n7258), .ZN(n5407) );
NAND2_X2 U4429 ( .A1(n5409), .A2(n5410), .ZN(w_d[313]) );
NAND2_X2 U4430 ( .A1(w_q[281]), .A2(n7200), .ZN(n5410) );
NAND2_X2 U4431 ( .A1(w_q[313]), .A2(n7258), .ZN(n5409) );
NAND2_X2 U4432 ( .A1(n5411), .A2(n5412), .ZN(w_d[312]) );
NAND2_X2 U4433 ( .A1(w_q[280]), .A2(n7200), .ZN(n5412) );
NAND2_X2 U4434 ( .A1(w_q[312]), .A2(n7258), .ZN(n5411) );
NAND2_X2 U4435 ( .A1(n5413), .A2(n5414), .ZN(w_d[311]) );
NAND2_X2 U4436 ( .A1(w_q[279]), .A2(n7200), .ZN(n5414) );
NAND2_X2 U4437 ( .A1(w_q[311]), .A2(n7258), .ZN(n5413) );
NAND2_X2 U4438 ( .A1(n5415), .A2(n5416), .ZN(w_d[310]) );
NAND2_X2 U4439 ( .A1(w_q[278]), .A2(n7200), .ZN(n5416) );
NAND2_X2 U4440 ( .A1(w_q[310]), .A2(n7258), .ZN(n5415) );
NAND2_X2 U4442 ( .A1(w[30]), .A2(n7159), .ZN(n5419) );
NAND2_X2 U4443 ( .A1(w_q[30]), .A2(n7258), .ZN(n5418) );
NAND2_X2 U4445 ( .A1(n5420), .A2(n5421), .ZN(w_d[309]) );
NAND2_X2 U4446 ( .A1(w_q[277]), .A2(n7200), .ZN(n5421) );
NAND2_X2 U4447 ( .A1(w_q[309]), .A2(n7258), .ZN(n5420) );
NAND2_X2 U4448 ( .A1(n5422), .A2(n5423), .ZN(w_d[308]) );
NAND2_X2 U4449 ( .A1(w_q[276]), .A2(n7199), .ZN(n5423) );
NAND2_X2 U4450 ( .A1(w_q[308]), .A2(n7258), .ZN(n5422) );
NAND2_X2 U4451 ( .A1(n5424), .A2(n5425), .ZN(w_d[307]) );
NAND2_X2 U4452 ( .A1(w_q[275]), .A2(n7199), .ZN(n5425) );
NAND2_X2 U4453 ( .A1(w_q[307]), .A2(n7257), .ZN(n5424) );
NAND2_X2 U4454 ( .A1(n5426), .A2(n5427), .ZN(w_d[306]) );
NAND2_X2 U4455 ( .A1(w_q[274]), .A2(n7199), .ZN(n5427) );
NAND2_X2 U4456 ( .A1(w_q[306]), .A2(n7257), .ZN(n5426) );
NAND2_X2 U4457 ( .A1(n5428), .A2(n5429), .ZN(w_d[305]) );
NAND2_X2 U4458 ( .A1(w_q[273]), .A2(n7199), .ZN(n5429) );
NAND2_X2 U4459 ( .A1(w_q[305]), .A2(n7257), .ZN(n5428) );
NAND2_X2 U4460 ( .A1(n5430), .A2(n5431), .ZN(w_d[304]) );
NAND2_X2 U4461 ( .A1(w_q[272]), .A2(n7199), .ZN(n5431) );
NAND2_X2 U4462 ( .A1(w_q[304]), .A2(n7257), .ZN(n5430) );
NAND2_X2 U4463 ( .A1(n5432), .A2(n5433), .ZN(w_d[303]) );
NAND2_X2 U4464 ( .A1(w_q[271]), .A2(n7199), .ZN(n5433) );
NAND2_X2 U4465 ( .A1(w_q[303]), .A2(n7257), .ZN(n5432) );
NAND2_X2 U4466 ( .A1(n5434), .A2(n5435), .ZN(w_d[302]) );
NAND2_X2 U4467 ( .A1(w_q[270]), .A2(n7199), .ZN(n5435) );
NAND2_X2 U4468 ( .A1(w_q[302]), .A2(n7257), .ZN(n5434) );
NAND2_X2 U4469 ( .A1(n5436), .A2(n5437), .ZN(w_d[301]) );
NAND2_X2 U4470 ( .A1(w_q[269]), .A2(n7199), .ZN(n5437) );
NAND2_X2 U4471 ( .A1(w_q[301]), .A2(n7257), .ZN(n5436) );
NAND2_X2 U4472 ( .A1(n5438), .A2(n5439), .ZN(w_d[300]) );
NAND2_X2 U4473 ( .A1(w_q[268]), .A2(n7199), .ZN(n5439) );
NAND2_X2 U4474 ( .A1(w_q[300]), .A2(n7257), .ZN(n5438) );
NAND2_X2 U4476 ( .A1(w[2]), .A2(n7159), .ZN(n5442) );
NAND2_X2 U4477 ( .A1(w_q[2]), .A2(n7257), .ZN(n5441) );
NAND2_X2 U4480 ( .A1(w[29]), .A2(n7159), .ZN(n5445) );
NAND2_X2 U4481 ( .A1(w_q[29]), .A2(n7257), .ZN(n5444) );
NAND2_X2 U4483 ( .A1(n5446), .A2(n5447), .ZN(w_d[299]) );
NAND2_X2 U4484 ( .A1(w_q[267]), .A2(n7199), .ZN(n5447) );
NAND2_X2 U4485 ( .A1(w_q[299]), .A2(n7257), .ZN(n5446) );
NAND2_X2 U4486 ( .A1(n5448), .A2(n5449), .ZN(w_d[298]) );
NAND2_X2 U4487 ( .A1(w_q[266]), .A2(n7199), .ZN(n5449) );
NAND2_X2 U4488 ( .A1(w_q[298]), .A2(n7256), .ZN(n5448) );
NAND2_X2 U4489 ( .A1(n5450), .A2(n5451), .ZN(w_d[297]) );
NAND2_X2 U4490 ( .A1(w_q[265]), .A2(n7198), .ZN(n5451) );
NAND2_X2 U4491 ( .A1(w_q[297]), .A2(n7256), .ZN(n5450) );
NAND2_X2 U4492 ( .A1(n5452), .A2(n5453), .ZN(w_d[296]) );
NAND2_X2 U4493 ( .A1(w_q[264]), .A2(n7198), .ZN(n5453) );
NAND2_X2 U4494 ( .A1(w_q[296]), .A2(n7256), .ZN(n5452) );
NAND2_X2 U4495 ( .A1(n5454), .A2(n5455), .ZN(w_d[295]) );
NAND2_X2 U4496 ( .A1(w_q[263]), .A2(n7198), .ZN(n5455) );
NAND2_X2 U4497 ( .A1(w_q[295]), .A2(n7256), .ZN(n5454) );
NAND2_X2 U4498 ( .A1(n5456), .A2(n5457), .ZN(w_d[294]) );
NAND2_X2 U4499 ( .A1(w_q[262]), .A2(n7198), .ZN(n5457) );
NAND2_X2 U4500 ( .A1(w_q[294]), .A2(n7256), .ZN(n5456) );
NAND2_X2 U4501 ( .A1(n5458), .A2(n5459), .ZN(w_d[293]) );
NAND2_X2 U4502 ( .A1(w_q[261]), .A2(n7198), .ZN(n5459) );
NAND2_X2 U4503 ( .A1(w_q[293]), .A2(n7256), .ZN(n5458) );
NAND2_X2 U4504 ( .A1(n5460), .A2(n5461), .ZN(w_d[292]) );
NAND2_X2 U4505 ( .A1(w_q[260]), .A2(n7198), .ZN(n5461) );
NAND2_X2 U4506 ( .A1(w_q[292]), .A2(n7256), .ZN(n5460) );
NAND2_X2 U4507 ( .A1(n5462), .A2(n5463), .ZN(w_d[291]) );
NAND2_X2 U4508 ( .A1(w_q[259]), .A2(n7198), .ZN(n5463) );
NAND2_X2 U4509 ( .A1(w_q[291]), .A2(n7256), .ZN(n5462) );
NAND2_X2 U4510 ( .A1(n5464), .A2(n5465), .ZN(w_d[290]) );
NAND2_X2 U4511 ( .A1(w_q[258]), .A2(n7198), .ZN(n5465) );
NAND2_X2 U4512 ( .A1(w_q[290]), .A2(n7256), .ZN(n5464) );
NAND2_X2 U4514 ( .A1(w[28]), .A2(n7159), .ZN(n5468) );
NAND2_X2 U4515 ( .A1(w_q[28]), .A2(n7256), .ZN(n5467) );
NAND2_X2 U4517 ( .A1(n5469), .A2(n5470), .ZN(w_d[289]) );
NAND2_X2 U4518 ( .A1(w_q[257]), .A2(n7198), .ZN(n5470) );
NAND2_X2 U4519 ( .A1(w_q[289]), .A2(n7256), .ZN(n5469) );
NAND2_X2 U4520 ( .A1(n5471), .A2(n5472), .ZN(w_d[288]) );
NAND2_X2 U4521 ( .A1(w_q[256]), .A2(n7198), .ZN(n5472) );
NAND2_X2 U4522 ( .A1(w_q[288]), .A2(n7255), .ZN(n5471) );
NAND2_X2 U4523 ( .A1(n5473), .A2(n5474), .ZN(w_d[287]) );
NAND2_X2 U4524 ( .A1(w_q[255]), .A2(n7198), .ZN(n5474) );
NAND2_X2 U4525 ( .A1(w_q[287]), .A2(n7255), .ZN(n5473) );
NAND2_X2 U4526 ( .A1(n5475), .A2(n5476), .ZN(w_d[286]) );
NAND2_X2 U4527 ( .A1(w_q[254]), .A2(n7197), .ZN(n5476) );
NAND2_X2 U4528 ( .A1(w_q[286]), .A2(n7255), .ZN(n5475) );
NAND2_X2 U4529 ( .A1(n5477), .A2(n5478), .ZN(w_d[285]) );
NAND2_X2 U4530 ( .A1(w_q[253]), .A2(n7197), .ZN(n5478) );
NAND2_X2 U4531 ( .A1(w_q[285]), .A2(n7255), .ZN(n5477) );
NAND2_X2 U4532 ( .A1(n5479), .A2(n5480), .ZN(w_d[284]) );
NAND2_X2 U4533 ( .A1(w_q[252]), .A2(n7197), .ZN(n5480) );
NAND2_X2 U4534 ( .A1(w_q[284]), .A2(n7255), .ZN(n5479) );
NAND2_X2 U4535 ( .A1(n5481), .A2(n5482), .ZN(w_d[283]) );
NAND2_X2 U4536 ( .A1(w_q[251]), .A2(n7197), .ZN(n5482) );
NAND2_X2 U4537 ( .A1(w_q[283]), .A2(n7255), .ZN(n5481) );
NAND2_X2 U4538 ( .A1(n5483), .A2(n5484), .ZN(w_d[282]) );
NAND2_X2 U4539 ( .A1(w_q[250]), .A2(n7197), .ZN(n5484) );
NAND2_X2 U4540 ( .A1(w_q[282]), .A2(n7255), .ZN(n5483) );
NAND2_X2 U4541 ( .A1(n5485), .A2(n5486), .ZN(w_d[281]) );
NAND2_X2 U4542 ( .A1(w_q[249]), .A2(n7197), .ZN(n5486) );
NAND2_X2 U4543 ( .A1(w_q[281]), .A2(n7255), .ZN(n5485) );
NAND2_X2 U4544 ( .A1(n5487), .A2(n5488), .ZN(w_d[280]) );
NAND2_X2 U4545 ( .A1(w_q[248]), .A2(n7197), .ZN(n5488) );
NAND2_X2 U4546 ( .A1(w_q[280]), .A2(n7255), .ZN(n5487) );
NAND2_X2 U4548 ( .A1(w[27]), .A2(n7159), .ZN(n5491) );
NAND2_X2 U4549 ( .A1(w_q[27]), .A2(n7255), .ZN(n5490) );
NAND2_X2 U4551 ( .A1(n5492), .A2(n5493), .ZN(w_d[279]) );
NAND2_X2 U4552 ( .A1(w_q[247]), .A2(n7197), .ZN(n5493) );
NAND2_X2 U4553 ( .A1(w_q[279]), .A2(n7255), .ZN(n5492) );
NAND2_X2 U4554 ( .A1(n5494), .A2(n5495), .ZN(w_d[278]) );
NAND2_X2 U4555 ( .A1(w_q[246]), .A2(n7197), .ZN(n5495) );
NAND2_X2 U4556 ( .A1(w_q[278]), .A2(n7254), .ZN(n5494) );
NAND2_X2 U4557 ( .A1(n5496), .A2(n5497), .ZN(w_d[277]) );
NAND2_X2 U4558 ( .A1(w_q[245]), .A2(n7197), .ZN(n5497) );
NAND2_X2 U4559 ( .A1(w_q[277]), .A2(n7254), .ZN(n5496) );
NAND2_X2 U4560 ( .A1(n5498), .A2(n5499), .ZN(w_d[276]) );
NAND2_X2 U4561 ( .A1(w_q[244]), .A2(n7197), .ZN(n5499) );
NAND2_X2 U4562 ( .A1(w_q[276]), .A2(n7254), .ZN(n5498) );
NAND2_X2 U4563 ( .A1(n5500), .A2(n5501), .ZN(w_d[275]) );
NAND2_X2 U4564 ( .A1(w_q[243]), .A2(n7196), .ZN(n5501) );
NAND2_X2 U4565 ( .A1(w_q[275]), .A2(n7254), .ZN(n5500) );
NAND2_X2 U4566 ( .A1(n5502), .A2(n5503), .ZN(w_d[274]) );
NAND2_X2 U4567 ( .A1(w_q[242]), .A2(n7196), .ZN(n5503) );
NAND2_X2 U4568 ( .A1(w_q[274]), .A2(n7254), .ZN(n5502) );
NAND2_X2 U4569 ( .A1(n5504), .A2(n5505), .ZN(w_d[273]) );
NAND2_X2 U4570 ( .A1(w_q[241]), .A2(n7196), .ZN(n5505) );
NAND2_X2 U4571 ( .A1(w_q[273]), .A2(n7254), .ZN(n5504) );
NAND2_X2 U4572 ( .A1(n5506), .A2(n5507), .ZN(w_d[272]) );
NAND2_X2 U4573 ( .A1(w_q[240]), .A2(n7196), .ZN(n5507) );
NAND2_X2 U4574 ( .A1(w_q[272]), .A2(n7254), .ZN(n5506) );
NAND2_X2 U4575 ( .A1(n5508), .A2(n5509), .ZN(w_d[271]) );
NAND2_X2 U4576 ( .A1(w_q[239]), .A2(n7196), .ZN(n5509) );
NAND2_X2 U4577 ( .A1(w_q[271]), .A2(n7254), .ZN(n5508) );
NAND2_X2 U4578 ( .A1(n5510), .A2(n5511), .ZN(w_d[270]) );
NAND2_X2 U4579 ( .A1(w_q[238]), .A2(n7196), .ZN(n5511) );
NAND2_X2 U4580 ( .A1(w_q[270]), .A2(n7254), .ZN(n5510) );
NAND2_X2 U4582 ( .A1(w[26]), .A2(n7160), .ZN(n5514) );
NAND2_X2 U4583 ( .A1(w_q[26]), .A2(n7254), .ZN(n5513) );
NAND2_X2 U4585 ( .A1(n5515), .A2(n5516), .ZN(w_d[269]) );
NAND2_X2 U4586 ( .A1(w_q[237]), .A2(n7196), .ZN(n5516) );
NAND2_X2 U4587 ( .A1(w_q[269]), .A2(n7254), .ZN(n5515) );
NAND2_X2 U4588 ( .A1(n5517), .A2(n5518), .ZN(w_d[268]) );
NAND2_X2 U4589 ( .A1(w_q[236]), .A2(n7196), .ZN(n5518) );
NAND2_X2 U4590 ( .A1(w_q[268]), .A2(n7253), .ZN(n5517) );
NAND2_X2 U4591 ( .A1(n5519), .A2(n5520), .ZN(w_d[267]) );
NAND2_X2 U4592 ( .A1(w_q[235]), .A2(n7196), .ZN(n5520) );
NAND2_X2 U4593 ( .A1(w_q[267]), .A2(n7253), .ZN(n5519) );
NAND2_X2 U4594 ( .A1(n5521), .A2(n5522), .ZN(w_d[266]) );
NAND2_X2 U4595 ( .A1(w_q[234]), .A2(n7196), .ZN(n5522) );
NAND2_X2 U4596 ( .A1(w_q[266]), .A2(n7253), .ZN(n5521) );
NAND2_X2 U4597 ( .A1(n5523), .A2(n5524), .ZN(w_d[265]) );
NAND2_X2 U4598 ( .A1(w_q[233]), .A2(n7196), .ZN(n5524) );
NAND2_X2 U4599 ( .A1(w_q[265]), .A2(n7253), .ZN(n5523) );
NAND2_X2 U4600 ( .A1(n5525), .A2(n5526), .ZN(w_d[264]) );
NAND2_X2 U4601 ( .A1(w_q[232]), .A2(n7195), .ZN(n5526) );
NAND2_X2 U4602 ( .A1(w_q[264]), .A2(n7253), .ZN(n5525) );
NAND2_X2 U4603 ( .A1(n5527), .A2(n5528), .ZN(w_d[263]) );
NAND2_X2 U4604 ( .A1(w_q[231]), .A2(n7195), .ZN(n5528) );
NAND2_X2 U4605 ( .A1(w_q[263]), .A2(n7253), .ZN(n5527) );
NAND2_X2 U4606 ( .A1(n5529), .A2(n5530), .ZN(w_d[262]) );
NAND2_X2 U4607 ( .A1(w_q[230]), .A2(n7195), .ZN(n5530) );
NAND2_X2 U4608 ( .A1(w_q[262]), .A2(n7253), .ZN(n5529) );
NAND2_X2 U4609 ( .A1(n5531), .A2(n5532), .ZN(w_d[261]) );
NAND2_X2 U4610 ( .A1(w_q[229]), .A2(n7195), .ZN(n5532) );
NAND2_X2 U4611 ( .A1(w_q[261]), .A2(n7253), .ZN(n5531) );
NAND2_X2 U4612 ( .A1(n5533), .A2(n5534), .ZN(w_d[260]) );
NAND2_X2 U4613 ( .A1(w_q[228]), .A2(n7195), .ZN(n5534) );
NAND2_X2 U4614 ( .A1(w_q[260]), .A2(n7253), .ZN(n5533) );
NAND2_X2 U4616 ( .A1(w[25]), .A2(n7160), .ZN(n5537) );
NAND2_X2 U4617 ( .A1(w_q[25]), .A2(n7253), .ZN(n5536) );
NAND2_X2 U4619 ( .A1(n5538), .A2(n5539), .ZN(w_d[259]) );
NAND2_X2 U4620 ( .A1(w_q[227]), .A2(n7195), .ZN(n5539) );
NAND2_X2 U4621 ( .A1(w_q[259]), .A2(n7253), .ZN(n5538) );
NAND2_X2 U4622 ( .A1(n5540), .A2(n5541), .ZN(w_d[258]) );
NAND2_X2 U4623 ( .A1(w_q[226]), .A2(n7195), .ZN(n5541) );
NAND2_X2 U4624 ( .A1(w_q[258]), .A2(n7252), .ZN(n5540) );
NAND2_X2 U4625 ( .A1(n5542), .A2(n5543), .ZN(w_d[257]) );
NAND2_X2 U4626 ( .A1(w_q[225]), .A2(n7195), .ZN(n5543) );
NAND2_X2 U4627 ( .A1(w_q[257]), .A2(n7252), .ZN(n5542) );
NAND2_X2 U4628 ( .A1(n5544), .A2(n5545), .ZN(w_d[256]) );
NAND2_X2 U4629 ( .A1(w_q[224]), .A2(n7195), .ZN(n5545) );
NAND2_X2 U4630 ( .A1(w_q[256]), .A2(n7252), .ZN(n5544) );
NAND2_X2 U4631 ( .A1(n5546), .A2(n5547), .ZN(w_d[255]) );
NAND2_X2 U4632 ( .A1(w_q[223]), .A2(n7195), .ZN(n5547) );
NAND2_X2 U4633 ( .A1(w_q[255]), .A2(n7252), .ZN(n5546) );
NAND2_X2 U4634 ( .A1(n5548), .A2(n5549), .ZN(w_d[254]) );
NAND2_X2 U4635 ( .A1(w_q[222]), .A2(n7195), .ZN(n5549) );
NAND2_X2 U4636 ( .A1(w_q[254]), .A2(n7252), .ZN(n5548) );
NAND2_X2 U4637 ( .A1(n5550), .A2(n5551), .ZN(w_d[253]) );
NAND2_X2 U4638 ( .A1(w_q[221]), .A2(n7194), .ZN(n5551) );
NAND2_X2 U4639 ( .A1(w_q[253]), .A2(n7252), .ZN(n5550) );
NAND2_X2 U4640 ( .A1(n5552), .A2(n5553), .ZN(w_d[252]) );
NAND2_X2 U4641 ( .A1(w_q[220]), .A2(n7194), .ZN(n5553) );
NAND2_X2 U4642 ( .A1(w_q[252]), .A2(n7252), .ZN(n5552) );
NAND2_X2 U4643 ( .A1(n5554), .A2(n5555), .ZN(w_d[251]) );
NAND2_X2 U4644 ( .A1(w_q[219]), .A2(n7194), .ZN(n5555) );
NAND2_X2 U4645 ( .A1(w_q[251]), .A2(n7252), .ZN(n5554) );
NAND2_X2 U4646 ( .A1(n5556), .A2(n5557), .ZN(w_d[250]) );
NAND2_X2 U4647 ( .A1(w_q[218]), .A2(n7194), .ZN(n5557) );
NAND2_X2 U4648 ( .A1(w_q[250]), .A2(n7252), .ZN(n5556) );
NAND2_X2 U4650 ( .A1(w[24]), .A2(n7160), .ZN(n5560) );
NAND2_X2 U4651 ( .A1(w_q[24]), .A2(n7252), .ZN(n5559) );
NAND2_X2 U4653 ( .A1(n5561), .A2(n5562), .ZN(w_d[249]) );
NAND2_X2 U4654 ( .A1(w_q[217]), .A2(n7194), .ZN(n5562) );
NAND2_X2 U4655 ( .A1(w_q[249]), .A2(n7252), .ZN(n5561) );
NAND2_X2 U4656 ( .A1(n5563), .A2(n5564), .ZN(w_d[248]) );
NAND2_X2 U4657 ( .A1(w_q[216]), .A2(n7194), .ZN(n5564) );
NAND2_X2 U4658 ( .A1(w_q[248]), .A2(n7234), .ZN(n5563) );
NAND2_X2 U4659 ( .A1(n5565), .A2(n5566), .ZN(w_d[247]) );
NAND2_X2 U4660 ( .A1(w_q[215]), .A2(n7194), .ZN(n5566) );
NAND2_X2 U4661 ( .A1(w_q[247]), .A2(n7233), .ZN(n5565) );
NAND2_X2 U4662 ( .A1(n5567), .A2(n5568), .ZN(w_d[246]) );
NAND2_X2 U4663 ( .A1(w_q[214]), .A2(n7194), .ZN(n5568) );
NAND2_X2 U4664 ( .A1(w_q[246]), .A2(n7235), .ZN(n5567) );
NAND2_X2 U4665 ( .A1(n5569), .A2(n5570), .ZN(w_d[245]) );
NAND2_X2 U4666 ( .A1(w_q[213]), .A2(n7194), .ZN(n5570) );
NAND2_X2 U4667 ( .A1(w_q[245]), .A2(n7236), .ZN(n5569) );
NAND2_X2 U4668 ( .A1(n5571), .A2(n5572), .ZN(w_d[244]) );
NAND2_X2 U4669 ( .A1(w_q[212]), .A2(n7194), .ZN(n5572) );
NAND2_X2 U4670 ( .A1(w_q[244]), .A2(n7231), .ZN(n5571) );
NAND2_X2 U4671 ( .A1(n5573), .A2(n5574), .ZN(w_d[243]) );
NAND2_X2 U4672 ( .A1(w_q[211]), .A2(n7194), .ZN(n5574) );
NAND2_X2 U4673 ( .A1(w_q[243]), .A2(n7234), .ZN(n5573) );
NAND2_X2 U4674 ( .A1(n5575), .A2(n5576), .ZN(w_d[242]) );
NAND2_X2 U4675 ( .A1(w_q[210]), .A2(n7193), .ZN(n5576) );
NAND2_X2 U4676 ( .A1(w_q[242]), .A2(n7233), .ZN(n5575) );
NAND2_X2 U4677 ( .A1(n5577), .A2(n5578), .ZN(w_d[241]) );
NAND2_X2 U4678 ( .A1(w_q[209]), .A2(n7193), .ZN(n5578) );
NAND2_X2 U4679 ( .A1(w_q[241]), .A2(n7232), .ZN(n5577) );
NAND2_X2 U4680 ( .A1(n5579), .A2(n5580), .ZN(w_d[240]) );
NAND2_X2 U4681 ( .A1(w_q[208]), .A2(n7193), .ZN(n5580) );
NAND2_X2 U4682 ( .A1(w_q[240]), .A2(n7230), .ZN(n5579) );
NAND2_X2 U4684 ( .A1(w[23]), .A2(n7160), .ZN(n5583) );
NAND2_X2 U4685 ( .A1(w_q[23]), .A2(n7274), .ZN(n5582) );
NAND2_X2 U4687 ( .A1(n5584), .A2(n5585), .ZN(w_d[239]) );
NAND2_X2 U4688 ( .A1(w_q[207]), .A2(n7193), .ZN(n5585) );
NAND2_X2 U4689 ( .A1(w_q[239]), .A2(n7231), .ZN(n5584) );
NAND2_X2 U4690 ( .A1(n5586), .A2(n5587), .ZN(w_d[238]) );
NAND2_X2 U4691 ( .A1(w_q[206]), .A2(n7193), .ZN(n5587) );
NAND2_X2 U4692 ( .A1(w_q[238]), .A2(n7232), .ZN(n5586) );
NAND2_X2 U4693 ( .A1(n5588), .A2(n5589), .ZN(w_d[237]) );
NAND2_X2 U4694 ( .A1(w_q[205]), .A2(n7193), .ZN(n5589) );
NAND2_X2 U4695 ( .A1(w_q[237]), .A2(n7230), .ZN(n5588) );
NAND2_X2 U4696 ( .A1(n5590), .A2(n5591), .ZN(w_d[236]) );
NAND2_X2 U4697 ( .A1(w_q[204]), .A2(n7193), .ZN(n5591) );
NAND2_X2 U4698 ( .A1(w_q[236]), .A2(n7238), .ZN(n5590) );
NAND2_X2 U4699 ( .A1(n5592), .A2(n5593), .ZN(w_d[235]) );
NAND2_X2 U4700 ( .A1(w_q[203]), .A2(n7193), .ZN(n5593) );
NAND2_X2 U4701 ( .A1(w_q[235]), .A2(n7231), .ZN(n5592) );
NAND2_X2 U4702 ( .A1(n5594), .A2(n5595), .ZN(w_d[234]) );
NAND2_X2 U4703 ( .A1(w_q[202]), .A2(n7193), .ZN(n5595) );
NAND2_X2 U4704 ( .A1(w_q[234]), .A2(n7233), .ZN(n5594) );
NAND2_X2 U4705 ( .A1(n5596), .A2(n5597), .ZN(w_d[233]) );
NAND2_X2 U4706 ( .A1(w_q[201]), .A2(n7193), .ZN(n5597) );
NAND2_X2 U4707 ( .A1(w_q[233]), .A2(n7235), .ZN(n5596) );
NAND2_X2 U4708 ( .A1(n5598), .A2(n5599), .ZN(w_d[232]) );
NAND2_X2 U4709 ( .A1(w_q[200]), .A2(n7193), .ZN(n5599) );
NAND2_X2 U4710 ( .A1(w_q[232]), .A2(n7232), .ZN(n5598) );
NAND2_X2 U4711 ( .A1(n5600), .A2(n5601), .ZN(w_d[231]) );
NAND2_X2 U4712 ( .A1(w_q[199]), .A2(n7192), .ZN(n5601) );
NAND2_X2 U4713 ( .A1(w_q[231]), .A2(n7230), .ZN(n5600) );
NAND2_X2 U4714 ( .A1(n5602), .A2(n5603), .ZN(w_d[230]) );
NAND2_X2 U4715 ( .A1(w_q[198]), .A2(n7192), .ZN(n5603) );
NAND2_X2 U4716 ( .A1(w_q[230]), .A2(n7234), .ZN(n5602) );
NAND2_X2 U4718 ( .A1(w[22]), .A2(n7160), .ZN(n5606) );
NAND2_X2 U4719 ( .A1(w_q[22]), .A2(n7267), .ZN(n5605) );
NAND2_X2 U4721 ( .A1(n5607), .A2(n5608), .ZN(w_d[229]) );
NAND2_X2 U4722 ( .A1(w_q[197]), .A2(n7192), .ZN(n5608) );
NAND2_X2 U4723 ( .A1(w_q[229]), .A2(n7238), .ZN(n5607) );
NAND2_X2 U4724 ( .A1(n5609), .A2(n5610), .ZN(w_d[228]) );
NAND2_X2 U4725 ( .A1(w_q[196]), .A2(n7192), .ZN(n5610) );
NAND2_X2 U4726 ( .A1(w_q[228]), .A2(n7251), .ZN(n5609) );
NAND2_X2 U4727 ( .A1(n5611), .A2(n5612), .ZN(w_d[227]) );
NAND2_X2 U4728 ( .A1(w_q[195]), .A2(n7192), .ZN(n5612) );
NAND2_X2 U4729 ( .A1(w_q[227]), .A2(n7251), .ZN(n5611) );
NAND2_X2 U4730 ( .A1(n5613), .A2(n5614), .ZN(w_d[226]) );
NAND2_X2 U4731 ( .A1(w_q[194]), .A2(n7192), .ZN(n5614) );
NAND2_X2 U4732 ( .A1(w_q[226]), .A2(n7251), .ZN(n5613) );
NAND2_X2 U4733 ( .A1(n5615), .A2(n5616), .ZN(w_d[225]) );
NAND2_X2 U4734 ( .A1(w_q[193]), .A2(n7192), .ZN(n5616) );
NAND2_X2 U4735 ( .A1(w_q[225]), .A2(n7251), .ZN(n5615) );
NAND2_X2 U4736 ( .A1(n5617), .A2(n5618), .ZN(w_d[224]) );
NAND2_X2 U4737 ( .A1(w_q[192]), .A2(n7192), .ZN(n5618) );
NAND2_X2 U4738 ( .A1(w_q[224]), .A2(n7251), .ZN(n5617) );
NAND2_X2 U4739 ( .A1(n5619), .A2(n5620), .ZN(w_d[223]) );
NAND2_X2 U4740 ( .A1(w_q[191]), .A2(n7192), .ZN(n5620) );
NAND2_X2 U4741 ( .A1(w_q[223]), .A2(n7251), .ZN(n5619) );
NAND2_X2 U4742 ( .A1(n5621), .A2(n5622), .ZN(w_d[222]) );
NAND2_X2 U4743 ( .A1(w_q[190]), .A2(n7192), .ZN(n5622) );
NAND2_X2 U4744 ( .A1(w_q[222]), .A2(n7251), .ZN(n5621) );
NAND2_X2 U4745 ( .A1(n5623), .A2(n5624), .ZN(w_d[221]) );
NAND2_X2 U4746 ( .A1(w_q[189]), .A2(n7192), .ZN(n5624) );
NAND2_X2 U4747 ( .A1(w_q[221]), .A2(n7251), .ZN(n5623) );
NAND2_X2 U4748 ( .A1(n5625), .A2(n5626), .ZN(w_d[220]) );
NAND2_X2 U4749 ( .A1(w_q[188]), .A2(n7191), .ZN(n5626) );
NAND2_X2 U4750 ( .A1(w_q[220]), .A2(n7251), .ZN(n5625) );
NAND2_X2 U4752 ( .A1(w[21]), .A2(n7160), .ZN(n5629) );
NAND2_X2 U4753 ( .A1(w_q[21]), .A2(n7251), .ZN(n5628) );
NAND2_X2 U4755 ( .A1(n5630), .A2(n5631), .ZN(w_d[219]) );
NAND2_X2 U4756 ( .A1(w_q[187]), .A2(n7191), .ZN(n5631) );
NAND2_X2 U4757 ( .A1(w_q[219]), .A2(n7251), .ZN(n5630) );
NAND2_X2 U4758 ( .A1(n5632), .A2(n5633), .ZN(w_d[218]) );
NAND2_X2 U4759 ( .A1(w_q[186]), .A2(n7191), .ZN(n5633) );
NAND2_X2 U4760 ( .A1(w_q[218]), .A2(n7250), .ZN(n5632) );
NAND2_X2 U4761 ( .A1(n5634), .A2(n5635), .ZN(w_d[217]) );
NAND2_X2 U4762 ( .A1(w_q[185]), .A2(n7191), .ZN(n5635) );
NAND2_X2 U4763 ( .A1(w_q[217]), .A2(n7250), .ZN(n5634) );
NAND2_X2 U4764 ( .A1(n5636), .A2(n5637), .ZN(w_d[216]) );
NAND2_X2 U4765 ( .A1(w_q[184]), .A2(n7191), .ZN(n5637) );
NAND2_X2 U4766 ( .A1(w_q[216]), .A2(n7250), .ZN(n5636) );
NAND2_X2 U4767 ( .A1(n5638), .A2(n5639), .ZN(w_d[215]) );
NAND2_X2 U4768 ( .A1(w_q[183]), .A2(n7191), .ZN(n5639) );
NAND2_X2 U4769 ( .A1(w_q[215]), .A2(n7250), .ZN(n5638) );
NAND2_X2 U4770 ( .A1(n5640), .A2(n5641), .ZN(w_d[214]) );
NAND2_X2 U4771 ( .A1(w_q[182]), .A2(n7191), .ZN(n5641) );
NAND2_X2 U4772 ( .A1(w_q[214]), .A2(n7250), .ZN(n5640) );
NAND2_X2 U4773 ( .A1(n5642), .A2(n5643), .ZN(w_d[213]) );
NAND2_X2 U4774 ( .A1(w_q[181]), .A2(n7191), .ZN(n5643) );
NAND2_X2 U4775 ( .A1(w_q[213]), .A2(n7250), .ZN(n5642) );
NAND2_X2 U4776 ( .A1(n5644), .A2(n5645), .ZN(w_d[212]) );
NAND2_X2 U4777 ( .A1(w_q[180]), .A2(n7191), .ZN(n5645) );
NAND2_X2 U4778 ( .A1(w_q[212]), .A2(n7250), .ZN(n5644) );
NAND2_X2 U4779 ( .A1(n5646), .A2(n5647), .ZN(w_d[211]) );
NAND2_X2 U4780 ( .A1(w_q[179]), .A2(n7191), .ZN(n5647) );
NAND2_X2 U4781 ( .A1(w_q[211]), .A2(n7250), .ZN(n5646) );
NAND2_X2 U4782 ( .A1(n5648), .A2(n5649), .ZN(w_d[210]) );
NAND2_X2 U4783 ( .A1(w_q[178]), .A2(n7191), .ZN(n5649) );
NAND2_X2 U4784 ( .A1(w_q[210]), .A2(n7250), .ZN(n5648) );
NAND2_X2 U4786 ( .A1(w[20]), .A2(n7160), .ZN(n5652) );
NAND2_X2 U4787 ( .A1(w_q[20]), .A2(n7250), .ZN(n5651) );
NAND2_X2 U4789 ( .A1(n5653), .A2(n5654), .ZN(w_d[209]) );
NAND2_X2 U4790 ( .A1(w_q[177]), .A2(n7190), .ZN(n5654) );
NAND2_X2 U4791 ( .A1(w_q[209]), .A2(n7250), .ZN(n5653) );
NAND2_X2 U4792 ( .A1(n5655), .A2(n5656), .ZN(w_d[208]) );
NAND2_X2 U4793 ( .A1(w_q[176]), .A2(n7190), .ZN(n5656) );
NAND2_X2 U4794 ( .A1(w_q[208]), .A2(n7249), .ZN(n5655) );
NAND2_X2 U4795 ( .A1(n5657), .A2(n5658), .ZN(w_d[207]) );
NAND2_X2 U4796 ( .A1(w_q[175]), .A2(n7190), .ZN(n5658) );
NAND2_X2 U4797 ( .A1(w_q[207]), .A2(n7249), .ZN(n5657) );
NAND2_X2 U4798 ( .A1(n5659), .A2(n5660), .ZN(w_d[206]) );
NAND2_X2 U4799 ( .A1(w_q[174]), .A2(n7190), .ZN(n5660) );
NAND2_X2 U4800 ( .A1(w_q[206]), .A2(n7249), .ZN(n5659) );
NAND2_X2 U4801 ( .A1(n5661), .A2(n5662), .ZN(w_d[205]) );
NAND2_X2 U4802 ( .A1(w_q[173]), .A2(n7190), .ZN(n5662) );
NAND2_X2 U4803 ( .A1(w_q[205]), .A2(n7249), .ZN(n5661) );
NAND2_X2 U4804 ( .A1(n5663), .A2(n5664), .ZN(w_d[204]) );
NAND2_X2 U4805 ( .A1(w_q[172]), .A2(n7190), .ZN(n5664) );
NAND2_X2 U4806 ( .A1(w_q[204]), .A2(n7249), .ZN(n5663) );
NAND2_X2 U4807 ( .A1(n5665), .A2(n5666), .ZN(w_d[203]) );
NAND2_X2 U4808 ( .A1(w_q[171]), .A2(n7190), .ZN(n5666) );
NAND2_X2 U4809 ( .A1(w_q[203]), .A2(n7249), .ZN(n5665) );
NAND2_X2 U4810 ( .A1(n5667), .A2(n5668), .ZN(w_d[202]) );
NAND2_X2 U4811 ( .A1(w_q[170]), .A2(n7190), .ZN(n5668) );
NAND2_X2 U4812 ( .A1(w_q[202]), .A2(n7249), .ZN(n5667) );
NAND2_X2 U4813 ( .A1(n5669), .A2(n5670), .ZN(w_d[201]) );
NAND2_X2 U4814 ( .A1(w_q[169]), .A2(n7190), .ZN(n5670) );
NAND2_X2 U4815 ( .A1(w_q[201]), .A2(n7249), .ZN(n5669) );
NAND2_X2 U4816 ( .A1(n5671), .A2(n5672), .ZN(w_d[200]) );
NAND2_X2 U4817 ( .A1(w_q[168]), .A2(n7190), .ZN(n5672) );
NAND2_X2 U4818 ( .A1(w_q[200]), .A2(n7249), .ZN(n5671) );
NAND2_X2 U4820 ( .A1(w[1]), .A2(n7160), .ZN(n5675) );
NAND2_X2 U4821 ( .A1(w_q[1]), .A2(n7249), .ZN(n5674) );
NAND2_X2 U4824 ( .A1(w[19]), .A2(n7160), .ZN(n5678) );
NAND2_X2 U4825 ( .A1(w_q[19]), .A2(n7249), .ZN(n5677) );
NAND2_X2 U4827 ( .A1(n5679), .A2(n5680), .ZN(w_d[199]) );
NAND2_X2 U4828 ( .A1(w_q[167]), .A2(n7190), .ZN(n5680) );
NAND2_X2 U4829 ( .A1(w_q[199]), .A2(n7248), .ZN(n5679) );
NAND2_X2 U4830 ( .A1(n5681), .A2(n5682), .ZN(w_d[198]) );
NAND2_X2 U4831 ( .A1(w_q[166]), .A2(n7189), .ZN(n5682) );
NAND2_X2 U4832 ( .A1(w_q[198]), .A2(n7248), .ZN(n5681) );
NAND2_X2 U4833 ( .A1(n5683), .A2(n5684), .ZN(w_d[197]) );
NAND2_X2 U4834 ( .A1(w_q[165]), .A2(n7189), .ZN(n5684) );
NAND2_X2 U4835 ( .A1(w_q[197]), .A2(n7248), .ZN(n5683) );
NAND2_X2 U4836 ( .A1(n5685), .A2(n5686), .ZN(w_d[196]) );
NAND2_X2 U4837 ( .A1(w_q[164]), .A2(n7189), .ZN(n5686) );
NAND2_X2 U4838 ( .A1(w_q[196]), .A2(n7248), .ZN(n5685) );
NAND2_X2 U4839 ( .A1(n5687), .A2(n5688), .ZN(w_d[195]) );
NAND2_X2 U4840 ( .A1(w_q[163]), .A2(n7189), .ZN(n5688) );
NAND2_X2 U4841 ( .A1(w_q[195]), .A2(n7248), .ZN(n5687) );
NAND2_X2 U4842 ( .A1(n5689), .A2(n5690), .ZN(w_d[194]) );
NAND2_X2 U4843 ( .A1(w_q[162]), .A2(n7189), .ZN(n5690) );
NAND2_X2 U4844 ( .A1(w_q[194]), .A2(n7248), .ZN(n5689) );
NAND2_X2 U4845 ( .A1(n5691), .A2(n5692), .ZN(w_d[193]) );
NAND2_X2 U4846 ( .A1(w_q[161]), .A2(n7189), .ZN(n5692) );
NAND2_X2 U4847 ( .A1(w_q[193]), .A2(n7248), .ZN(n5691) );
NAND2_X2 U4848 ( .A1(n5693), .A2(n5694), .ZN(w_d[192]) );
NAND2_X2 U4849 ( .A1(w_q[160]), .A2(n7189), .ZN(n5694) );
NAND2_X2 U4850 ( .A1(w_q[192]), .A2(n7248), .ZN(n5693) );
NAND2_X2 U4851 ( .A1(n5695), .A2(n5696), .ZN(w_d[191]) );
NAND2_X2 U4852 ( .A1(w_q[159]), .A2(n7189), .ZN(n5696) );
NAND2_X2 U4853 ( .A1(w_q[191]), .A2(n7248), .ZN(n5695) );
NAND2_X2 U4854 ( .A1(n5697), .A2(n5698), .ZN(w_d[190]) );
NAND2_X2 U4855 ( .A1(w_q[158]), .A2(n7189), .ZN(n5698) );
NAND2_X2 U4856 ( .A1(w_q[190]), .A2(n7248), .ZN(n5697) );
NAND2_X2 U4858 ( .A1(w[18]), .A2(n7160), .ZN(n5701) );
NAND2_X2 U4859 ( .A1(w_q[18]), .A2(n7248), .ZN(n5700) );
NAND2_X2 U4861 ( .A1(n5702), .A2(n5703), .ZN(w_d[189]) );
NAND2_X2 U4862 ( .A1(w_q[157]), .A2(n7189), .ZN(n5703) );
NAND2_X2 U4863 ( .A1(w_q[189]), .A2(n7247), .ZN(n5702) );
NAND2_X2 U4864 ( .A1(n5704), .A2(n5705), .ZN(w_d[188]) );
NAND2_X2 U4865 ( .A1(w_q[156]), .A2(n7189), .ZN(n5705) );
NAND2_X2 U4866 ( .A1(w_q[188]), .A2(n7247), .ZN(n5704) );
NAND2_X2 U4867 ( .A1(n5706), .A2(n5707), .ZN(w_d[187]) );
NAND2_X2 U4868 ( .A1(w_q[155]), .A2(n7188), .ZN(n5707) );
NAND2_X2 U4869 ( .A1(w_q[187]), .A2(n7247), .ZN(n5706) );
NAND2_X2 U4870 ( .A1(n5708), .A2(n5709), .ZN(w_d[186]) );
NAND2_X2 U4871 ( .A1(w_q[154]), .A2(n7188), .ZN(n5709) );
NAND2_X2 U4872 ( .A1(w_q[186]), .A2(n7247), .ZN(n5708) );
NAND2_X2 U4873 ( .A1(n5710), .A2(n5711), .ZN(w_d[185]) );
NAND2_X2 U4874 ( .A1(w_q[153]), .A2(n7188), .ZN(n5711) );
NAND2_X2 U4875 ( .A1(w_q[185]), .A2(n7247), .ZN(n5710) );
NAND2_X2 U4876 ( .A1(n5712), .A2(n5713), .ZN(w_d[184]) );
NAND2_X2 U4877 ( .A1(w_q[152]), .A2(n7188), .ZN(n5713) );
NAND2_X2 U4878 ( .A1(w_q[184]), .A2(n7247), .ZN(n5712) );
NAND2_X2 U4879 ( .A1(n5714), .A2(n5715), .ZN(w_d[183]) );
NAND2_X2 U4880 ( .A1(w_q[151]), .A2(n7188), .ZN(n5715) );
NAND2_X2 U4881 ( .A1(w_q[183]), .A2(n7247), .ZN(n5714) );
NAND2_X2 U4882 ( .A1(n5716), .A2(n5717), .ZN(w_d[182]) );
NAND2_X2 U4883 ( .A1(w_q[150]), .A2(n7188), .ZN(n5717) );
NAND2_X2 U4884 ( .A1(w_q[182]), .A2(n7247), .ZN(n5716) );
NAND2_X2 U4885 ( .A1(n5718), .A2(n5719), .ZN(w_d[181]) );
NAND2_X2 U4886 ( .A1(w_q[149]), .A2(n7188), .ZN(n5719) );
NAND2_X2 U4887 ( .A1(w_q[181]), .A2(n7247), .ZN(n5718) );
NAND2_X2 U4888 ( .A1(n5720), .A2(n5721), .ZN(w_d[180]) );
NAND2_X2 U4889 ( .A1(w_q[148]), .A2(n7188), .ZN(n5721) );
NAND2_X2 U4890 ( .A1(w_q[180]), .A2(n7247), .ZN(n5720) );
NAND2_X2 U4892 ( .A1(w[17]), .A2(n7160), .ZN(n5724) );
NAND2_X2 U4893 ( .A1(w_q[17]), .A2(n7247), .ZN(n5723) );
NAND2_X2 U4895 ( .A1(n5725), .A2(n5726), .ZN(w_d[179]) );
NAND2_X2 U4896 ( .A1(w_q[147]), .A2(n7188), .ZN(n5726) );
NAND2_X2 U4897 ( .A1(w_q[179]), .A2(n7246), .ZN(n5725) );
NAND2_X2 U4898 ( .A1(n5727), .A2(n5728), .ZN(w_d[178]) );
NAND2_X2 U4899 ( .A1(w_q[146]), .A2(n7188), .ZN(n5728) );
NAND2_X2 U4900 ( .A1(w_q[178]), .A2(n7246), .ZN(n5727) );
NAND2_X2 U4901 ( .A1(n5729), .A2(n5730), .ZN(w_d[177]) );
NAND2_X2 U4902 ( .A1(w_q[145]), .A2(n7188), .ZN(n5730) );
NAND2_X2 U4903 ( .A1(w_q[177]), .A2(n7246), .ZN(n5729) );
NAND2_X2 U4904 ( .A1(n5731), .A2(n5732), .ZN(w_d[176]) );
NAND2_X2 U4905 ( .A1(w_q[144]), .A2(n7187), .ZN(n5732) );
NAND2_X2 U4906 ( .A1(w_q[176]), .A2(n7246), .ZN(n5731) );
NAND2_X2 U4907 ( .A1(n5733), .A2(n5734), .ZN(w_d[175]) );
NAND2_X2 U4908 ( .A1(w_q[143]), .A2(n7187), .ZN(n5734) );
NAND2_X2 U4909 ( .A1(w_q[175]), .A2(n7246), .ZN(n5733) );
NAND2_X2 U4910 ( .A1(n5735), .A2(n5736), .ZN(w_d[174]) );
NAND2_X2 U4911 ( .A1(w_q[142]), .A2(n7187), .ZN(n5736) );
NAND2_X2 U4912 ( .A1(w_q[174]), .A2(n7246), .ZN(n5735) );
NAND2_X2 U4913 ( .A1(n5737), .A2(n5738), .ZN(w_d[173]) );
NAND2_X2 U4914 ( .A1(w_q[141]), .A2(n7187), .ZN(n5738) );
NAND2_X2 U4915 ( .A1(w_q[173]), .A2(n7246), .ZN(n5737) );
NAND2_X2 U4916 ( .A1(n5739), .A2(n5740), .ZN(w_d[172]) );
NAND2_X2 U4917 ( .A1(w_q[140]), .A2(n7187), .ZN(n5740) );
NAND2_X2 U4918 ( .A1(w_q[172]), .A2(n7246), .ZN(n5739) );
NAND2_X2 U4919 ( .A1(n5741), .A2(n5742), .ZN(w_d[171]) );
NAND2_X2 U4920 ( .A1(w_q[139]), .A2(n7187), .ZN(n5742) );
NAND2_X2 U4921 ( .A1(w_q[171]), .A2(n7246), .ZN(n5741) );
NAND2_X2 U4922 ( .A1(n5743), .A2(n5744), .ZN(w_d[170]) );
NAND2_X2 U4923 ( .A1(w_q[138]), .A2(n7187), .ZN(n5744) );
NAND2_X2 U4924 ( .A1(w_q[170]), .A2(n7246), .ZN(n5743) );
NAND2_X2 U4926 ( .A1(w[16]), .A2(n7160), .ZN(n5747) );
NAND2_X2 U4927 ( .A1(w_q[16]), .A2(n7246), .ZN(n5746) );
NAND2_X2 U4929 ( .A1(n5748), .A2(n5749), .ZN(w_d[169]) );
NAND2_X2 U4930 ( .A1(w_q[137]), .A2(n7187), .ZN(n5749) );
NAND2_X2 U4931 ( .A1(w_q[169]), .A2(n7245), .ZN(n5748) );
NAND2_X2 U4932 ( .A1(n5750), .A2(n5751), .ZN(w_d[168]) );
NAND2_X2 U4933 ( .A1(w_q[136]), .A2(n7187), .ZN(n5751) );
NAND2_X2 U4934 ( .A1(w_q[168]), .A2(n7245), .ZN(n5750) );
NAND2_X2 U4935 ( .A1(n5752), .A2(n5753), .ZN(w_d[167]) );
NAND2_X2 U4936 ( .A1(w_q[135]), .A2(n7187), .ZN(n5753) );
NAND2_X2 U4937 ( .A1(w_q[167]), .A2(n7245), .ZN(n5752) );
NAND2_X2 U4938 ( .A1(n5754), .A2(n5755), .ZN(w_d[166]) );
NAND2_X2 U4939 ( .A1(w_q[134]), .A2(n7187), .ZN(n5755) );
NAND2_X2 U4940 ( .A1(w_q[166]), .A2(n7245), .ZN(n5754) );
NAND2_X2 U4941 ( .A1(n5756), .A2(n5757), .ZN(w_d[165]) );
NAND2_X2 U4942 ( .A1(w_q[133]), .A2(n7186), .ZN(n5757) );
NAND2_X2 U4943 ( .A1(w_q[165]), .A2(n7245), .ZN(n5756) );
NAND2_X2 U4944 ( .A1(n5758), .A2(n5759), .ZN(w_d[164]) );
NAND2_X2 U4945 ( .A1(w_q[132]), .A2(n7186), .ZN(n5759) );
NAND2_X2 U4946 ( .A1(w_q[164]), .A2(n7245), .ZN(n5758) );
NAND2_X2 U4947 ( .A1(n5760), .A2(n5761), .ZN(w_d[163]) );
NAND2_X2 U4948 ( .A1(w_q[131]), .A2(n7186), .ZN(n5761) );
NAND2_X2 U4949 ( .A1(w_q[163]), .A2(n7245), .ZN(n5760) );
NAND2_X2 U4950 ( .A1(n5762), .A2(n5763), .ZN(w_d[162]) );
NAND2_X2 U4951 ( .A1(w_q[130]), .A2(n7186), .ZN(n5763) );
NAND2_X2 U4952 ( .A1(w_q[162]), .A2(n7245), .ZN(n5762) );
NAND2_X2 U4953 ( .A1(n5764), .A2(n5765), .ZN(w_d[161]) );
NAND2_X2 U4954 ( .A1(w_q[129]), .A2(n7186), .ZN(n5765) );
NAND2_X2 U4955 ( .A1(w_q[161]), .A2(n7245), .ZN(n5764) );
NAND2_X2 U4956 ( .A1(n5766), .A2(n5767), .ZN(w_d[160]) );
NAND2_X2 U4957 ( .A1(w_q[128]), .A2(n7186), .ZN(n5767) );
NAND2_X2 U4958 ( .A1(w_q[160]), .A2(n7245), .ZN(n5766) );
NAND2_X2 U4960 ( .A1(w[15]), .A2(n7160), .ZN(n5770) );
NAND2_X2 U4961 ( .A1(w_q[15]), .A2(n7245), .ZN(n5769) );
NAND2_X2 U4963 ( .A1(n5771), .A2(n5772), .ZN(w_d[159]) );
NAND2_X2 U4964 ( .A1(w_q[127]), .A2(n7186), .ZN(n5772) );
NAND2_X2 U4965 ( .A1(w_q[159]), .A2(n7244), .ZN(n5771) );
NAND2_X2 U4966 ( .A1(n5773), .A2(n5774), .ZN(w_d[158]) );
NAND2_X2 U4967 ( .A1(w_q[126]), .A2(n7186), .ZN(n5774) );
NAND2_X2 U4968 ( .A1(w_q[158]), .A2(n7244), .ZN(n5773) );
NAND2_X2 U4969 ( .A1(n5775), .A2(n5776), .ZN(w_d[157]) );
NAND2_X2 U4970 ( .A1(w_q[125]), .A2(n7186), .ZN(n5776) );
NAND2_X2 U4971 ( .A1(w_q[157]), .A2(n7244), .ZN(n5775) );
NAND2_X2 U4972 ( .A1(n5777), .A2(n5778), .ZN(w_d[156]) );
NAND2_X2 U4973 ( .A1(w_q[124]), .A2(n7186), .ZN(n5778) );
NAND2_X2 U4974 ( .A1(w_q[156]), .A2(n7244), .ZN(n5777) );
NAND2_X2 U4975 ( .A1(n5779), .A2(n5780), .ZN(w_d[155]) );
NAND2_X2 U4976 ( .A1(w_q[123]), .A2(n7186), .ZN(n5780) );
NAND2_X2 U4977 ( .A1(w_q[155]), .A2(n7244), .ZN(n5779) );
NAND2_X2 U4978 ( .A1(n5781), .A2(n5782), .ZN(w_d[154]) );
NAND2_X2 U4979 ( .A1(w_q[122]), .A2(n7185), .ZN(n5782) );
NAND2_X2 U4980 ( .A1(w_q[154]), .A2(n7244), .ZN(n5781) );
NAND2_X2 U4981 ( .A1(n5783), .A2(n5784), .ZN(w_d[153]) );
NAND2_X2 U4982 ( .A1(w_q[121]), .A2(n7185), .ZN(n5784) );
NAND2_X2 U4983 ( .A1(w_q[153]), .A2(n7244), .ZN(n5783) );
NAND2_X2 U4984 ( .A1(n5785), .A2(n5786), .ZN(w_d[152]) );
NAND2_X2 U4985 ( .A1(w_q[120]), .A2(n7185), .ZN(n5786) );
NAND2_X2 U4986 ( .A1(w_q[152]), .A2(n7244), .ZN(n5785) );
NAND2_X2 U4987 ( .A1(n5787), .A2(n5788), .ZN(w_d[151]) );
NAND2_X2 U4988 ( .A1(w_q[119]), .A2(n7185), .ZN(n5788) );
NAND2_X2 U4989 ( .A1(w_q[151]), .A2(n7244), .ZN(n5787) );
NAND2_X2 U4990 ( .A1(n5789), .A2(n5790), .ZN(w_d[150]) );
NAND2_X2 U4991 ( .A1(w_q[118]), .A2(n7185), .ZN(n5790) );
NAND2_X2 U4992 ( .A1(w_q[150]), .A2(n7244), .ZN(n5789) );
NAND2_X2 U4994 ( .A1(w[14]), .A2(n7160), .ZN(n5793) );
NAND2_X2 U4995 ( .A1(w_q[14]), .A2(n7244), .ZN(n5792) );
NAND2_X2 U4997 ( .A1(n5794), .A2(n5795), .ZN(w_d[149]) );
NAND2_X2 U4998 ( .A1(w_q[117]), .A2(n7185), .ZN(n5795) );
NAND2_X2 U4999 ( .A1(w_q[149]), .A2(n7243), .ZN(n5794) );
NAND2_X2 U5000 ( .A1(n5796), .A2(n5797), .ZN(w_d[148]) );
NAND2_X2 U5001 ( .A1(w_q[116]), .A2(n7185), .ZN(n5797) );
NAND2_X2 U5002 ( .A1(w_q[148]), .A2(n7243), .ZN(n5796) );
NAND2_X2 U5003 ( .A1(n5798), .A2(n5799), .ZN(w_d[147]) );
NAND2_X2 U5004 ( .A1(w_q[115]), .A2(n7185), .ZN(n5799) );
NAND2_X2 U5005 ( .A1(w_q[147]), .A2(n7243), .ZN(n5798) );
NAND2_X2 U5006 ( .A1(n5800), .A2(n5801), .ZN(w_d[146]) );
NAND2_X2 U5007 ( .A1(w_q[114]), .A2(n7185), .ZN(n5801) );
NAND2_X2 U5008 ( .A1(w_q[146]), .A2(n7243), .ZN(n5800) );
NAND2_X2 U5009 ( .A1(n5802), .A2(n5803), .ZN(w_d[145]) );
NAND2_X2 U5010 ( .A1(w_q[113]), .A2(n7185), .ZN(n5803) );
NAND2_X2 U5011 ( .A1(w_q[145]), .A2(n7243), .ZN(n5802) );
NAND2_X2 U5012 ( .A1(n5804), .A2(n5805), .ZN(w_d[144]) );
NAND2_X2 U5013 ( .A1(w_q[112]), .A2(n7185), .ZN(n5805) );
NAND2_X2 U5014 ( .A1(w_q[144]), .A2(n7243), .ZN(n5804) );
NAND2_X2 U5015 ( .A1(n5806), .A2(n5807), .ZN(w_d[143]) );
NAND2_X2 U5016 ( .A1(w_q[111]), .A2(n7184), .ZN(n5807) );
NAND2_X2 U5017 ( .A1(w_q[143]), .A2(n7243), .ZN(n5806) );
NAND2_X2 U5018 ( .A1(n5808), .A2(n5809), .ZN(w_d[142]) );
NAND2_X2 U5019 ( .A1(w_q[110]), .A2(n7184), .ZN(n5809) );
NAND2_X2 U5020 ( .A1(w_q[142]), .A2(n7243), .ZN(n5808) );
NAND2_X2 U5021 ( .A1(n5810), .A2(n5811), .ZN(w_d[141]) );
NAND2_X2 U5022 ( .A1(w_q[109]), .A2(n7184), .ZN(n5811) );
NAND2_X2 U5023 ( .A1(w_q[141]), .A2(n7243), .ZN(n5810) );
NAND2_X2 U5024 ( .A1(n5812), .A2(n5813), .ZN(w_d[140]) );
NAND2_X2 U5025 ( .A1(w_q[108]), .A2(n7184), .ZN(n5813) );
NAND2_X2 U5026 ( .A1(w_q[140]), .A2(n7243), .ZN(n5812) );
NAND2_X2 U5028 ( .A1(w[13]), .A2(n7160), .ZN(n5816) );
NAND2_X2 U5029 ( .A1(w_q[13]), .A2(n7243), .ZN(n5815) );
NAND2_X2 U5031 ( .A1(n5817), .A2(n5818), .ZN(w_d[139]) );
NAND2_X2 U5032 ( .A1(w_q[107]), .A2(n7184), .ZN(n5818) );
NAND2_X2 U5033 ( .A1(w_q[139]), .A2(n7242), .ZN(n5817) );
NAND2_X2 U5034 ( .A1(n5819), .A2(n5820), .ZN(w_d[138]) );
NAND2_X2 U5035 ( .A1(w_q[106]), .A2(n7184), .ZN(n5820) );
NAND2_X2 U5036 ( .A1(w_q[138]), .A2(n7242), .ZN(n5819) );
NAND2_X2 U5037 ( .A1(n5821), .A2(n5822), .ZN(w_d[137]) );
NAND2_X2 U5038 ( .A1(w_q[105]), .A2(n7184), .ZN(n5822) );
NAND2_X2 U5039 ( .A1(w_q[137]), .A2(n7242), .ZN(n5821) );
NAND2_X2 U5040 ( .A1(n5823), .A2(n5824), .ZN(w_d[136]) );
NAND2_X2 U5041 ( .A1(w_q[104]), .A2(n7184), .ZN(n5824) );
NAND2_X2 U5042 ( .A1(w_q[136]), .A2(n7242), .ZN(n5823) );
NAND2_X2 U5043 ( .A1(n5825), .A2(n5826), .ZN(w_d[135]) );
NAND2_X2 U5044 ( .A1(w_q[103]), .A2(n7184), .ZN(n5826) );
NAND2_X2 U5045 ( .A1(w_q[135]), .A2(n7242), .ZN(n5825) );
NAND2_X2 U5046 ( .A1(n5827), .A2(n5828), .ZN(w_d[134]) );
NAND2_X2 U5047 ( .A1(w_q[102]), .A2(n7184), .ZN(n5828) );
NAND2_X2 U5048 ( .A1(w_q[134]), .A2(n7242), .ZN(n5827) );
NAND2_X2 U5049 ( .A1(n5829), .A2(n5830), .ZN(w_d[133]) );
NAND2_X2 U5050 ( .A1(w_q[101]), .A2(n7184), .ZN(n5830) );
NAND2_X2 U5051 ( .A1(w_q[133]), .A2(n7242), .ZN(n5829) );
NAND2_X2 U5052 ( .A1(n5831), .A2(n5832), .ZN(w_d[132]) );
NAND2_X2 U5053 ( .A1(w_q[100]), .A2(n7183), .ZN(n5832) );
NAND2_X2 U5054 ( .A1(w_q[132]), .A2(n7242), .ZN(n5831) );
NAND2_X2 U5055 ( .A1(n5833), .A2(n5834), .ZN(w_d[131]) );
NAND2_X2 U5056 ( .A1(w_q[99]), .A2(n7183), .ZN(n5834) );
NAND2_X2 U5057 ( .A1(w_q[131]), .A2(n7242), .ZN(n5833) );
NAND2_X2 U5058 ( .A1(n5835), .A2(n5836), .ZN(w_d[130]) );
NAND2_X2 U5059 ( .A1(w_q[98]), .A2(n7183), .ZN(n5836) );
NAND2_X2 U5060 ( .A1(w_q[130]), .A2(n7242), .ZN(n5835) );
NAND2_X2 U5062 ( .A1(w[12]), .A2(n7160), .ZN(n5839) );
NAND2_X2 U5063 ( .A1(w_q[12]), .A2(n7242), .ZN(n5838) );
NAND2_X2 U5065 ( .A1(n5840), .A2(n5841), .ZN(w_d[129]) );
NAND2_X2 U5066 ( .A1(w_q[97]), .A2(n7183), .ZN(n5841) );
NAND2_X2 U5067 ( .A1(w_q[129]), .A2(n7241), .ZN(n5840) );
NAND2_X2 U5068 ( .A1(n5842), .A2(n5843), .ZN(w_d[128]) );
NAND2_X2 U5069 ( .A1(w_q[96]), .A2(n7183), .ZN(n5843) );
NAND2_X2 U5070 ( .A1(w_q[128]), .A2(n7241), .ZN(n5842) );
NAND2_X2 U5071 ( .A1(n5844), .A2(n5845), .ZN(w_d[127]) );
NAND2_X2 U5072 ( .A1(w_q[95]), .A2(n7183), .ZN(n5845) );
NAND2_X2 U5073 ( .A1(w_q[127]), .A2(n7241), .ZN(n5844) );
NAND2_X2 U5074 ( .A1(n5846), .A2(n5847), .ZN(w_d[126]) );
NAND2_X2 U5075 ( .A1(w_q[94]), .A2(n7183), .ZN(n5847) );
NAND2_X2 U5076 ( .A1(w_q[126]), .A2(n7241), .ZN(n5846) );
NAND2_X2 U5077 ( .A1(n5848), .A2(n5849), .ZN(w_d[125]) );
NAND2_X2 U5078 ( .A1(w_q[93]), .A2(n7183), .ZN(n5849) );
NAND2_X2 U5079 ( .A1(w_q[125]), .A2(n7241), .ZN(n5848) );
NAND2_X2 U5080 ( .A1(n5850), .A2(n5851), .ZN(w_d[124]) );
NAND2_X2 U5081 ( .A1(w_q[92]), .A2(n7183), .ZN(n5851) );
NAND2_X2 U5082 ( .A1(w_q[124]), .A2(n7241), .ZN(n5850) );
NAND2_X2 U5083 ( .A1(n5852), .A2(n5853), .ZN(w_d[123]) );
NAND2_X2 U5084 ( .A1(w_q[91]), .A2(n7183), .ZN(n5853) );
NAND2_X2 U5085 ( .A1(w_q[123]), .A2(n7241), .ZN(n5852) );
NAND2_X2 U5086 ( .A1(n5854), .A2(n5855), .ZN(w_d[122]) );
NAND2_X2 U5087 ( .A1(w_q[90]), .A2(n7183), .ZN(n5855) );
NAND2_X2 U5088 ( .A1(w_q[122]), .A2(n7241), .ZN(n5854) );
NAND2_X2 U5089 ( .A1(n5856), .A2(n5857), .ZN(w_d[121]) );
NAND2_X2 U5090 ( .A1(w_q[89]), .A2(n7216), .ZN(n5857) );
NAND2_X2 U5091 ( .A1(w_q[121]), .A2(n7241), .ZN(n5856) );
NAND2_X2 U5092 ( .A1(n5858), .A2(n5859), .ZN(w_d[120]) );
NAND2_X2 U5093 ( .A1(w_q[88]), .A2(n7216), .ZN(n5859) );
NAND2_X2 U5094 ( .A1(w_q[120]), .A2(n7241), .ZN(n5858) );
NAND2_X2 U5096 ( .A1(w[11]), .A2(n7160), .ZN(n5862) );
NAND2_X2 U5097 ( .A1(w_q[11]), .A2(n7241), .ZN(n5861) );
NAND2_X2 U5099 ( .A1(n5863), .A2(n5864), .ZN(w_d[119]) );
NAND2_X2 U5100 ( .A1(w_q[87]), .A2(n7216), .ZN(n5864) );
NAND2_X2 U5101 ( .A1(w_q[119]), .A2(n7240), .ZN(n5863) );
NAND2_X2 U5102 ( .A1(n5865), .A2(n5866), .ZN(w_d[118]) );
NAND2_X2 U5103 ( .A1(w_q[86]), .A2(n7182), .ZN(n5866) );
NAND2_X2 U5104 ( .A1(w_q[118]), .A2(n7240), .ZN(n5865) );
NAND2_X2 U5105 ( .A1(n5867), .A2(n5868), .ZN(w_d[117]) );
NAND2_X2 U5106 ( .A1(w_q[85]), .A2(n7226), .ZN(n5868) );
NAND2_X2 U5107 ( .A1(w_q[117]), .A2(n7240), .ZN(n5867) );
NAND2_X2 U5108 ( .A1(n5869), .A2(n5870), .ZN(w_d[116]) );
NAND2_X2 U5109 ( .A1(w_q[84]), .A2(n7216), .ZN(n5870) );
NAND2_X2 U5110 ( .A1(w_q[116]), .A2(n7240), .ZN(n5869) );
NAND2_X2 U5111 ( .A1(n5871), .A2(n5872), .ZN(w_d[115]) );
NAND2_X2 U5112 ( .A1(w_q[83]), .A2(n7216), .ZN(n5872) );
NAND2_X2 U5113 ( .A1(w_q[115]), .A2(n7240), .ZN(n5871) );
NAND2_X2 U5114 ( .A1(n5873), .A2(n5874), .ZN(w_d[114]) );
NAND2_X2 U5115 ( .A1(w_q[82]), .A2(n7226), .ZN(n5874) );
NAND2_X2 U5116 ( .A1(w_q[114]), .A2(n7240), .ZN(n5873) );
NAND2_X2 U5117 ( .A1(n5875), .A2(n5876), .ZN(w_d[113]) );
NAND2_X2 U5118 ( .A1(w_q[81]), .A2(n7214), .ZN(n5876) );
NAND2_X2 U5119 ( .A1(w_q[113]), .A2(n7240), .ZN(n5875) );
NAND2_X2 U5120 ( .A1(n5877), .A2(n5878), .ZN(w_d[112]) );
NAND2_X2 U5121 ( .A1(w_q[80]), .A2(n7183), .ZN(n5878) );
NAND2_X2 U5122 ( .A1(w_q[112]), .A2(n7240), .ZN(n5877) );
NAND2_X2 U5123 ( .A1(n5879), .A2(n5880), .ZN(w_d[111]) );
NAND2_X2 U5124 ( .A1(w_q[79]), .A2(n7184), .ZN(n5880) );
NAND2_X2 U5125 ( .A1(w_q[111]), .A2(n7240), .ZN(n5879) );
NAND2_X2 U5126 ( .A1(n5881), .A2(n5882), .ZN(w_d[110]) );
NAND2_X2 U5127 ( .A1(w_q[78]), .A2(n7182), .ZN(n5882) );
NAND2_X2 U5128 ( .A1(w_q[110]), .A2(n7240), .ZN(n5881) );
NAND2_X2 U5130 ( .A1(w[10]), .A2(n7160), .ZN(n5885) );
NAND2_X2 U5131 ( .A1(w_q[10]), .A2(n7240), .ZN(n5884) );
NAND2_X2 U5133 ( .A1(n5886), .A2(n5887), .ZN(w_d[109]) );
NAND2_X2 U5134 ( .A1(w_q[77]), .A2(n7182), .ZN(n5887) );
NAND2_X2 U5135 ( .A1(w_q[109]), .A2(n7239), .ZN(n5886) );
NAND2_X2 U5136 ( .A1(n5888), .A2(n5889), .ZN(w_d[108]) );
NAND2_X2 U5137 ( .A1(w_q[76]), .A2(n7182), .ZN(n5889) );
NAND2_X2 U5138 ( .A1(w_q[108]), .A2(n7239), .ZN(n5888) );
NAND2_X2 U5139 ( .A1(n5890), .A2(n5891), .ZN(w_d[107]) );
NAND2_X2 U5140 ( .A1(w_q[75]), .A2(n7182), .ZN(n5891) );
NAND2_X2 U5141 ( .A1(w_q[107]), .A2(n7239), .ZN(n5890) );
NAND2_X2 U5142 ( .A1(n5892), .A2(n5893), .ZN(w_d[106]) );
NAND2_X2 U5143 ( .A1(w_q[74]), .A2(n7182), .ZN(n5893) );
NAND2_X2 U5144 ( .A1(w_q[106]), .A2(n7239), .ZN(n5892) );
NAND2_X2 U5145 ( .A1(n5894), .A2(n5895), .ZN(w_d[105]) );
NAND2_X2 U5146 ( .A1(w_q[73]), .A2(n7182), .ZN(n5895) );
NAND2_X2 U5147 ( .A1(w_q[105]), .A2(n7239), .ZN(n5894) );
NAND2_X2 U5148 ( .A1(n5896), .A2(n5897), .ZN(w_d[104]) );
NAND2_X2 U5149 ( .A1(w_q[72]), .A2(n7182), .ZN(n5897) );
NAND2_X2 U5150 ( .A1(w_q[104]), .A2(n7239), .ZN(n5896) );
NAND2_X2 U5151 ( .A1(n5898), .A2(n5899), .ZN(w_d[103]) );
NAND2_X2 U5152 ( .A1(w_q[71]), .A2(n7182), .ZN(n5899) );
NAND2_X2 U5153 ( .A1(w_q[103]), .A2(n7239), .ZN(n5898) );
NAND2_X2 U5154 ( .A1(n5900), .A2(n5901), .ZN(w_d[102]) );
NAND2_X2 U5155 ( .A1(w_q[70]), .A2(n7182), .ZN(n5901) );
NAND2_X2 U5156 ( .A1(w_q[102]), .A2(n7239), .ZN(n5900) );
NAND2_X2 U5157 ( .A1(n5902), .A2(n5903), .ZN(w_d[101]) );
NAND2_X2 U5158 ( .A1(w_q[69]), .A2(n7182), .ZN(n5903) );
NAND2_X2 U5159 ( .A1(w_q[101]), .A2(n7239), .ZN(n5902) );
NAND2_X2 U5160 ( .A1(n5904), .A2(n5905), .ZN(w_d[100]) );
NAND2_X2 U5161 ( .A1(w_q[68]), .A2(n7182), .ZN(n5905) );
NAND2_X2 U5163 ( .A1(w_q[100]), .A2(n7239), .ZN(n5904) );
NAND2_X2 U5165 ( .A1(w[0]), .A2(n7160), .ZN(n5908) );
NAND2_X2 U5166 ( .A1(w_q[0]), .A2(n7239), .ZN(n5907) );
NAND2_X2 U5170 ( .A1(n5909), .A2(n5910), .ZN(rnd_d[9]) );
NAND2_X2 U5171 ( .A1(sha1_round_wire[9]), .A2(n7160), .ZN(n5910) );
NAND2_X2 U5172 ( .A1(n5911), .A2(n5912), .ZN(rnd_d[99]) );
NAND2_X2 U5173 ( .A1(sha1_round_wire[99]), .A2(n7160), .ZN(n5912) );
NAND2_X2 U5174 ( .A1(n5913), .A2(n5914), .ZN(rnd_d[98]) );
NAND2_X2 U5175 ( .A1(sha1_round_wire[98]), .A2(n7160), .ZN(n5914) );
NAND2_X2 U5176 ( .A1(n5915), .A2(n5916), .ZN(rnd_d[97]) );
NAND2_X2 U5177 ( .A1(sha1_round_wire[97]), .A2(n7160), .ZN(n5916) );
NAND2_X2 U5178 ( .A1(n5917), .A2(n5918), .ZN(rnd_d[96]) );
NAND2_X2 U5179 ( .A1(sha1_round_wire[96]), .A2(n7160), .ZN(n5918) );
NAND2_X2 U5180 ( .A1(n5919), .A2(n5920), .ZN(rnd_d[95]) );
NAND2_X2 U5181 ( .A1(sha1_round_wire[95]), .A2(n7160), .ZN(n5920) );
NAND2_X2 U5182 ( .A1(n5921), .A2(n5922), .ZN(rnd_d[94]) );
NAND2_X2 U5183 ( .A1(sha1_round_wire[94]), .A2(n7160), .ZN(n5922) );
NAND2_X2 U5184 ( .A1(n5923), .A2(n5924), .ZN(rnd_d[93]) );
NAND2_X2 U5185 ( .A1(sha1_round_wire[93]), .A2(n7160), .ZN(n5924) );
NAND2_X2 U5186 ( .A1(n5925), .A2(n5926), .ZN(rnd_d[92]) );
NAND2_X2 U5187 ( .A1(sha1_round_wire[92]), .A2(n7161), .ZN(n5926) );
NAND2_X2 U5188 ( .A1(n5927), .A2(n5928), .ZN(rnd_d[91]) );
NAND2_X2 U5189 ( .A1(sha1_round_wire[91]), .A2(n7161), .ZN(n5928) );
NAND2_X2 U5190 ( .A1(n5929), .A2(n5930), .ZN(rnd_d[90]) );
NAND2_X2 U5191 ( .A1(sha1_round_wire[90]), .A2(n7161), .ZN(n5930) );
NAND2_X2 U5192 ( .A1(n5931), .A2(n5932), .ZN(rnd_d[8]) );
NAND2_X2 U5193 ( .A1(sha1_round_wire[8]), .A2(n7161), .ZN(n5932) );
NAND2_X2 U5194 ( .A1(n5933), .A2(n5934), .ZN(rnd_d[89]) );
NAND2_X2 U5195 ( .A1(sha1_round_wire[89]), .A2(n7161), .ZN(n5934) );
NAND2_X2 U5196 ( .A1(n5935), .A2(n5936), .ZN(rnd_d[88]) );
NAND2_X2 U5197 ( .A1(sha1_round_wire[88]), .A2(n7161), .ZN(n5936) );
NAND2_X2 U5198 ( .A1(n5937), .A2(n5938), .ZN(rnd_d[87]) );
NAND2_X2 U5199 ( .A1(sha1_round_wire[87]), .A2(n7161), .ZN(n5938) );
NAND2_X2 U5200 ( .A1(n5939), .A2(n5940), .ZN(rnd_d[86]) );
NAND2_X2 U5201 ( .A1(sha1_round_wire[86]), .A2(n7161), .ZN(n5940) );
NAND2_X2 U5202 ( .A1(n5941), .A2(n5942), .ZN(rnd_d[85]) );
NAND2_X2 U5203 ( .A1(sha1_round_wire[85]), .A2(n7161), .ZN(n5942) );
NAND2_X2 U5204 ( .A1(n5943), .A2(n5944), .ZN(rnd_d[84]) );
NAND2_X2 U5205 ( .A1(sha1_round_wire[84]), .A2(n7161), .ZN(n5944) );
NAND2_X2 U5206 ( .A1(n5945), .A2(n5946), .ZN(rnd_d[83]) );
NAND2_X2 U5207 ( .A1(sha1_round_wire[83]), .A2(n7161), .ZN(n5946) );
NAND2_X2 U5208 ( .A1(n5947), .A2(n5948), .ZN(rnd_d[82]) );
NAND2_X2 U5209 ( .A1(sha1_round_wire[82]), .A2(n7161), .ZN(n5948) );
NAND2_X2 U5210 ( .A1(n5949), .A2(n5950), .ZN(rnd_d[81]) );
NAND2_X2 U5211 ( .A1(sha1_round_wire[81]), .A2(n7161), .ZN(n5950) );
NAND2_X2 U5212 ( .A1(n5951), .A2(n5952), .ZN(rnd_d[80]) );
NAND2_X2 U5213 ( .A1(sha1_round_wire[80]), .A2(n7161), .ZN(n5952) );
NAND2_X2 U5214 ( .A1(n5953), .A2(n5954), .ZN(rnd_d[7]) );
NAND2_X2 U5215 ( .A1(sha1_round_wire[7]), .A2(n7161), .ZN(n5954) );
NAND2_X2 U5216 ( .A1(n5955), .A2(n5956), .ZN(rnd_d[79]) );
NAND2_X2 U5217 ( .A1(sha1_round_wire[79]), .A2(n7161), .ZN(n5956) );
NAND2_X2 U5218 ( .A1(n5957), .A2(n5958), .ZN(rnd_d[78]) );
NAND2_X2 U5219 ( .A1(sha1_round_wire[78]), .A2(n7161), .ZN(n5958) );
NAND2_X2 U5220 ( .A1(n5959), .A2(n5960), .ZN(rnd_d[77]) );
NAND2_X2 U5221 ( .A1(sha1_round_wire[77]), .A2(n7161), .ZN(n5960) );
NAND2_X2 U5222 ( .A1(n5961), .A2(n5962), .ZN(rnd_d[76]) );
NAND2_X2 U5223 ( .A1(sha1_round_wire[76]), .A2(n7161), .ZN(n5962) );
NAND2_X2 U5224 ( .A1(n5963), .A2(n5964), .ZN(rnd_d[75]) );
NAND2_X2 U5225 ( .A1(sha1_round_wire[75]), .A2(n7161), .ZN(n5964) );
NAND2_X2 U5226 ( .A1(n5965), .A2(n5966), .ZN(rnd_d[74]) );
NAND2_X2 U5227 ( .A1(sha1_round_wire[74]), .A2(n7161), .ZN(n5966) );
NAND2_X2 U5228 ( .A1(n5967), .A2(n5968), .ZN(rnd_d[73]) );
NAND2_X2 U5229 ( .A1(sha1_round_wire[73]), .A2(n7161), .ZN(n5968) );
NAND2_X2 U5230 ( .A1(n5969), .A2(n5970), .ZN(rnd_d[72]) );
NAND2_X2 U5231 ( .A1(sha1_round_wire[72]), .A2(n7161), .ZN(n5970) );
NAND2_X2 U5232 ( .A1(n5971), .A2(n5972), .ZN(rnd_d[71]) );
NAND2_X2 U5233 ( .A1(sha1_round_wire[71]), .A2(n7161), .ZN(n5972) );
NAND2_X2 U5234 ( .A1(n5973), .A2(n5974), .ZN(rnd_d[70]) );
NAND2_X2 U5235 ( .A1(sha1_round_wire[70]), .A2(n7161), .ZN(n5974) );
NAND2_X2 U5236 ( .A1(n5975), .A2(n5976), .ZN(rnd_d[6]) );
NAND2_X2 U5237 ( .A1(sha1_round_wire[6]), .A2(n7161), .ZN(n5976) );
NAND2_X2 U5238 ( .A1(n5977), .A2(n5978), .ZN(rnd_d[69]) );
NAND2_X2 U5239 ( .A1(sha1_round_wire[69]), .A2(n7161), .ZN(n5978) );
NAND2_X2 U5240 ( .A1(n5979), .A2(n5980), .ZN(rnd_d[68]) );
NAND2_X2 U5241 ( .A1(sha1_round_wire[68]), .A2(n7162), .ZN(n5980) );
NAND2_X2 U5242 ( .A1(n5981), .A2(n5982), .ZN(rnd_d[67]) );
NAND2_X2 U5243 ( .A1(sha1_round_wire[67]), .A2(n7162), .ZN(n5982) );
NAND2_X2 U5244 ( .A1(n5983), .A2(n5984), .ZN(rnd_d[66]) );
NAND2_X2 U5245 ( .A1(sha1_round_wire[66]), .A2(n7162), .ZN(n5984) );
NAND2_X2 U5246 ( .A1(n5985), .A2(n5986), .ZN(rnd_d[65]) );
NAND2_X2 U5247 ( .A1(sha1_round_wire[65]), .A2(n7162), .ZN(n5986) );
NAND2_X2 U5248 ( .A1(n5987), .A2(n5988), .ZN(rnd_d[64]) );
NAND2_X2 U5249 ( .A1(sha1_round_wire[64]), .A2(n7162), .ZN(n5988) );
NAND2_X2 U5250 ( .A1(n5989), .A2(n5990), .ZN(rnd_d[63]) );
NAND2_X2 U5251 ( .A1(sha1_round_wire[63]), .A2(n7162), .ZN(n5990) );
NAND2_X2 U5252 ( .A1(n5991), .A2(n5992), .ZN(rnd_d[62]) );
NAND2_X2 U5253 ( .A1(sha1_round_wire[62]), .A2(n7162), .ZN(n5992) );
NAND2_X2 U5254 ( .A1(n5993), .A2(n5994), .ZN(rnd_d[61]) );
NAND2_X2 U5255 ( .A1(sha1_round_wire[61]), .A2(n7162), .ZN(n5994) );
NAND2_X2 U5256 ( .A1(n5995), .A2(n5996), .ZN(rnd_d[60]) );
NAND2_X2 U5257 ( .A1(sha1_round_wire[60]), .A2(n7162), .ZN(n5996) );
NAND2_X2 U5258 ( .A1(n5997), .A2(n5998), .ZN(rnd_d[5]) );
NAND2_X2 U5259 ( .A1(sha1_round_wire[5]), .A2(n7162), .ZN(n5998) );
NAND2_X2 U5260 ( .A1(n5999), .A2(n6000), .ZN(rnd_d[59]) );
NAND2_X2 U5261 ( .A1(sha1_round_wire[59]), .A2(n7162), .ZN(n6000) );
NAND2_X2 U5262 ( .A1(n6001), .A2(n6002), .ZN(rnd_d[58]) );
NAND2_X2 U5263 ( .A1(sha1_round_wire[58]), .A2(n7162), .ZN(n6002) );
NAND2_X2 U5264 ( .A1(n6003), .A2(n6004), .ZN(rnd_d[57]) );
NAND2_X2 U5265 ( .A1(sha1_round_wire[57]), .A2(n7162), .ZN(n6004) );
NAND2_X2 U5266 ( .A1(n6005), .A2(n6006), .ZN(rnd_d[56]) );
NAND2_X2 U5267 ( .A1(sha1_round_wire[56]), .A2(n7162), .ZN(n6006) );
NAND2_X2 U5268 ( .A1(n6007), .A2(n6008), .ZN(rnd_d[55]) );
NAND2_X2 U5269 ( .A1(sha1_round_wire[55]), .A2(n7162), .ZN(n6008) );
NAND2_X2 U5270 ( .A1(n6009), .A2(n6010), .ZN(rnd_d[54]) );
NAND2_X2 U5271 ( .A1(sha1_round_wire[54]), .A2(n7162), .ZN(n6010) );
NAND2_X2 U5272 ( .A1(n6011), .A2(n6012), .ZN(rnd_d[53]) );
NAND2_X2 U5273 ( .A1(sha1_round_wire[53]), .A2(n7162), .ZN(n6012) );
NAND2_X2 U5274 ( .A1(n6013), .A2(n6014), .ZN(rnd_d[52]) );
NAND2_X2 U5275 ( .A1(sha1_round_wire[52]), .A2(n7162), .ZN(n6014) );
NAND2_X2 U5276 ( .A1(n6015), .A2(n6016), .ZN(rnd_d[51]) );
NAND2_X2 U5277 ( .A1(sha1_round_wire[51]), .A2(n7162), .ZN(n6016) );
NAND2_X2 U5278 ( .A1(n6017), .A2(n6018), .ZN(rnd_d[50]) );
NAND2_X2 U5279 ( .A1(sha1_round_wire[50]), .A2(n7162), .ZN(n6018) );
NAND2_X2 U5280 ( .A1(n6019), .A2(n6020), .ZN(rnd_d[4]) );
NAND2_X2 U5281 ( .A1(sha1_round_wire[4]), .A2(n7162), .ZN(n6020) );
NAND2_X2 U5282 ( .A1(n6021), .A2(n6022), .ZN(rnd_d[49]) );
NAND2_X2 U5283 ( .A1(sha1_round_wire[49]), .A2(n7162), .ZN(n6022) );
NAND2_X2 U5284 ( .A1(n6023), .A2(n6024), .ZN(rnd_d[48]) );
NAND2_X2 U5285 ( .A1(sha1_round_wire[48]), .A2(n7162), .ZN(n6024) );
NAND2_X2 U5286 ( .A1(n6025), .A2(n6026), .ZN(rnd_d[47]) );
NAND2_X2 U5287 ( .A1(sha1_round_wire[47]), .A2(n7162), .ZN(n6026) );
NAND2_X2 U5288 ( .A1(n6027), .A2(n6028), .ZN(rnd_d[46]) );
NAND2_X2 U5289 ( .A1(sha1_round_wire[46]), .A2(n7162), .ZN(n6028) );
NAND2_X2 U5290 ( .A1(n6029), .A2(n6030), .ZN(rnd_d[45]) );
NAND2_X2 U5291 ( .A1(sha1_round_wire[45]), .A2(n7162), .ZN(n6030) );
NAND2_X2 U5292 ( .A1(n6031), .A2(n6032), .ZN(rnd_d[44]) );
NAND2_X2 U5293 ( .A1(sha1_round_wire[44]), .A2(n7163), .ZN(n6032) );
NAND2_X2 U5294 ( .A1(n6033), .A2(n6034), .ZN(rnd_d[43]) );
NAND2_X2 U5295 ( .A1(sha1_round_wire[43]), .A2(n7163), .ZN(n6034) );
NAND2_X2 U5296 ( .A1(n6035), .A2(n6036), .ZN(rnd_d[42]) );
NAND2_X2 U5297 ( .A1(sha1_round_wire[42]), .A2(n7163), .ZN(n6036) );
NAND2_X2 U5298 ( .A1(n6037), .A2(n6038), .ZN(rnd_d[41]) );
NAND2_X2 U5299 ( .A1(sha1_round_wire[41]), .A2(n7163), .ZN(n6038) );
NAND2_X2 U5300 ( .A1(n6039), .A2(n6040), .ZN(rnd_d[40]) );
NAND2_X2 U5301 ( .A1(sha1_round_wire[40]), .A2(n7163), .ZN(n6040) );
NAND2_X2 U5302 ( .A1(n6041), .A2(n6042), .ZN(rnd_d[3]) );
NAND2_X2 U5303 ( .A1(sha1_round_wire[3]), .A2(n7163), .ZN(n6042) );
NAND2_X2 U5304 ( .A1(n6043), .A2(n6044), .ZN(rnd_d[39]) );
NAND2_X2 U5305 ( .A1(sha1_round_wire[39]), .A2(n7163), .ZN(n6044) );
NAND2_X2 U5306 ( .A1(n6045), .A2(n6046), .ZN(rnd_d[38]) );
NAND2_X2 U5307 ( .A1(sha1_round_wire[38]), .A2(n7163), .ZN(n6046) );
NAND2_X2 U5308 ( .A1(n6047), .A2(n6048), .ZN(rnd_d[37]) );
NAND2_X2 U5309 ( .A1(sha1_round_wire[37]), .A2(n7163), .ZN(n6048) );
NAND2_X2 U5310 ( .A1(n6049), .A2(n6050), .ZN(rnd_d[36]) );
NAND2_X2 U5311 ( .A1(sha1_round_wire[36]), .A2(n7163), .ZN(n6050) );
NAND2_X2 U5312 ( .A1(n6051), .A2(n6052), .ZN(rnd_d[35]) );
NAND2_X2 U5313 ( .A1(sha1_round_wire[35]), .A2(n7163), .ZN(n6052) );
NAND2_X2 U5314 ( .A1(n6053), .A2(n6054), .ZN(rnd_d[34]) );
NAND2_X2 U5315 ( .A1(sha1_round_wire[34]), .A2(n7163), .ZN(n6054) );
NAND2_X2 U5316 ( .A1(n6055), .A2(n6056), .ZN(rnd_d[33]) );
NAND2_X2 U5317 ( .A1(sha1_round_wire[33]), .A2(n7163), .ZN(n6056) );
NAND2_X2 U5318 ( .A1(n6057), .A2(n6058), .ZN(rnd_d[32]) );
NAND2_X2 U5319 ( .A1(sha1_round_wire[32]), .A2(n7163), .ZN(n6058) );
NAND2_X2 U5320 ( .A1(n6059), .A2(n6060), .ZN(rnd_d[31]) );
NAND2_X2 U5321 ( .A1(sha1_round_wire[31]), .A2(n7163), .ZN(n6060) );
NAND2_X2 U5322 ( .A1(n6061), .A2(n6062), .ZN(rnd_d[30]) );
NAND2_X2 U5323 ( .A1(sha1_round_wire[30]), .A2(n7163), .ZN(n6062) );
NAND2_X2 U5324 ( .A1(n6063), .A2(n6064), .ZN(rnd_d[2]) );
NAND2_X2 U5325 ( .A1(sha1_round_wire[2]), .A2(n7163), .ZN(n6064) );
NAND2_X2 U5326 ( .A1(n6065), .A2(n6066), .ZN(rnd_d[29]) );
NAND2_X2 U5327 ( .A1(sha1_round_wire[29]), .A2(n7163), .ZN(n6066) );
NAND2_X2 U5328 ( .A1(n6067), .A2(n6068), .ZN(rnd_d[28]) );
NAND2_X2 U5329 ( .A1(sha1_round_wire[28]), .A2(n7163), .ZN(n6068) );
NAND2_X2 U5330 ( .A1(n6069), .A2(n6070), .ZN(rnd_d[27]) );
NAND2_X2 U5331 ( .A1(sha1_round_wire[27]), .A2(n7163), .ZN(n6070) );
NAND2_X2 U5332 ( .A1(n6071), .A2(n6072), .ZN(rnd_d[26]) );
NAND2_X2 U5333 ( .A1(sha1_round_wire[26]), .A2(n7163), .ZN(n6072) );
NAND2_X2 U5334 ( .A1(n6073), .A2(n6074), .ZN(rnd_d[25]) );
NAND2_X2 U5335 ( .A1(sha1_round_wire[25]), .A2(n7163), .ZN(n6074) );
NAND2_X2 U5336 ( .A1(n6075), .A2(n6076), .ZN(rnd_d[24]) );
NAND2_X2 U5337 ( .A1(sha1_round_wire[24]), .A2(n7163), .ZN(n6076) );
NAND2_X2 U5338 ( .A1(n6077), .A2(n6078), .ZN(rnd_d[23]) );
NAND2_X2 U5339 ( .A1(sha1_round_wire[23]), .A2(n7163), .ZN(n6078) );
NAND2_X2 U5340 ( .A1(n6079), .A2(n6080), .ZN(rnd_d[22]) );
NAND2_X2 U5341 ( .A1(sha1_round_wire[22]), .A2(n7163), .ZN(n6080) );
NAND2_X2 U5342 ( .A1(n6081), .A2(n6082), .ZN(rnd_d[21]) );
NAND2_X2 U5343 ( .A1(sha1_round_wire[21]), .A2(n7163), .ZN(n6082) );
NAND2_X2 U5344 ( .A1(n6083), .A2(n6084), .ZN(rnd_d[20]) );
NAND2_X2 U5345 ( .A1(sha1_round_wire[20]), .A2(n7163), .ZN(n6084) );
NAND2_X2 U5346 ( .A1(n6085), .A2(n6086), .ZN(rnd_d[1]) );
NAND2_X2 U5347 ( .A1(sha1_round_wire[1]), .A2(n7164), .ZN(n6086) );
NAND2_X2 U5348 ( .A1(n6087), .A2(n6088), .ZN(rnd_d[19]) );
NAND2_X2 U5349 ( .A1(sha1_round_wire[19]), .A2(n7164), .ZN(n6088) );
NAND2_X2 U5350 ( .A1(n6089), .A2(n6090), .ZN(rnd_d[18]) );
NAND2_X2 U5351 ( .A1(sha1_round_wire[18]), .A2(n7164), .ZN(n6090) );
NAND2_X2 U5352 ( .A1(n6091), .A2(n6092), .ZN(rnd_d[17]) );
NAND2_X2 U5353 ( .A1(sha1_round_wire[17]), .A2(n7164), .ZN(n6092) );
NAND2_X2 U5354 ( .A1(n6093), .A2(n6094), .ZN(rnd_d[16]) );
NAND2_X2 U5355 ( .A1(sha1_round_wire[16]), .A2(n7164), .ZN(n6094) );
NAND2_X2 U5356 ( .A1(n6095), .A2(n6096), .ZN(rnd_d[15]) );
NAND2_X2 U5357 ( .A1(sha1_round_wire[15]), .A2(n7164), .ZN(n6096) );
NAND2_X2 U5378 ( .A1(n6117), .A2(n6118), .ZN(rnd_d[14]) );
NAND2_X2 U5379 ( .A1(sha1_round_wire[14]), .A2(n7164), .ZN(n6118) );
NAND2_X2 U5400 ( .A1(n6139), .A2(n6140), .ZN(rnd_d[13]) );
NAND2_X2 U5401 ( .A1(sha1_round_wire[13]), .A2(n7164), .ZN(n6140) );
NAND2_X2 U5406 ( .A1(n6145), .A2(n6146), .ZN(rnd_d[137]) );
NAND2_X2 U5407 ( .A1(sha1_round_wire[137]), .A2(n7164), .ZN(n6146) );
NAND2_X2 U5408 ( .A1(n6147), .A2(n6148), .ZN(rnd_d[136]) );
NAND2_X2 U5409 ( .A1(sha1_round_wire[136]), .A2(n7164), .ZN(n6148) );
NAND2_X2 U5410 ( .A1(n6149), .A2(n6150), .ZN(rnd_d[135]) );
NAND2_X2 U5411 ( .A1(sha1_round_wire[135]), .A2(n7164), .ZN(n6150) );
NAND2_X2 U5412 ( .A1(n6151), .A2(n6152), .ZN(rnd_d[134]) );
NAND2_X2 U5413 ( .A1(sha1_round_wire[134]), .A2(n7164), .ZN(n6152) );
NAND2_X2 U5414 ( .A1(n6153), .A2(n6154), .ZN(rnd_d[133]) );
NAND2_X2 U5415 ( .A1(sha1_round_wire[133]), .A2(n7164), .ZN(n6154) );
NAND2_X2 U5416 ( .A1(n6155), .A2(n6156), .ZN(rnd_d[132]) );
NAND2_X2 U5417 ( .A1(sha1_round_wire[132]), .A2(n7164), .ZN(n6156) );
NAND2_X2 U5418 ( .A1(n6157), .A2(n6158), .ZN(rnd_d[131]) );
NAND2_X2 U5419 ( .A1(sha1_round_wire[131]), .A2(n7164), .ZN(n6158) );
NAND2_X2 U5420 ( .A1(n6159), .A2(n6160), .ZN(rnd_d[130]) );
NAND2_X2 U5421 ( .A1(sha1_round_wire[130]), .A2(n7164), .ZN(n6160) );
NAND2_X2 U5422 ( .A1(n6161), .A2(n6162), .ZN(rnd_d[12]) );
NAND2_X2 U5423 ( .A1(sha1_round_wire[12]), .A2(n7164), .ZN(n6162) );
NAND2_X2 U5424 ( .A1(n6163), .A2(n6164), .ZN(rnd_d[129]) );
NAND2_X2 U5425 ( .A1(sha1_round_wire[129]), .A2(n7164), .ZN(n6164) );
NAND2_X2 U5426 ( .A1(n6165), .A2(n6166), .ZN(rnd_d[128]) );
NAND2_X2 U5427 ( .A1(sha1_round_wire[128]), .A2(n7164), .ZN(n6166) );
NAND2_X2 U5428 ( .A1(n6167), .A2(n6168), .ZN(rnd_d[127]) );
NAND2_X2 U5429 ( .A1(sha1_round_wire[127]), .A2(n7164), .ZN(n6168) );
NAND2_X2 U5430 ( .A1(n6169), .A2(n6170), .ZN(rnd_d[126]) );
NAND2_X2 U5431 ( .A1(sha1_round_wire[126]), .A2(n7164), .ZN(n6170) );
NAND2_X2 U5432 ( .A1(n6171), .A2(n6172), .ZN(rnd_d[125]) );
NAND2_X2 U5433 ( .A1(sha1_round_wire[125]), .A2(n7164), .ZN(n6172) );
NAND2_X2 U5434 ( .A1(n6173), .A2(n6174), .ZN(rnd_d[124]) );
NAND2_X2 U5435 ( .A1(sha1_round_wire[124]), .A2(n7164), .ZN(n6174) );
NAND2_X2 U5436 ( .A1(n6175), .A2(n6176), .ZN(rnd_d[123]) );
NAND2_X2 U5437 ( .A1(sha1_round_wire[123]), .A2(n7164), .ZN(n6176) );
NAND2_X2 U5438 ( .A1(n6177), .A2(n6178), .ZN(rnd_d[122]) );
NAND2_X2 U5439 ( .A1(sha1_round_wire[122]), .A2(n7164), .ZN(n6178) );
NAND2_X2 U5440 ( .A1(n6179), .A2(n6180), .ZN(rnd_d[121]) );
NAND2_X2 U5441 ( .A1(sha1_round_wire[121]), .A2(n7164), .ZN(n6180) );
NAND2_X2 U5442 ( .A1(n6181), .A2(n6182), .ZN(rnd_d[120]) );
NAND2_X2 U5443 ( .A1(sha1_round_wire[120]), .A2(n7164), .ZN(n6182) );
NAND2_X2 U5444 ( .A1(n6183), .A2(n6184), .ZN(rnd_d[11]) );
NAND2_X2 U5445 ( .A1(sha1_round_wire[11]), .A2(n7165), .ZN(n6184) );
NAND2_X2 U5446 ( .A1(n6185), .A2(n6186), .ZN(rnd_d[119]) );
NAND2_X2 U5447 ( .A1(sha1_round_wire[119]), .A2(n7165), .ZN(n6186) );
NAND2_X2 U5448 ( .A1(n6187), .A2(n6188), .ZN(rnd_d[118]) );
NAND2_X2 U5449 ( .A1(sha1_round_wire[118]), .A2(n7165), .ZN(n6188) );
NAND2_X2 U5450 ( .A1(n6189), .A2(n6190), .ZN(rnd_d[117]) );
NAND2_X2 U5451 ( .A1(sha1_round_wire[117]), .A2(n7165), .ZN(n6190) );
NAND2_X2 U5452 ( .A1(n6191), .A2(n6192), .ZN(rnd_d[116]) );
NAND2_X2 U5453 ( .A1(sha1_round_wire[116]), .A2(n7165), .ZN(n6192) );
NAND2_X2 U5454 ( .A1(n6193), .A2(n6194), .ZN(rnd_d[115]) );
NAND2_X2 U5455 ( .A1(sha1_round_wire[115]), .A2(n7165), .ZN(n6194) );
NAND2_X2 U5456 ( .A1(n6195), .A2(n6196), .ZN(rnd_d[114]) );
NAND2_X2 U5457 ( .A1(sha1_round_wire[114]), .A2(n7165), .ZN(n6196) );
NAND2_X2 U5458 ( .A1(n6197), .A2(n6198), .ZN(rnd_d[113]) );
NAND2_X2 U5459 ( .A1(sha1_round_wire[113]), .A2(n7155), .ZN(n6198) );
NAND2_X2 U5460 ( .A1(n6199), .A2(n6200), .ZN(rnd_d[112]) );
NAND2_X2 U5461 ( .A1(sha1_round_wire[112]), .A2(n7152), .ZN(n6200) );
NAND2_X2 U5462 ( .A1(n6201), .A2(n6202), .ZN(rnd_d[111]) );
NAND2_X2 U5463 ( .A1(sha1_round_wire[111]), .A2(n7152), .ZN(n6202) );
NAND2_X2 U5464 ( .A1(n6203), .A2(n6204), .ZN(rnd_d[110]) );
NAND2_X2 U5465 ( .A1(sha1_round_wire[110]), .A2(n7152), .ZN(n6204) );
NAND2_X2 U5466 ( .A1(n6205), .A2(n6206), .ZN(rnd_d[10]) );
NAND2_X2 U5467 ( .A1(sha1_round_wire[10]), .A2(n7152), .ZN(n6206) );
NAND2_X2 U5468 ( .A1(n6207), .A2(n6208), .ZN(rnd_d[109]) );
NAND2_X2 U5469 ( .A1(sha1_round_wire[109]), .A2(n7152), .ZN(n6208) );
NAND2_X2 U5470 ( .A1(n6209), .A2(n6210), .ZN(rnd_d[108]) );
NAND2_X2 U5471 ( .A1(sha1_round_wire[108]), .A2(n7152), .ZN(n6210) );
NAND2_X2 U5472 ( .A1(n6211), .A2(n6212), .ZN(rnd_d[107]) );
NAND2_X2 U5473 ( .A1(sha1_round_wire[107]), .A2(n7152), .ZN(n6212) );
NAND2_X2 U5474 ( .A1(n6213), .A2(n6214), .ZN(rnd_d[106]) );
NAND2_X2 U5475 ( .A1(sha1_round_wire[106]), .A2(n7152), .ZN(n6214) );
NAND2_X2 U5476 ( .A1(n6215), .A2(n6216), .ZN(rnd_d[105]) );
NAND2_X2 U5477 ( .A1(sha1_round_wire[105]), .A2(n7152), .ZN(n6216) );
NAND2_X2 U5478 ( .A1(n6217), .A2(n6218), .ZN(rnd_d[104]) );
NAND2_X2 U5479 ( .A1(sha1_round_wire[104]), .A2(n7152), .ZN(n6218) );
NAND2_X2 U5480 ( .A1(n6219), .A2(n6220), .ZN(rnd_d[103]) );
NAND2_X2 U5481 ( .A1(sha1_round_wire[103]), .A2(n7152), .ZN(n6220) );
NAND2_X2 U5482 ( .A1(n6221), .A2(n6222), .ZN(rnd_d[102]) );
NAND2_X2 U5483 ( .A1(sha1_round_wire[102]), .A2(n7152), .ZN(n6222) );
NAND2_X2 U5484 ( .A1(n6223), .A2(n6224), .ZN(rnd_d[101]) );
NAND2_X2 U5485 ( .A1(sha1_round_wire[101]), .A2(n7152), .ZN(n6224) );
NAND2_X2 U5486 ( .A1(n6225), .A2(n6226), .ZN(rnd_d[100]) );
NAND2_X2 U5487 ( .A1(sha1_round_wire[100]), .A2(n7152), .ZN(n6226) );
NAND2_X2 U5488 ( .A1(n6227), .A2(n6228), .ZN(rnd_d[0]) );
NAND2_X2 U5489 ( .A1(sha1_round_wire[0]), .A2(n7152), .ZN(n6228) );
XNOR2_X2 U5494 ( .A(n6232), .B(n7398), .ZN(n6233) );
NAND2_X2 U5500 ( .A1(n6237), .A2(n6238), .ZN(rnd_cnt_d[2]) );
NAND4_X2 U5501 ( .A1(n7396), .A2(rnd_cnt_q[1]), .A3(rnd_cnt_q[0]), .A4(n7400), .ZN(n6238) );
NAND2_X2 U5503 ( .A1(n7397), .A2(n6240), .ZN(n6239) );
NAND2_X2 U5504 ( .A1(n7396), .A2(n7401), .ZN(n6240) );
NAND2_X2 U5505 ( .A1(n6241), .A2(n6242), .ZN(rnd_cnt_d[1]) );
NAND2_X2 U5507 ( .A1(rnd_cnt_d[0]), .A2(rnd_cnt_q[1]), .ZN(n6241) );
AND2_X2 U5509 ( .A1(state[0]), .A2(state[1]), .ZN(out_valid) );
NAND2_X2 U5514 ( .A1(n7176), .A2(n7402), .ZN(n6247) );
AND2_X2 U5517 ( .A1(rnd_cnt_q[3]), .A2(n6236), .ZN(n5038) );
NAND2_X2 U6001 ( .A1(n5909), .A2(n6569), .ZN(cv_d[9]) );
NAND2_X2 U6002 ( .A1(cv_q[9]), .A2(n7152), .ZN(n6569) );
NAND2_X2 U6004 ( .A1(cv[9]), .A2(n7124), .ZN(n6571) );
NAND2_X2 U6005 ( .A1(cv_next[9]), .A2(n7139), .ZN(n6570) );
NAND2_X2 U6006 ( .A1(n5911), .A2(n6574), .ZN(cv_d[99]) );
NAND2_X2 U6007 ( .A1(cv_q[99]), .A2(n7152), .ZN(n6574) );
NAND2_X2 U6009 ( .A1(cv[99]), .A2(n7124), .ZN(n6576) );
NAND2_X2 U6010 ( .A1(cv_next[99]), .A2(n7139), .ZN(n6575) );
NAND2_X2 U6011 ( .A1(n5913), .A2(n6577), .ZN(cv_d[98]) );
NAND2_X2 U6012 ( .A1(cv_q[98]), .A2(n7152), .ZN(n6577) );
NAND2_X2 U6014 ( .A1(cv[98]), .A2(n7124), .ZN(n6579) );
NAND2_X2 U6015 ( .A1(cv_next[98]), .A2(n7139), .ZN(n6578) );
NAND2_X2 U6016 ( .A1(n5915), .A2(n6580), .ZN(cv_d[97]) );
NAND2_X2 U6017 ( .A1(cv_q[97]), .A2(n7153), .ZN(n6580) );
NAND2_X2 U6019 ( .A1(cv[97]), .A2(n7124), .ZN(n6582) );
NAND2_X2 U6020 ( .A1(cv_next[97]), .A2(n7139), .ZN(n6581) );
NAND2_X2 U6021 ( .A1(n5917), .A2(n6583), .ZN(cv_d[96]) );
NAND2_X2 U6022 ( .A1(cv_q[96]), .A2(n7152), .ZN(n6583) );
NAND2_X2 U6024 ( .A1(cv[96]), .A2(n7124), .ZN(n6585) );
NAND2_X2 U6025 ( .A1(cv_next[96]), .A2(n7139), .ZN(n6584) );
NAND2_X2 U6026 ( .A1(n5919), .A2(n6586), .ZN(cv_d[95]) );
NAND2_X2 U6027 ( .A1(cv_q[95]), .A2(n7152), .ZN(n6586) );
NAND2_X2 U6029 ( .A1(cv[95]), .A2(n7124), .ZN(n6588) );
NAND2_X2 U6030 ( .A1(cv_next[95]), .A2(n7139), .ZN(n6587) );
NAND2_X2 U6031 ( .A1(n5921), .A2(n6589), .ZN(cv_d[94]) );
NAND2_X2 U6032 ( .A1(cv_q[94]), .A2(n7153), .ZN(n6589) );
NAND2_X2 U6034 ( .A1(cv[94]), .A2(n7124), .ZN(n6591) );
NAND2_X2 U6035 ( .A1(cv_next[94]), .A2(n7139), .ZN(n6590) );
NAND2_X2 U6036 ( .A1(n5923), .A2(n6592), .ZN(cv_d[93]) );
NAND2_X2 U6037 ( .A1(cv_q[93]), .A2(n7153), .ZN(n6592) );
NAND2_X2 U6039 ( .A1(cv[93]), .A2(n7124), .ZN(n6594) );
NAND2_X2 U6040 ( .A1(cv_next[93]), .A2(n7139), .ZN(n6593) );
NAND2_X2 U6041 ( .A1(n5925), .A2(n6595), .ZN(cv_d[92]) );
NAND2_X2 U6042 ( .A1(cv_q[92]), .A2(n7153), .ZN(n6595) );
NAND2_X2 U6044 ( .A1(cv[92]), .A2(n7124), .ZN(n6597) );
NAND2_X2 U6045 ( .A1(cv_next[92]), .A2(n7139), .ZN(n6596) );
NAND2_X2 U6046 ( .A1(n5927), .A2(n6598), .ZN(cv_d[91]) );
NAND2_X2 U6047 ( .A1(cv_q[91]), .A2(n7153), .ZN(n6598) );
NAND2_X2 U6049 ( .A1(cv[91]), .A2(n7124), .ZN(n6600) );
NAND2_X2 U6050 ( .A1(cv_next[91]), .A2(n7139), .ZN(n6599) );
NAND2_X2 U6051 ( .A1(n5929), .A2(n6601), .ZN(cv_d[90]) );
NAND2_X2 U6052 ( .A1(cv_q[90]), .A2(n7153), .ZN(n6601) );
NAND2_X2 U6054 ( .A1(cv[90]), .A2(n7124), .ZN(n6603) );
NAND2_X2 U6055 ( .A1(cv_next[90]), .A2(n7139), .ZN(n6602) );
NAND2_X2 U6056 ( .A1(n5931), .A2(n6604), .ZN(cv_d[8]) );
NAND2_X2 U6057 ( .A1(cv_q[8]), .A2(n7153), .ZN(n6604) );
NAND2_X2 U6059 ( .A1(cv[8]), .A2(n7125), .ZN(n6606) );
NAND2_X2 U6060 ( .A1(cv_next[8]), .A2(n7140), .ZN(n6605) );
NAND2_X2 U6061 ( .A1(n5933), .A2(n6607), .ZN(cv_d[89]) );
NAND2_X2 U6062 ( .A1(cv_q[89]), .A2(n7153), .ZN(n6607) );
NAND2_X2 U6064 ( .A1(cv[89]), .A2(n7125), .ZN(n6609) );
NAND2_X2 U6065 ( .A1(cv_next[89]), .A2(n7140), .ZN(n6608) );
NAND2_X2 U6066 ( .A1(n5935), .A2(n6610), .ZN(cv_d[88]) );
NAND2_X2 U6067 ( .A1(cv_q[88]), .A2(n7153), .ZN(n6610) );
NAND2_X2 U6069 ( .A1(cv[88]), .A2(n7125), .ZN(n6612) );
NAND2_X2 U6070 ( .A1(cv_next[88]), .A2(n7140), .ZN(n6611) );
NAND2_X2 U6071 ( .A1(n5937), .A2(n6613), .ZN(cv_d[87]) );
NAND2_X2 U6072 ( .A1(cv_q[87]), .A2(n7153), .ZN(n6613) );
NAND2_X2 U6074 ( .A1(cv[87]), .A2(n7125), .ZN(n6615) );
NAND2_X2 U6075 ( .A1(cv_next[87]), .A2(n7140), .ZN(n6614) );
NAND2_X2 U6076 ( .A1(n5939), .A2(n6616), .ZN(cv_d[86]) );
NAND2_X2 U6077 ( .A1(cv_q[86]), .A2(n7153), .ZN(n6616) );
NAND2_X2 U6079 ( .A1(cv[86]), .A2(n7125), .ZN(n6618) );
NAND2_X2 U6080 ( .A1(cv_next[86]), .A2(n7140), .ZN(n6617) );
NAND2_X2 U6081 ( .A1(n5941), .A2(n6619), .ZN(cv_d[85]) );
NAND2_X2 U6082 ( .A1(cv_q[85]), .A2(n7153), .ZN(n6619) );
NAND2_X2 U6084 ( .A1(cv[85]), .A2(n7125), .ZN(n6621) );
NAND2_X2 U6085 ( .A1(cv_next[85]), .A2(n7140), .ZN(n6620) );
NAND2_X2 U6086 ( .A1(n5943), .A2(n6622), .ZN(cv_d[84]) );
NAND2_X2 U6087 ( .A1(cv_q[84]), .A2(n7153), .ZN(n6622) );
NAND2_X2 U6089 ( .A1(cv[84]), .A2(n7125), .ZN(n6624) );
NAND2_X2 U6090 ( .A1(cv_next[84]), .A2(n7140), .ZN(n6623) );
NAND2_X2 U6091 ( .A1(n5945), .A2(n6625), .ZN(cv_d[83]) );
NAND2_X2 U6092 ( .A1(cv_q[83]), .A2(n7153), .ZN(n6625) );
NAND2_X2 U6094 ( .A1(cv[83]), .A2(n7125), .ZN(n6627) );
NAND2_X2 U6095 ( .A1(cv_next[83]), .A2(n7140), .ZN(n6626) );
NAND2_X2 U6096 ( .A1(n5947), .A2(n6628), .ZN(cv_d[82]) );
NAND2_X2 U6097 ( .A1(cv_q[82]), .A2(n7153), .ZN(n6628) );
NAND2_X2 U6099 ( .A1(cv[82]), .A2(n7125), .ZN(n6630) );
NAND2_X2 U6100 ( .A1(cv_next[82]), .A2(n7140), .ZN(n6629) );
NAND2_X2 U6101 ( .A1(n5949), .A2(n6631), .ZN(cv_d[81]) );
NAND2_X2 U6102 ( .A1(cv_q[81]), .A2(n7153), .ZN(n6631) );
NAND2_X2 U6104 ( .A1(cv[81]), .A2(n7125), .ZN(n6633) );
NAND2_X2 U6105 ( .A1(cv_next[81]), .A2(n7140), .ZN(n6632) );
NAND2_X2 U6106 ( .A1(n5951), .A2(n6634), .ZN(cv_d[80]) );
NAND2_X2 U6107 ( .A1(cv_q[80]), .A2(n7153), .ZN(n6634) );
NAND2_X2 U6109 ( .A1(cv[80]), .A2(n7125), .ZN(n6636) );
NAND2_X2 U6110 ( .A1(cv_next[80]), .A2(n7140), .ZN(n6635) );
NAND2_X2 U6111 ( .A1(n5953), .A2(n6637), .ZN(cv_d[7]) );
NAND2_X2 U6112 ( .A1(cv_q[7]), .A2(n7153), .ZN(n6637) );
NAND2_X2 U6114 ( .A1(cv[7]), .A2(n7126), .ZN(n6639) );
NAND2_X2 U6115 ( .A1(cv_next[7]), .A2(n7141), .ZN(n6638) );
NAND2_X2 U6116 ( .A1(n5955), .A2(n6640), .ZN(cv_d[79]) );
NAND2_X2 U6117 ( .A1(cv_q[79]), .A2(n7153), .ZN(n6640) );
NAND2_X2 U6119 ( .A1(cv[79]), .A2(n7126), .ZN(n6642) );
NAND2_X2 U6120 ( .A1(cv_next[79]), .A2(n7141), .ZN(n6641) );
NAND2_X2 U6121 ( .A1(n5957), .A2(n6643), .ZN(cv_d[78]) );
NAND2_X2 U6122 ( .A1(cv_q[78]), .A2(n7153), .ZN(n6643) );
NAND2_X2 U6124 ( .A1(cv[78]), .A2(n7126), .ZN(n6645) );
NAND2_X2 U6125 ( .A1(cv_next[78]), .A2(n7141), .ZN(n6644) );
NAND2_X2 U6126 ( .A1(n5959), .A2(n6646), .ZN(cv_d[77]) );
NAND2_X2 U6127 ( .A1(cv_q[77]), .A2(n7153), .ZN(n6646) );
NAND2_X2 U6129 ( .A1(cv[77]), .A2(n7126), .ZN(n6648) );
NAND2_X2 U6130 ( .A1(cv_next[77]), .A2(n7141), .ZN(n6647) );
NAND2_X2 U6131 ( .A1(n5961), .A2(n6649), .ZN(cv_d[76]) );
NAND2_X2 U6132 ( .A1(cv_q[76]), .A2(n7153), .ZN(n6649) );
NAND2_X2 U6134 ( .A1(cv[76]), .A2(n7126), .ZN(n6651) );
NAND2_X2 U6135 ( .A1(cv_next[76]), .A2(n7141), .ZN(n6650) );
NAND2_X2 U6136 ( .A1(n5963), .A2(n6652), .ZN(cv_d[75]) );
NAND2_X2 U6137 ( .A1(cv_q[75]), .A2(n7153), .ZN(n6652) );
NAND2_X2 U6139 ( .A1(cv[75]), .A2(n7126), .ZN(n6654) );
NAND2_X2 U6140 ( .A1(cv_next[75]), .A2(n7141), .ZN(n6653) );
NAND2_X2 U6141 ( .A1(n5965), .A2(n6655), .ZN(cv_d[74]) );
NAND2_X2 U6142 ( .A1(cv_q[74]), .A2(n7153), .ZN(n6655) );
NAND2_X2 U6144 ( .A1(cv[74]), .A2(n7126), .ZN(n6657) );
NAND2_X2 U6145 ( .A1(cv_next[74]), .A2(n7141), .ZN(n6656) );
NAND2_X2 U6146 ( .A1(n5967), .A2(n6658), .ZN(cv_d[73]) );
NAND2_X2 U6147 ( .A1(cv_q[73]), .A2(n7153), .ZN(n6658) );
NAND2_X2 U6149 ( .A1(cv[73]), .A2(n7126), .ZN(n6660) );
NAND2_X2 U6150 ( .A1(cv_next[73]), .A2(n7141), .ZN(n6659) );
NAND2_X2 U6151 ( .A1(n5969), .A2(n6661), .ZN(cv_d[72]) );
NAND2_X2 U6152 ( .A1(cv_q[72]), .A2(n7154), .ZN(n6661) );
NAND2_X2 U6154 ( .A1(cv[72]), .A2(n7126), .ZN(n6663) );
NAND2_X2 U6155 ( .A1(cv_next[72]), .A2(n7141), .ZN(n6662) );
NAND2_X2 U6156 ( .A1(n5971), .A2(n6664), .ZN(cv_d[71]) );
NAND2_X2 U6157 ( .A1(cv_q[71]), .A2(n7153), .ZN(n6664) );
NAND2_X2 U6159 ( .A1(cv[71]), .A2(n7126), .ZN(n6666) );
NAND2_X2 U6160 ( .A1(cv_next[71]), .A2(n7141), .ZN(n6665) );
NAND2_X2 U6161 ( .A1(n5973), .A2(n6667), .ZN(cv_d[70]) );
NAND2_X2 U6162 ( .A1(cv_q[70]), .A2(n7153), .ZN(n6667) );
NAND2_X2 U6164 ( .A1(cv[70]), .A2(n7126), .ZN(n6669) );
NAND2_X2 U6165 ( .A1(cv_next[70]), .A2(n7141), .ZN(n6668) );
NAND2_X2 U6166 ( .A1(n5975), .A2(n6670), .ZN(cv_d[6]) );
NAND2_X2 U6167 ( .A1(cv_q[6]), .A2(n7154), .ZN(n6670) );
NAND2_X2 U6169 ( .A1(cv[6]), .A2(n7127), .ZN(n6672) );
NAND2_X2 U6170 ( .A1(cv_next[6]), .A2(n7142), .ZN(n6671) );
NAND2_X2 U6171 ( .A1(n5977), .A2(n6673), .ZN(cv_d[69]) );
NAND2_X2 U6172 ( .A1(cv_q[69]), .A2(n7154), .ZN(n6673) );
NAND2_X2 U6174 ( .A1(cv[69]), .A2(n7127), .ZN(n6675) );
NAND2_X2 U6175 ( .A1(cv_next[69]), .A2(n7142), .ZN(n6674) );
NAND2_X2 U6176 ( .A1(n5979), .A2(n6676), .ZN(cv_d[68]) );
NAND2_X2 U6177 ( .A1(cv_q[68]), .A2(n7154), .ZN(n6676) );
NAND2_X2 U6179 ( .A1(cv[68]), .A2(n7127), .ZN(n6678) );
NAND2_X2 U6180 ( .A1(cv_next[68]), .A2(n7142), .ZN(n6677) );
NAND2_X2 U6181 ( .A1(n5981), .A2(n6679), .ZN(cv_d[67]) );
NAND2_X2 U6182 ( .A1(cv_q[67]), .A2(n7154), .ZN(n6679) );
NAND2_X2 U6184 ( .A1(cv[67]), .A2(n7127), .ZN(n6681) );
NAND2_X2 U6185 ( .A1(cv_next[67]), .A2(n7142), .ZN(n6680) );
NAND2_X2 U6186 ( .A1(n5983), .A2(n6682), .ZN(cv_d[66]) );
NAND2_X2 U6187 ( .A1(cv_q[66]), .A2(n7154), .ZN(n6682) );
NAND2_X2 U6189 ( .A1(cv[66]), .A2(n7127), .ZN(n6684) );
NAND2_X2 U6190 ( .A1(cv_next[66]), .A2(n7142), .ZN(n6683) );
NAND2_X2 U6191 ( .A1(n5985), .A2(n6685), .ZN(cv_d[65]) );
NAND2_X2 U6192 ( .A1(cv_q[65]), .A2(n7154), .ZN(n6685) );
NAND2_X2 U6194 ( .A1(cv[65]), .A2(n7127), .ZN(n6687) );
NAND2_X2 U6195 ( .A1(cv_next[65]), .A2(n7142), .ZN(n6686) );
NAND2_X2 U6196 ( .A1(n5987), .A2(n6688), .ZN(cv_d[64]) );
NAND2_X2 U6197 ( .A1(cv_q[64]), .A2(n7154), .ZN(n6688) );
NAND2_X2 U6199 ( .A1(cv[64]), .A2(n7127), .ZN(n6690) );
NAND2_X2 U6200 ( .A1(cv_next[64]), .A2(n7142), .ZN(n6689) );
NAND2_X2 U6201 ( .A1(n5989), .A2(n6691), .ZN(cv_d[63]) );
NAND2_X2 U6202 ( .A1(cv_q[63]), .A2(n7154), .ZN(n6691) );
NAND2_X2 U6204 ( .A1(cv[63]), .A2(n7127), .ZN(n6693) );
NAND2_X2 U6205 ( .A1(cv_next[63]), .A2(n7142), .ZN(n6692) );
NAND2_X2 U6206 ( .A1(n5991), .A2(n6694), .ZN(cv_d[62]) );
NAND2_X2 U6207 ( .A1(cv_q[62]), .A2(n7154), .ZN(n6694) );
NAND2_X2 U6209 ( .A1(cv[62]), .A2(n7127), .ZN(n6696) );
NAND2_X2 U6210 ( .A1(cv_next[62]), .A2(n7142), .ZN(n6695) );
NAND2_X2 U6211 ( .A1(n5993), .A2(n6697), .ZN(cv_d[61]) );
NAND2_X2 U6212 ( .A1(cv_q[61]), .A2(n7154), .ZN(n6697) );
NAND2_X2 U6214 ( .A1(cv[61]), .A2(n7127), .ZN(n6699) );
NAND2_X2 U6215 ( .A1(cv_next[61]), .A2(n7142), .ZN(n6698) );
NAND2_X2 U6216 ( .A1(n5995), .A2(n6700), .ZN(cv_d[60]) );
NAND2_X2 U6217 ( .A1(cv_q[60]), .A2(n7154), .ZN(n6700) );
NAND2_X2 U6219 ( .A1(cv[60]), .A2(n7127), .ZN(n6702) );
NAND2_X2 U6220 ( .A1(cv_next[60]), .A2(n7142), .ZN(n6701) );
NAND2_X2 U6221 ( .A1(n5997), .A2(n6703), .ZN(cv_d[5]) );
NAND2_X2 U6222 ( .A1(cv_q[5]), .A2(n7154), .ZN(n6703) );
NAND2_X2 U6224 ( .A1(cv[5]), .A2(n7128), .ZN(n6705) );
NAND2_X2 U6225 ( .A1(cv_next[5]), .A2(n7143), .ZN(n6704) );
NAND2_X2 U6226 ( .A1(n5999), .A2(n6706), .ZN(cv_d[59]) );
NAND2_X2 U6227 ( .A1(cv_q[59]), .A2(n7154), .ZN(n6706) );
NAND2_X2 U6229 ( .A1(cv[59]), .A2(n7128), .ZN(n6708) );
NAND2_X2 U6230 ( .A1(cv_next[59]), .A2(n7143), .ZN(n6707) );
NAND2_X2 U6231 ( .A1(n6001), .A2(n6709), .ZN(cv_d[58]) );
NAND2_X2 U6232 ( .A1(cv_q[58]), .A2(n7154), .ZN(n6709) );
NAND2_X2 U6234 ( .A1(cv[58]), .A2(n7128), .ZN(n6711) );
NAND2_X2 U6235 ( .A1(cv_next[58]), .A2(n7143), .ZN(n6710) );
NAND2_X2 U6236 ( .A1(n6003), .A2(n6712), .ZN(cv_d[57]) );
NAND2_X2 U6237 ( .A1(cv_q[57]), .A2(n7154), .ZN(n6712) );
NAND2_X2 U6239 ( .A1(cv[57]), .A2(n7128), .ZN(n6714) );
NAND2_X2 U6240 ( .A1(cv_next[57]), .A2(n7143), .ZN(n6713) );
NAND2_X2 U6241 ( .A1(n6005), .A2(n6715), .ZN(cv_d[56]) );
NAND2_X2 U6242 ( .A1(cv_q[56]), .A2(n7154), .ZN(n6715) );
NAND2_X2 U6244 ( .A1(cv[56]), .A2(n7128), .ZN(n6717) );
NAND2_X2 U6245 ( .A1(cv_next[56]), .A2(n7143), .ZN(n6716) );
NAND2_X2 U6246 ( .A1(n6007), .A2(n6718), .ZN(cv_d[55]) );
NAND2_X2 U6247 ( .A1(cv_q[55]), .A2(n7154), .ZN(n6718) );
NAND2_X2 U6249 ( .A1(cv[55]), .A2(n7128), .ZN(n6720) );
NAND2_X2 U6250 ( .A1(cv_next[55]), .A2(n7143), .ZN(n6719) );
NAND2_X2 U6251 ( .A1(n6009), .A2(n6721), .ZN(cv_d[54]) );
NAND2_X2 U6252 ( .A1(cv_q[54]), .A2(n7154), .ZN(n6721) );
NAND2_X2 U6254 ( .A1(cv[54]), .A2(n7128), .ZN(n6723) );
NAND2_X2 U6255 ( .A1(cv_next[54]), .A2(n7143), .ZN(n6722) );
NAND2_X2 U6256 ( .A1(n6011), .A2(n6724), .ZN(cv_d[53]) );
NAND2_X2 U6257 ( .A1(cv_q[53]), .A2(n7154), .ZN(n6724) );
NAND2_X2 U6259 ( .A1(cv[53]), .A2(n7128), .ZN(n6726) );
NAND2_X2 U6260 ( .A1(cv_next[53]), .A2(n7143), .ZN(n6725) );
NAND2_X2 U6261 ( .A1(n6013), .A2(n6727), .ZN(cv_d[52]) );
NAND2_X2 U6262 ( .A1(cv_q[52]), .A2(n7154), .ZN(n6727) );
NAND2_X2 U6264 ( .A1(cv[52]), .A2(n7128), .ZN(n6729) );
NAND2_X2 U6265 ( .A1(cv_next[52]), .A2(n7143), .ZN(n6728) );
NAND2_X2 U6266 ( .A1(n6015), .A2(n6730), .ZN(cv_d[51]) );
NAND2_X2 U6267 ( .A1(cv_q[51]), .A2(n7154), .ZN(n6730) );
NAND2_X2 U6269 ( .A1(cv[51]), .A2(n7128), .ZN(n6732) );
NAND2_X2 U6270 ( .A1(cv_next[51]), .A2(n7143), .ZN(n6731) );
NAND2_X2 U6271 ( .A1(n6017), .A2(n6733), .ZN(cv_d[50]) );
NAND2_X2 U6272 ( .A1(cv_q[50]), .A2(n7154), .ZN(n6733) );
NAND2_X2 U6274 ( .A1(cv[50]), .A2(n7128), .ZN(n6735) );
NAND2_X2 U6275 ( .A1(cv_next[50]), .A2(n7143), .ZN(n6734) );
NAND2_X2 U6276 ( .A1(n6019), .A2(n6736), .ZN(cv_d[4]) );
NAND2_X2 U6277 ( .A1(cv_q[4]), .A2(n7154), .ZN(n6736) );
NAND2_X2 U6279 ( .A1(cv[4]), .A2(n7129), .ZN(n6738) );
NAND2_X2 U6280 ( .A1(cv_next[4]), .A2(n7144), .ZN(n6737) );
NAND2_X2 U6281 ( .A1(n6021), .A2(n6739), .ZN(cv_d[49]) );
NAND2_X2 U6282 ( .A1(cv_q[49]), .A2(n7154), .ZN(n6739) );
NAND2_X2 U6284 ( .A1(cv[49]), .A2(n7129), .ZN(n6741) );
NAND2_X2 U6285 ( .A1(cv_next[49]), .A2(n7144), .ZN(n6740) );
NAND2_X2 U6286 ( .A1(n6023), .A2(n6742), .ZN(cv_d[48]) );
NAND2_X2 U6287 ( .A1(cv_q[48]), .A2(n7154), .ZN(n6742) );
NAND2_X2 U6289 ( .A1(cv[48]), .A2(n7129), .ZN(n6744) );
NAND2_X2 U6290 ( .A1(cv_next[48]), .A2(n7144), .ZN(n6743) );
NAND2_X2 U6291 ( .A1(n6025), .A2(n6745), .ZN(cv_d[47]) );
NAND2_X2 U6292 ( .A1(cv_q[47]), .A2(n7154), .ZN(n6745) );
NAND2_X2 U6294 ( .A1(cv[47]), .A2(n7129), .ZN(n6747) );
NAND2_X2 U6295 ( .A1(cv_next[47]), .A2(n7144), .ZN(n6746) );
NAND2_X2 U6296 ( .A1(n6027), .A2(n6748), .ZN(cv_d[46]) );
NAND2_X2 U6297 ( .A1(cv_q[46]), .A2(n7155), .ZN(n6748) );
NAND2_X2 U6299 ( .A1(cv[46]), .A2(n7129), .ZN(n6750) );
NAND2_X2 U6300 ( .A1(cv_next[46]), .A2(n7144), .ZN(n6749) );
NAND2_X2 U6301 ( .A1(n6029), .A2(n6751), .ZN(cv_d[45]) );
NAND2_X2 U6302 ( .A1(cv_q[45]), .A2(n7155), .ZN(n6751) );
NAND2_X2 U6304 ( .A1(cv[45]), .A2(n7129), .ZN(n6753) );
NAND2_X2 U6305 ( .A1(cv_next[45]), .A2(n7144), .ZN(n6752) );
NAND2_X2 U6306 ( .A1(n6031), .A2(n6754), .ZN(cv_d[44]) );
NAND2_X2 U6307 ( .A1(cv_q[44]), .A2(n7155), .ZN(n6754) );
NAND2_X2 U6309 ( .A1(cv[44]), .A2(n7129), .ZN(n6756) );
NAND2_X2 U6310 ( .A1(cv_next[44]), .A2(n7144), .ZN(n6755) );
NAND2_X2 U6311 ( .A1(n6033), .A2(n6757), .ZN(cv_d[43]) );
NAND2_X2 U6312 ( .A1(cv_q[43]), .A2(n7155), .ZN(n6757) );
NAND2_X2 U6314 ( .A1(cv[43]), .A2(n7129), .ZN(n6759) );
NAND2_X2 U6315 ( .A1(cv_next[43]), .A2(n7144), .ZN(n6758) );
NAND2_X2 U6316 ( .A1(n6035), .A2(n6760), .ZN(cv_d[42]) );
NAND2_X2 U6317 ( .A1(cv_q[42]), .A2(n7155), .ZN(n6760) );
NAND2_X2 U6319 ( .A1(cv[42]), .A2(n7129), .ZN(n6762) );
NAND2_X2 U6320 ( .A1(cv_next[42]), .A2(n7144), .ZN(n6761) );
NAND2_X2 U6321 ( .A1(n6037), .A2(n6763), .ZN(cv_d[41]) );
NAND2_X2 U6322 ( .A1(cv_q[41]), .A2(n7155), .ZN(n6763) );
NAND2_X2 U6324 ( .A1(cv[41]), .A2(n7129), .ZN(n6765) );
NAND2_X2 U6325 ( .A1(cv_next[41]), .A2(n7144), .ZN(n6764) );
NAND2_X2 U6326 ( .A1(n6039), .A2(n6766), .ZN(cv_d[40]) );
NAND2_X2 U6327 ( .A1(cv_q[40]), .A2(n7155), .ZN(n6766) );
NAND2_X2 U6329 ( .A1(cv[40]), .A2(n7129), .ZN(n6768) );
NAND2_X2 U6330 ( .A1(cv_next[40]), .A2(n7144), .ZN(n6767) );
NAND2_X2 U6331 ( .A1(n6041), .A2(n6769), .ZN(cv_d[3]) );
NAND2_X2 U6332 ( .A1(cv_q[3]), .A2(n7155), .ZN(n6769) );
NAND2_X2 U6334 ( .A1(cv[3]), .A2(n7130), .ZN(n6771) );
NAND2_X2 U6335 ( .A1(cv_next[3]), .A2(n7145), .ZN(n6770) );
NAND2_X2 U6336 ( .A1(n6043), .A2(n6772), .ZN(cv_d[39]) );
NAND2_X2 U6337 ( .A1(cv_q[39]), .A2(n7155), .ZN(n6772) );
NAND2_X2 U6339 ( .A1(cv[39]), .A2(n7130), .ZN(n6774) );
NAND2_X2 U6340 ( .A1(cv_next[39]), .A2(n7145), .ZN(n6773) );
NAND2_X2 U6341 ( .A1(n6045), .A2(n6775), .ZN(cv_d[38]) );
NAND2_X2 U6342 ( .A1(cv_q[38]), .A2(n7155), .ZN(n6775) );
NAND2_X2 U6344 ( .A1(cv[38]), .A2(n7130), .ZN(n6777) );
NAND2_X2 U6345 ( .A1(cv_next[38]), .A2(n7145), .ZN(n6776) );
NAND2_X2 U6346 ( .A1(n6047), .A2(n6778), .ZN(cv_d[37]) );
NAND2_X2 U6347 ( .A1(cv_q[37]), .A2(n7155), .ZN(n6778) );
NAND2_X2 U6349 ( .A1(cv[37]), .A2(n7130), .ZN(n6780) );
NAND2_X2 U6350 ( .A1(cv_next[37]), .A2(n7145), .ZN(n6779) );
NAND2_X2 U6351 ( .A1(n6049), .A2(n6781), .ZN(cv_d[36]) );
NAND2_X2 U6352 ( .A1(cv_q[36]), .A2(n7155), .ZN(n6781) );
NAND2_X2 U6354 ( .A1(cv[36]), .A2(n7130), .ZN(n6783) );
NAND2_X2 U6355 ( .A1(cv_next[36]), .A2(n7145), .ZN(n6782) );
NAND2_X2 U6356 ( .A1(n6051), .A2(n6784), .ZN(cv_d[35]) );
NAND2_X2 U6357 ( .A1(cv_q[35]), .A2(n7155), .ZN(n6784) );
NAND2_X2 U6359 ( .A1(cv[35]), .A2(n7130), .ZN(n6786) );
NAND2_X2 U6360 ( .A1(cv_next[35]), .A2(n7145), .ZN(n6785) );
NAND2_X2 U6361 ( .A1(n6053), .A2(n6787), .ZN(cv_d[34]) );
NAND2_X2 U6362 ( .A1(cv_q[34]), .A2(n7155), .ZN(n6787) );
NAND2_X2 U6364 ( .A1(cv[34]), .A2(n7130), .ZN(n6789) );
NAND2_X2 U6365 ( .A1(cv_next[34]), .A2(n7145), .ZN(n6788) );
NAND2_X2 U6366 ( .A1(n6055), .A2(n6790), .ZN(cv_d[33]) );
NAND2_X2 U6367 ( .A1(cv_q[33]), .A2(n7155), .ZN(n6790) );
NAND2_X2 U6369 ( .A1(cv[33]), .A2(n7130), .ZN(n6792) );
NAND2_X2 U6370 ( .A1(cv_next[33]), .A2(n7145), .ZN(n6791) );
NAND2_X2 U6371 ( .A1(n6057), .A2(n6793), .ZN(cv_d[32]) );
NAND2_X2 U6372 ( .A1(cv_q[32]), .A2(n7155), .ZN(n6793) );
NAND2_X2 U6374 ( .A1(cv[32]), .A2(n7130), .ZN(n6795) );
NAND2_X2 U6375 ( .A1(cv_next[32]), .A2(n7145), .ZN(n6794) );
NAND2_X2 U6376 ( .A1(n6059), .A2(n6796), .ZN(cv_d[31]) );
NAND2_X2 U6377 ( .A1(cv_q[31]), .A2(n7155), .ZN(n6796) );
NAND2_X2 U6379 ( .A1(cv[31]), .A2(n7130), .ZN(n6798) );
NAND2_X2 U6380 ( .A1(cv_next[31]), .A2(n7145), .ZN(n6797) );
NAND2_X2 U6381 ( .A1(n6061), .A2(n6799), .ZN(cv_d[30]) );
NAND2_X2 U6382 ( .A1(cv_q[30]), .A2(n7155), .ZN(n6799) );
NAND2_X2 U6384 ( .A1(cv[30]), .A2(n7130), .ZN(n6801) );
NAND2_X2 U6385 ( .A1(cv_next[30]), .A2(n7145), .ZN(n6800) );
NAND2_X2 U6386 ( .A1(n6063), .A2(n6802), .ZN(cv_d[2]) );
NAND2_X2 U6387 ( .A1(cv_q[2]), .A2(n7155), .ZN(n6802) );
NAND2_X2 U6389 ( .A1(cv[2]), .A2(n7131), .ZN(n6804) );
NAND2_X2 U6390 ( .A1(cv_next[2]), .A2(n7146), .ZN(n6803) );
NAND2_X2 U6391 ( .A1(n6065), .A2(n6805), .ZN(cv_d[29]) );
NAND2_X2 U6392 ( .A1(cv_q[29]), .A2(n7155), .ZN(n6805) );
NAND2_X2 U6394 ( .A1(cv[29]), .A2(n7131), .ZN(n6807) );
NAND2_X2 U6395 ( .A1(cv_next[29]), .A2(n7146), .ZN(n6806) );
NAND2_X2 U6396 ( .A1(n6067), .A2(n6808), .ZN(cv_d[28]) );
NAND2_X2 U6397 ( .A1(cv_q[28]), .A2(n7155), .ZN(n6808) );
NAND2_X2 U6399 ( .A1(cv[28]), .A2(n7131), .ZN(n6810) );
NAND2_X2 U6400 ( .A1(cv_next[28]), .A2(n7146), .ZN(n6809) );
NAND2_X2 U6401 ( .A1(n6069), .A2(n6811), .ZN(cv_d[27]) );
NAND2_X2 U6402 ( .A1(cv_q[27]), .A2(n7155), .ZN(n6811) );
NAND2_X2 U6404 ( .A1(cv[27]), .A2(n7131), .ZN(n6813) );
NAND2_X2 U6405 ( .A1(cv_next[27]), .A2(n7146), .ZN(n6812) );
NAND2_X2 U6406 ( .A1(n6071), .A2(n6814), .ZN(cv_d[26]) );
NAND2_X2 U6407 ( .A1(cv_q[26]), .A2(n7155), .ZN(n6814) );
NAND2_X2 U6409 ( .A1(cv[26]), .A2(n7131), .ZN(n6816) );
NAND2_X2 U6410 ( .A1(cv_next[26]), .A2(n7146), .ZN(n6815) );
NAND2_X2 U6411 ( .A1(n6073), .A2(n6817), .ZN(cv_d[25]) );
NAND2_X2 U6412 ( .A1(cv_q[25]), .A2(n7155), .ZN(n6817) );
NAND2_X2 U6414 ( .A1(cv[25]), .A2(n7131), .ZN(n6819) );
NAND2_X2 U6415 ( .A1(cv_next[25]), .A2(n7146), .ZN(n6818) );
NAND2_X2 U6416 ( .A1(n6075), .A2(n6820), .ZN(cv_d[24]) );
NAND2_X2 U6417 ( .A1(cv_q[24]), .A2(n7155), .ZN(n6820) );
NAND2_X2 U6419 ( .A1(cv[24]), .A2(n7131), .ZN(n6822) );
NAND2_X2 U6420 ( .A1(cv_next[24]), .A2(n7146), .ZN(n6821) );
NAND2_X2 U6421 ( .A1(n6077), .A2(n6823), .ZN(cv_d[23]) );
NAND2_X2 U6422 ( .A1(cv_q[23]), .A2(n7155), .ZN(n6823) );
NAND2_X2 U6424 ( .A1(cv[23]), .A2(n7131), .ZN(n6825) );
NAND2_X2 U6425 ( .A1(cv_next[23]), .A2(n7146), .ZN(n6824) );
NAND2_X2 U6426 ( .A1(n6079), .A2(n6826), .ZN(cv_d[22]) );
NAND2_X2 U6427 ( .A1(cv_q[22]), .A2(n7156), .ZN(n6826) );
NAND2_X2 U6429 ( .A1(cv[22]), .A2(n7131), .ZN(n6828) );
NAND2_X2 U6430 ( .A1(cv_next[22]), .A2(n7146), .ZN(n6827) );
NAND2_X2 U6431 ( .A1(n6081), .A2(n6829), .ZN(cv_d[21]) );
NAND2_X2 U6432 ( .A1(cv_q[21]), .A2(n7156), .ZN(n6829) );
NAND2_X2 U6434 ( .A1(cv[21]), .A2(n7131), .ZN(n6831) );
NAND2_X2 U6435 ( .A1(cv_next[21]), .A2(n7146), .ZN(n6830) );
NAND2_X2 U6436 ( .A1(n6083), .A2(n6832), .ZN(cv_d[20]) );
NAND2_X2 U6437 ( .A1(cv_q[20]), .A2(n7156), .ZN(n6832) );
NAND2_X2 U6439 ( .A1(cv[20]), .A2(n7131), .ZN(n6834) );
NAND2_X2 U6440 ( .A1(cv_next[20]), .A2(n7146), .ZN(n6833) );
NAND2_X2 U6441 ( .A1(n6085), .A2(n6835), .ZN(cv_d[1]) );
NAND2_X2 U6442 ( .A1(cv_q[1]), .A2(n7156), .ZN(n6835) );
NAND2_X2 U6444 ( .A1(cv[1]), .A2(n7132), .ZN(n6837) );
NAND2_X2 U6445 ( .A1(cv_next[1]), .A2(n7147), .ZN(n6836) );
NAND2_X2 U6446 ( .A1(n6087), .A2(n6838), .ZN(cv_d[19]) );
NAND2_X2 U6447 ( .A1(cv_q[19]), .A2(n7156), .ZN(n6838) );
NAND2_X2 U6449 ( .A1(cv[19]), .A2(n7132), .ZN(n6840) );
NAND2_X2 U6450 ( .A1(cv_next[19]), .A2(n7147), .ZN(n6839) );
NAND2_X2 U6451 ( .A1(n6089), .A2(n6841), .ZN(cv_d[18]) );
NAND2_X2 U6452 ( .A1(cv_q[18]), .A2(n7156), .ZN(n6841) );
NAND2_X2 U6454 ( .A1(cv[18]), .A2(n7132), .ZN(n6843) );
NAND2_X2 U6455 ( .A1(cv_next[18]), .A2(n7147), .ZN(n6842) );
NAND2_X2 U6456 ( .A1(n6091), .A2(n6844), .ZN(cv_d[17]) );
NAND2_X2 U6457 ( .A1(cv_q[17]), .A2(n7156), .ZN(n6844) );
NAND2_X2 U6459 ( .A1(cv[17]), .A2(n7132), .ZN(n6846) );
NAND2_X2 U6460 ( .A1(cv_next[17]), .A2(n7147), .ZN(n6845) );
NAND2_X2 U6461 ( .A1(n6093), .A2(n6847), .ZN(cv_d[16]) );
NAND2_X2 U6462 ( .A1(cv_q[16]), .A2(n7156), .ZN(n6847) );
NAND2_X2 U6464 ( .A1(cv[16]), .A2(n7132), .ZN(n6849) );
NAND2_X2 U6465 ( .A1(cv_next[16]), .A2(n7147), .ZN(n6848) );
NAND2_X2 U6466 ( .A1(n6095), .A2(n6850), .ZN(cv_d[15]) );
NAND2_X2 U6467 ( .A1(cv_q[15]), .A2(n7156), .ZN(n6850) );
NAND2_X2 U6469 ( .A1(cv[15]), .A2(n7132), .ZN(n6852) );
NAND2_X2 U6470 ( .A1(cv_next[15]), .A2(n7147), .ZN(n6851) );
NAND2_X2 U6471 ( .A1(n7373), .A2(n6853), .ZN(cv_d[159]) );
NAND2_X2 U6472 ( .A1(cv_q[159]), .A2(n7156), .ZN(n6853) );
NAND2_X2 U6477 ( .A1(cv_q[158]), .A2(n7156), .ZN(n6856) );
NAND2_X2 U6481 ( .A1(n7375), .A2(n6859), .ZN(cv_d[157]) );
NAND2_X2 U6482 ( .A1(cv_q[157]), .A2(n7156), .ZN(n6859) );
NAND2_X2 U6486 ( .A1(n7376), .A2(n6862), .ZN(cv_d[156]) );
NAND2_X2 U6487 ( .A1(cv_q[156]), .A2(n7156), .ZN(n6862) );
NAND2_X2 U6492 ( .A1(cv_q[155]), .A2(n7156), .ZN(n6865) );
NAND2_X2 U6497 ( .A1(cv_q[154]), .A2(n7156), .ZN(n6868) );
NAND2_X2 U6502 ( .A1(cv_q[153]), .A2(n7156), .ZN(n6871) );
NAND2_X2 U6506 ( .A1(n7380), .A2(n6874), .ZN(cv_d[152]) );
NAND2_X2 U6507 ( .A1(cv_q[152]), .A2(n7156), .ZN(n6874) );
NAND2_X2 U6511 ( .A1(n7381), .A2(n6877), .ZN(cv_d[151]) );
NAND2_X2 U6512 ( .A1(cv_q[151]), .A2(n7156), .ZN(n6877) );
NAND2_X2 U6516 ( .A1(n7382), .A2(n6880), .ZN(cv_d[150]) );
NAND2_X2 U6517 ( .A1(cv_q[150]), .A2(n7156), .ZN(n6880) );
NAND2_X2 U6521 ( .A1(n6117), .A2(n6883), .ZN(cv_d[14]) );
NAND2_X2 U6522 ( .A1(cv_q[14]), .A2(n7156), .ZN(n6883) );
NAND2_X2 U6524 ( .A1(cv[14]), .A2(n7132), .ZN(n6885) );
NAND2_X2 U6525 ( .A1(cv_next[14]), .A2(n7147), .ZN(n6884) );
NAND2_X2 U6527 ( .A1(cv_q[149]), .A2(n7156), .ZN(n6886) );
NAND2_X2 U6531 ( .A1(n7384), .A2(n6889), .ZN(cv_d[148]) );
NAND2_X2 U6532 ( .A1(cv_q[148]), .A2(n7156), .ZN(n6889) );
NAND2_X2 U6536 ( .A1(n7385), .A2(n6892), .ZN(cv_d[147]) );
NAND2_X2 U6537 ( .A1(cv_q[147]), .A2(n7156), .ZN(n6892) );
NAND2_X2 U6541 ( .A1(n7386), .A2(n6895), .ZN(cv_d[146]) );
NAND2_X2 U6542 ( .A1(cv_q[146]), .A2(n7156), .ZN(n6895) );
NAND2_X2 U6546 ( .A1(n7387), .A2(n6898), .ZN(cv_d[145]) );
NAND2_X2 U6547 ( .A1(cv_q[145]), .A2(n7156), .ZN(n6898) );
NAND2_X2 U6551 ( .A1(n7388), .A2(n6901), .ZN(cv_d[144]) );
NAND2_X2 U6552 ( .A1(cv_q[144]), .A2(n7156), .ZN(n6901) );
NAND2_X2 U6556 ( .A1(n7389), .A2(n6904), .ZN(cv_d[143]) );
NAND2_X2 U6557 ( .A1(cv_q[143]), .A2(n7156), .ZN(n6904) );
NAND2_X2 U6561 ( .A1(n7390), .A2(n6907), .ZN(cv_d[142]) );
NAND2_X2 U6562 ( .A1(cv_q[142]), .A2(n7157), .ZN(n6907) );
NAND2_X2 U6566 ( .A1(n7391), .A2(n6910), .ZN(cv_d[141]) );
NAND2_X2 U6567 ( .A1(cv_q[141]), .A2(n7157), .ZN(n6910) );
NAND2_X2 U6571 ( .A1(n7392), .A2(n6913), .ZN(cv_d[140]) );
NAND2_X2 U6572 ( .A1(cv_q[140]), .A2(n7157), .ZN(n6913) );
NAND2_X2 U6576 ( .A1(n6139), .A2(n6916), .ZN(cv_d[13]) );
NAND2_X2 U6577 ( .A1(cv_q[13]), .A2(n7157), .ZN(n6916) );
NAND2_X2 U6579 ( .A1(cv[13]), .A2(n7132), .ZN(n6918) );
NAND2_X2 U6580 ( .A1(cv_next[13]), .A2(n7147), .ZN(n6917) );
NAND2_X2 U6581 ( .A1(n7393), .A2(n6919), .ZN(cv_d[139]) );
NAND2_X2 U6582 ( .A1(cv_q[139]), .A2(n7157), .ZN(n6919) );
NAND2_X2 U6586 ( .A1(n7394), .A2(n6922), .ZN(cv_d[138]) );
NAND2_X2 U6587 ( .A1(cv_q[138]), .A2(n7157), .ZN(n6922) );
NAND2_X2 U6591 ( .A1(n6145), .A2(n6925), .ZN(cv_d[137]) );
NAND2_X2 U6592 ( .A1(cv_q[137]), .A2(n7157), .ZN(n6925) );
NAND2_X2 U6594 ( .A1(cv[137]), .A2(n7132), .ZN(n6927) );
NAND2_X2 U6595 ( .A1(cv_next[137]), .A2(n7147), .ZN(n6926) );
NAND2_X2 U6596 ( .A1(n6147), .A2(n6928), .ZN(cv_d[136]) );
NAND2_X2 U6597 ( .A1(cv_q[136]), .A2(n7157), .ZN(n6928) );
NAND2_X2 U6599 ( .A1(cv[136]), .A2(n7132), .ZN(n6930) );
NAND2_X2 U6600 ( .A1(cv_next[136]), .A2(n7147), .ZN(n6929) );
NAND2_X2 U6601 ( .A1(n6149), .A2(n6931), .ZN(cv_d[135]) );
NAND2_X2 U6602 ( .A1(cv_q[135]), .A2(n7157), .ZN(n6931) );
NAND2_X2 U6604 ( .A1(cv[135]), .A2(n7132), .ZN(n6933) );
NAND2_X2 U6605 ( .A1(cv_next[135]), .A2(n7147), .ZN(n6932) );
NAND2_X2 U6606 ( .A1(n6151), .A2(n6934), .ZN(cv_d[134]) );
NAND2_X2 U6607 ( .A1(cv_q[134]), .A2(n7157), .ZN(n6934) );
NAND2_X2 U6609 ( .A1(cv[134]), .A2(n7133), .ZN(n6936) );
NAND2_X2 U6610 ( .A1(cv_next[134]), .A2(n7148), .ZN(n6935) );
NAND2_X2 U6611 ( .A1(n6153), .A2(n6937), .ZN(cv_d[133]) );
NAND2_X2 U6612 ( .A1(cv_q[133]), .A2(n7157), .ZN(n6937) );
NAND2_X2 U6614 ( .A1(cv[133]), .A2(n7133), .ZN(n6939) );
NAND2_X2 U6615 ( .A1(cv_next[133]), .A2(n7148), .ZN(n6938) );
NAND2_X2 U6616 ( .A1(n6155), .A2(n6940), .ZN(cv_d[132]) );
NAND2_X2 U6617 ( .A1(cv_q[132]), .A2(n7157), .ZN(n6940) );
NAND2_X2 U6619 ( .A1(cv[132]), .A2(n7133), .ZN(n6942) );
NAND2_X2 U6620 ( .A1(cv_next[132]), .A2(n7148), .ZN(n6941) );
NAND2_X2 U6621 ( .A1(n6157), .A2(n6943), .ZN(cv_d[131]) );
NAND2_X2 U6622 ( .A1(cv_q[131]), .A2(n7157), .ZN(n6943) );
NAND2_X2 U6624 ( .A1(cv[131]), .A2(n7133), .ZN(n6945) );
NAND2_X2 U6625 ( .A1(cv_next[131]), .A2(n7148), .ZN(n6944) );
NAND2_X2 U6626 ( .A1(n6159), .A2(n6946), .ZN(cv_d[130]) );
NAND2_X2 U6627 ( .A1(cv_q[130]), .A2(n7157), .ZN(n6946) );
NAND2_X2 U6629 ( .A1(cv[130]), .A2(n7133), .ZN(n6948) );
NAND2_X2 U6630 ( .A1(cv_next[130]), .A2(n7148), .ZN(n6947) );
NAND2_X2 U6631 ( .A1(n6161), .A2(n6949), .ZN(cv_d[12]) );
NAND2_X2 U6632 ( .A1(cv_q[12]), .A2(n7157), .ZN(n6949) );
NAND2_X2 U6634 ( .A1(cv[12]), .A2(n7133), .ZN(n6951) );
NAND2_X2 U6635 ( .A1(cv_next[12]), .A2(n7148), .ZN(n6950) );
NAND2_X2 U6636 ( .A1(n6163), .A2(n6952), .ZN(cv_d[129]) );
NAND2_X2 U6637 ( .A1(cv_q[129]), .A2(n7157), .ZN(n6952) );
NAND2_X2 U6639 ( .A1(cv[129]), .A2(n7133), .ZN(n6954) );
NAND2_X2 U6640 ( .A1(cv_next[129]), .A2(n7148), .ZN(n6953) );
NAND2_X2 U6641 ( .A1(n6165), .A2(n6955), .ZN(cv_d[128]) );
NAND2_X2 U6642 ( .A1(cv_q[128]), .A2(n7157), .ZN(n6955) );
NAND2_X2 U6644 ( .A1(cv[128]), .A2(n7133), .ZN(n6957) );
NAND2_X2 U6645 ( .A1(cv_next[128]), .A2(n7148), .ZN(n6956) );
NAND2_X2 U6646 ( .A1(n6167), .A2(n6958), .ZN(cv_d[127]) );
NAND2_X2 U6647 ( .A1(cv_q[127]), .A2(n7157), .ZN(n6958) );
NAND2_X2 U6649 ( .A1(cv[127]), .A2(n7133), .ZN(n6960) );
NAND2_X2 U6650 ( .A1(cv_next[127]), .A2(n7148), .ZN(n6959) );
NAND2_X2 U6651 ( .A1(n6169), .A2(n6961), .ZN(cv_d[126]) );
NAND2_X2 U6652 ( .A1(cv_q[126]), .A2(n7157), .ZN(n6961) );
NAND2_X2 U6654 ( .A1(cv[126]), .A2(n7133), .ZN(n6963) );
NAND2_X2 U6655 ( .A1(cv_next[126]), .A2(n7148), .ZN(n6962) );
NAND2_X2 U6656 ( .A1(n6171), .A2(n6964), .ZN(cv_d[125]) );
NAND2_X2 U6657 ( .A1(cv_q[125]), .A2(n7157), .ZN(n6964) );
NAND2_X2 U6659 ( .A1(cv[125]), .A2(n7133), .ZN(n6966) );
NAND2_X2 U6660 ( .A1(cv_next[125]), .A2(n7148), .ZN(n6965) );
NAND2_X2 U6661 ( .A1(n6173), .A2(n6967), .ZN(cv_d[124]) );
NAND2_X2 U6662 ( .A1(cv_q[124]), .A2(n7157), .ZN(n6967) );
NAND2_X2 U6664 ( .A1(cv[124]), .A2(n7134), .ZN(n6969) );
NAND2_X2 U6665 ( .A1(cv_next[124]), .A2(n7149), .ZN(n6968) );
NAND2_X2 U6666 ( .A1(n6175), .A2(n6970), .ZN(cv_d[123]) );
NAND2_X2 U6667 ( .A1(cv_q[123]), .A2(n7157), .ZN(n6970) );
NAND2_X2 U6669 ( .A1(cv[123]), .A2(n7134), .ZN(n6972) );
NAND2_X2 U6670 ( .A1(cv_next[123]), .A2(n7149), .ZN(n6971) );
NAND2_X2 U6671 ( .A1(n6177), .A2(n6973), .ZN(cv_d[122]) );
NAND2_X2 U6672 ( .A1(cv_q[122]), .A2(n7157), .ZN(n6973) );
NAND2_X2 U6674 ( .A1(cv[122]), .A2(n7134), .ZN(n6975) );
NAND2_X2 U6675 ( .A1(cv_next[122]), .A2(n7149), .ZN(n6974) );
NAND2_X2 U6676 ( .A1(n6179), .A2(n6976), .ZN(cv_d[121]) );
NAND2_X2 U6677 ( .A1(cv_q[121]), .A2(n7157), .ZN(n6976) );
NAND2_X2 U6679 ( .A1(cv[121]), .A2(n7134), .ZN(n6978) );
NAND2_X2 U6680 ( .A1(cv_next[121]), .A2(n7149), .ZN(n6977) );
NAND2_X2 U6681 ( .A1(n6181), .A2(n6979), .ZN(cv_d[120]) );
NAND2_X2 U6682 ( .A1(cv_q[120]), .A2(n7157), .ZN(n6979) );
NAND2_X2 U6684 ( .A1(cv[120]), .A2(n7134), .ZN(n6981) );
NAND2_X2 U6685 ( .A1(cv_next[120]), .A2(n7149), .ZN(n6980) );
NAND2_X2 U6686 ( .A1(n6183), .A2(n6982), .ZN(cv_d[11]) );
NAND2_X2 U6687 ( .A1(cv_q[11]), .A2(n7157), .ZN(n6982) );
NAND2_X2 U6689 ( .A1(cv[11]), .A2(n7134), .ZN(n6984) );
NAND2_X2 U6690 ( .A1(cv_next[11]), .A2(n7149), .ZN(n6983) );
NAND2_X2 U6691 ( .A1(n6185), .A2(n6985), .ZN(cv_d[119]) );
NAND2_X2 U6692 ( .A1(cv_q[119]), .A2(n7157), .ZN(n6985) );
NAND2_X2 U6694 ( .A1(cv[119]), .A2(n7134), .ZN(n6987) );
NAND2_X2 U6695 ( .A1(cv_next[119]), .A2(n7149), .ZN(n6986) );
NAND2_X2 U6696 ( .A1(n6187), .A2(n6988), .ZN(cv_d[118]) );
NAND2_X2 U6697 ( .A1(cv_q[118]), .A2(n7158), .ZN(n6988) );
NAND2_X2 U6699 ( .A1(cv[118]), .A2(n7134), .ZN(n6990) );
NAND2_X2 U6700 ( .A1(cv_next[118]), .A2(n7149), .ZN(n6989) );
NAND2_X2 U6701 ( .A1(n6189), .A2(n6991), .ZN(cv_d[117]) );
NAND2_X2 U6702 ( .A1(cv_q[117]), .A2(n7158), .ZN(n6991) );
NAND2_X2 U6704 ( .A1(cv[117]), .A2(n7134), .ZN(n6993) );
NAND2_X2 U6705 ( .A1(cv_next[117]), .A2(n7149), .ZN(n6992) );
NAND2_X2 U6706 ( .A1(n6191), .A2(n6994), .ZN(cv_d[116]) );
NAND2_X2 U6707 ( .A1(cv_q[116]), .A2(n7158), .ZN(n6994) );
NAND2_X2 U6709 ( .A1(cv[116]), .A2(n7134), .ZN(n6996) );
NAND2_X2 U6710 ( .A1(cv_next[116]), .A2(n7149), .ZN(n6995) );
NAND2_X2 U6711 ( .A1(n6193), .A2(n6997), .ZN(cv_d[115]) );
NAND2_X2 U6712 ( .A1(cv_q[115]), .A2(n7158), .ZN(n6997) );
NAND2_X2 U6714 ( .A1(cv[115]), .A2(n7134), .ZN(n6999) );
NAND2_X2 U6715 ( .A1(cv_next[115]), .A2(n7149), .ZN(n6998) );
NAND2_X2 U6716 ( .A1(n6195), .A2(n7000), .ZN(cv_d[114]) );
NAND2_X2 U6717 ( .A1(cv_q[114]), .A2(n7158), .ZN(n7000) );
NAND2_X2 U6719 ( .A1(cv[114]), .A2(n7135), .ZN(n7002) );
NAND2_X2 U6720 ( .A1(cv_next[114]), .A2(n7150), .ZN(n7001) );
NAND2_X2 U6721 ( .A1(n6197), .A2(n7003), .ZN(cv_d[113]) );
NAND2_X2 U6722 ( .A1(cv_q[113]), .A2(n7158), .ZN(n7003) );
NAND2_X2 U6724 ( .A1(cv[113]), .A2(n7135), .ZN(n7005) );
NAND2_X2 U6725 ( .A1(cv_next[113]), .A2(n7150), .ZN(n7004) );
NAND2_X2 U6726 ( .A1(n6199), .A2(n7006), .ZN(cv_d[112]) );
NAND2_X2 U6727 ( .A1(cv_q[112]), .A2(n7158), .ZN(n7006) );
NAND2_X2 U6729 ( .A1(cv[112]), .A2(n7135), .ZN(n7008) );
NAND2_X2 U6730 ( .A1(cv_next[112]), .A2(n7150), .ZN(n7007) );
NAND2_X2 U6731 ( .A1(n6201), .A2(n7009), .ZN(cv_d[111]) );
NAND2_X2 U6732 ( .A1(cv_q[111]), .A2(n7158), .ZN(n7009) );
NAND2_X2 U6734 ( .A1(cv[111]), .A2(n7135), .ZN(n7011) );
NAND2_X2 U6735 ( .A1(cv_next[111]), .A2(n7150), .ZN(n7010) );
NAND2_X2 U6736 ( .A1(n6203), .A2(n7012), .ZN(cv_d[110]) );
NAND2_X2 U6737 ( .A1(cv_q[110]), .A2(n7158), .ZN(n7012) );
NAND2_X2 U6739 ( .A1(cv[110]), .A2(n7135), .ZN(n7014) );
NAND2_X2 U6740 ( .A1(cv_next[110]), .A2(n7150), .ZN(n7013) );
NAND2_X2 U6741 ( .A1(n6205), .A2(n7015), .ZN(cv_d[10]) );
NAND2_X2 U6742 ( .A1(cv_q[10]), .A2(n7158), .ZN(n7015) );
NAND2_X2 U6744 ( .A1(cv[10]), .A2(n7135), .ZN(n7017) );
NAND2_X2 U6745 ( .A1(cv_next[10]), .A2(n7150), .ZN(n7016) );
NAND2_X2 U6746 ( .A1(n6207), .A2(n7018), .ZN(cv_d[109]) );
NAND2_X2 U6747 ( .A1(cv_q[109]), .A2(n7158), .ZN(n7018) );
NAND2_X2 U6749 ( .A1(cv[109]), .A2(n7135), .ZN(n7020) );
NAND2_X2 U6750 ( .A1(cv_next[109]), .A2(n7150), .ZN(n7019) );
NAND2_X2 U6751 ( .A1(n6209), .A2(n7021), .ZN(cv_d[108]) );
NAND2_X2 U6752 ( .A1(cv_q[108]), .A2(n7158), .ZN(n7021) );
NAND2_X2 U6754 ( .A1(cv[108]), .A2(n7135), .ZN(n7023) );
NAND2_X2 U6755 ( .A1(cv_next[108]), .A2(n7150), .ZN(n7022) );
NAND2_X2 U6756 ( .A1(n6211), .A2(n7024), .ZN(cv_d[107]) );
NAND2_X2 U6757 ( .A1(cv_q[107]), .A2(n7158), .ZN(n7024) );
NAND2_X2 U6759 ( .A1(cv[107]), .A2(n7135), .ZN(n7026) );
NAND2_X2 U6760 ( .A1(cv_next[107]), .A2(n7150), .ZN(n7025) );
NAND2_X2 U6761 ( .A1(n6213), .A2(n7027), .ZN(cv_d[106]) );
NAND2_X2 U6762 ( .A1(cv_q[106]), .A2(n7158), .ZN(n7027) );
NAND2_X2 U6764 ( .A1(cv[106]), .A2(n7135), .ZN(n7029) );
NAND2_X2 U6765 ( .A1(cv_next[106]), .A2(n7150), .ZN(n7028) );
NAND2_X2 U6766 ( .A1(n6215), .A2(n7030), .ZN(cv_d[105]) );
NAND2_X2 U6767 ( .A1(cv_q[105]), .A2(n7158), .ZN(n7030) );
NAND2_X2 U6769 ( .A1(cv[105]), .A2(n7135), .ZN(n7032) );
NAND2_X2 U6770 ( .A1(cv_next[105]), .A2(n7150), .ZN(n7031) );
NAND2_X2 U6771 ( .A1(n6217), .A2(n7033), .ZN(cv_d[104]) );
NAND2_X2 U6772 ( .A1(cv_q[104]), .A2(n7158), .ZN(n7033) );
NAND2_X2 U6774 ( .A1(cv[104]), .A2(n7136), .ZN(n7035) );
NAND2_X2 U6775 ( .A1(cv_next[104]), .A2(n7151), .ZN(n7034) );
NAND2_X2 U6776 ( .A1(n6219), .A2(n7036), .ZN(cv_d[103]) );
NAND2_X2 U6777 ( .A1(cv_q[103]), .A2(n7158), .ZN(n7036) );
NAND2_X2 U6779 ( .A1(cv[103]), .A2(n7136), .ZN(n7038) );
NAND2_X2 U6780 ( .A1(cv_next[103]), .A2(n7151), .ZN(n7037) );
NAND2_X2 U6781 ( .A1(n6221), .A2(n7039), .ZN(cv_d[102]) );
NAND2_X2 U6782 ( .A1(cv_q[102]), .A2(n7158), .ZN(n7039) );
NAND2_X2 U6784 ( .A1(cv[102]), .A2(n7136), .ZN(n7041) );
NAND2_X2 U6785 ( .A1(cv_next[102]), .A2(n7151), .ZN(n7040) );
NAND2_X2 U6786 ( .A1(n6223), .A2(n7042), .ZN(cv_d[101]) );
NAND2_X2 U6787 ( .A1(cv_q[101]), .A2(n7158), .ZN(n7042) );
NAND2_X2 U6789 ( .A1(cv[101]), .A2(n7136), .ZN(n7044) );
NAND2_X2 U6790 ( .A1(cv_next[101]), .A2(n7151), .ZN(n7043) );
NAND2_X2 U6791 ( .A1(n6225), .A2(n7045), .ZN(cv_d[100]) );
NAND2_X2 U6792 ( .A1(cv_q[100]), .A2(n7158), .ZN(n7045) );
NAND2_X2 U6794 ( .A1(cv[100]), .A2(n7136), .ZN(n7047) );
NAND2_X2 U6795 ( .A1(cv_next[100]), .A2(n7151), .ZN(n7046) );
NAND2_X2 U6796 ( .A1(n6227), .A2(n7048), .ZN(cv_d[0]) );
NAND2_X2 U6797 ( .A1(cv_q[0]), .A2(n7158), .ZN(n7048) );
NAND2_X2 U6799 ( .A1(cv[0]), .A2(n7136), .ZN(n7050) );
NAND2_X2 U6801 ( .A1(cv_next[0]), .A2(n7151), .ZN(n7049) );
NAND2_X2 U6803 ( .A1(state[0]), .A2(n7395), .ZN(busy) );
NAND2_X1 U6818 ( .A1(n7377), .A2(n6865), .ZN(cv_d[155]) );
NAND2_X4 U6819 ( .A1(n7372), .A2(n7373), .ZN(rnd_d[159]) );
INV_X8 U6820 ( .A(n7118), .ZN(n7119) );
NAND2_X4 U6821 ( .A1(sha1_round_wire[151]), .A2(n7159), .ZN(n7340) );
NAND2_X4 U6822 ( .A1(sha1_round_wire[159]), .A2(n7159), .ZN(n7372) );
NAND2_X2 U6823 ( .A1(n7381), .A2(n7340), .ZN(rnd_d[151]) );
NAND2_X2 U6824 ( .A1(sha1_round_wire[157]), .A2(n7159), .ZN(n7364) );
INV_X8 U6825 ( .A(rnd_cnt_q[2]), .ZN(n7118) );
NAND2_X2 U6826 ( .A1(n7356), .A2(n7377), .ZN(rnd_d[155]) );
INV_X1 U6827 ( .A(n7331), .ZN(n7383) );
INV_X1 U6828 ( .A(n7351), .ZN(n7378) );
INV_X1 U6829 ( .A(n7367), .ZN(n7374) );
INV_X1 U6830 ( .A(n7347), .ZN(n7379) );
AND2_X1 U6831 ( .A1(n7049), .A2(n7050), .ZN(n6227) );
AND2_X1 U6832 ( .A1(n6836), .A2(n6837), .ZN(n6085) );
AND2_X1 U6833 ( .A1(n6803), .A2(n6804), .ZN(n6063) );
AND2_X1 U6834 ( .A1(n6770), .A2(n6771), .ZN(n6041) );
AND2_X1 U6835 ( .A1(n6737), .A2(n6738), .ZN(n6019) );
AND2_X1 U6836 ( .A1(n6704), .A2(n6705), .ZN(n5997) );
AND2_X1 U6837 ( .A1(n6671), .A2(n6672), .ZN(n5975) );
AND2_X1 U6838 ( .A1(n6638), .A2(n6639), .ZN(n5953) );
AND2_X1 U6839 ( .A1(n6605), .A2(n6606), .ZN(n5931) );
AND2_X1 U6840 ( .A1(n6570), .A2(n6571), .ZN(n5909) );
AND2_X1 U6841 ( .A1(n7016), .A2(n7017), .ZN(n6205) );
AND2_X1 U6842 ( .A1(n6983), .A2(n6984), .ZN(n6183) );
AND2_X1 U6843 ( .A1(n6950), .A2(n6951), .ZN(n6161) );
AND2_X1 U6844 ( .A1(n6917), .A2(n6918), .ZN(n6139) );
AND2_X1 U6845 ( .A1(n6884), .A2(n6885), .ZN(n6117) );
AND2_X1 U6846 ( .A1(n6851), .A2(n6852), .ZN(n6095) );
AND2_X1 U6847 ( .A1(n6848), .A2(n6849), .ZN(n6093) );
AND2_X1 U6848 ( .A1(n6845), .A2(n6846), .ZN(n6091) );
AND2_X1 U6849 ( .A1(n6842), .A2(n6843), .ZN(n6089) );
AND2_X1 U6850 ( .A1(n6839), .A2(n6840), .ZN(n6087) );
AND2_X1 U6851 ( .A1(n6833), .A2(n6834), .ZN(n6083) );
AND2_X1 U6852 ( .A1(n6830), .A2(n6831), .ZN(n6081) );
AND2_X1 U6853 ( .A1(n6827), .A2(n6828), .ZN(n6079) );
AND2_X1 U6854 ( .A1(n6824), .A2(n6825), .ZN(n6077) );
AND2_X1 U6855 ( .A1(n6821), .A2(n6822), .ZN(n6075) );
AND2_X1 U6856 ( .A1(n6818), .A2(n6819), .ZN(n6073) );
AND2_X1 U6857 ( .A1(n6815), .A2(n6816), .ZN(n6071) );
AND2_X1 U6858 ( .A1(n6812), .A2(n6813), .ZN(n6069) );
AND2_X1 U6859 ( .A1(n6809), .A2(n6810), .ZN(n6067) );
AND2_X1 U6860 ( .A1(n6806), .A2(n6807), .ZN(n6065) );
AND2_X1 U6861 ( .A1(n6800), .A2(n6801), .ZN(n6061) );
AND2_X1 U6862 ( .A1(n6797), .A2(n6798), .ZN(n6059) );
AND2_X1 U6863 ( .A1(n6794), .A2(n6795), .ZN(n6057) );
AND2_X1 U6864 ( .A1(n6791), .A2(n6792), .ZN(n6055) );
AND2_X1 U6865 ( .A1(n6788), .A2(n6789), .ZN(n6053) );
AND2_X1 U6866 ( .A1(n6785), .A2(n6786), .ZN(n6051) );
AND2_X1 U6867 ( .A1(n6782), .A2(n6783), .ZN(n6049) );
AND2_X1 U6868 ( .A1(n6779), .A2(n6780), .ZN(n6047) );
AND2_X1 U6869 ( .A1(n6776), .A2(n6777), .ZN(n6045) );
AND2_X1 U6870 ( .A1(n6773), .A2(n6774), .ZN(n6043) );
AND2_X1 U6871 ( .A1(n6767), .A2(n6768), .ZN(n6039) );
AND2_X1 U6872 ( .A1(n6764), .A2(n6765), .ZN(n6037) );
AND2_X1 U6873 ( .A1(n6761), .A2(n6762), .ZN(n6035) );
AND2_X1 U6874 ( .A1(n6758), .A2(n6759), .ZN(n6033) );
AND2_X1 U6875 ( .A1(n6755), .A2(n6756), .ZN(n6031) );
AND2_X1 U6876 ( .A1(n6752), .A2(n6753), .ZN(n6029) );
AND2_X1 U6877 ( .A1(n6749), .A2(n6750), .ZN(n6027) );
AND2_X1 U6878 ( .A1(n6746), .A2(n6747), .ZN(n6025) );
AND2_X1 U6879 ( .A1(n6743), .A2(n6744), .ZN(n6023) );
AND2_X1 U6880 ( .A1(n6740), .A2(n6741), .ZN(n6021) );
AND2_X1 U6881 ( .A1(n6734), .A2(n6735), .ZN(n6017) );
AND2_X1 U6882 ( .A1(n6731), .A2(n6732), .ZN(n6015) );
AND2_X1 U6883 ( .A1(n6728), .A2(n6729), .ZN(n6013) );
AND2_X1 U6884 ( .A1(n6725), .A2(n6726), .ZN(n6011) );
AND2_X1 U6885 ( .A1(n6722), .A2(n6723), .ZN(n6009) );
AND2_X1 U6886 ( .A1(n6719), .A2(n6720), .ZN(n6007) );
AND2_X1 U6887 ( .A1(n6716), .A2(n6717), .ZN(n6005) );
AND2_X1 U6888 ( .A1(n6713), .A2(n6714), .ZN(n6003) );
AND2_X1 U6889 ( .A1(n6710), .A2(n6711), .ZN(n6001) );
AND2_X1 U6890 ( .A1(n6707), .A2(n6708), .ZN(n5999) );
AND2_X1 U6891 ( .A1(n6701), .A2(n6702), .ZN(n5995) );
AND2_X1 U6892 ( .A1(n6698), .A2(n6699), .ZN(n5993) );
AND2_X1 U6893 ( .A1(n6695), .A2(n6696), .ZN(n5991) );
AND2_X1 U6894 ( .A1(n6692), .A2(n6693), .ZN(n5989) );
AND2_X1 U6895 ( .A1(n6689), .A2(n6690), .ZN(n5987) );
AND2_X1 U6896 ( .A1(n6686), .A2(n6687), .ZN(n5985) );
AND2_X1 U6897 ( .A1(n6683), .A2(n6684), .ZN(n5983) );
AND2_X1 U6898 ( .A1(n6680), .A2(n6681), .ZN(n5981) );
AND2_X1 U6899 ( .A1(n6677), .A2(n6678), .ZN(n5979) );
AND2_X1 U6900 ( .A1(n6674), .A2(n6675), .ZN(n5977) );
AND2_X1 U6901 ( .A1(n6668), .A2(n6669), .ZN(n5973) );
AND2_X1 U6902 ( .A1(n6665), .A2(n6666), .ZN(n5971) );
AND2_X1 U6903 ( .A1(n6662), .A2(n6663), .ZN(n5969) );
AND2_X1 U6904 ( .A1(n6659), .A2(n6660), .ZN(n5967) );
AND2_X1 U6905 ( .A1(n6656), .A2(n6657), .ZN(n5965) );
AND2_X1 U6906 ( .A1(n6653), .A2(n6654), .ZN(n5963) );
AND2_X1 U6907 ( .A1(n6650), .A2(n6651), .ZN(n5961) );
AND2_X1 U6908 ( .A1(n6647), .A2(n6648), .ZN(n5959) );
AND2_X1 U6909 ( .A1(n6644), .A2(n6645), .ZN(n5957) );
AND2_X1 U6910 ( .A1(n6641), .A2(n6642), .ZN(n5955) );
AND2_X1 U6911 ( .A1(n6635), .A2(n6636), .ZN(n5951) );
AND2_X1 U6912 ( .A1(n6632), .A2(n6633), .ZN(n5949) );
AND2_X1 U6913 ( .A1(n6629), .A2(n6630), .ZN(n5947) );
AND2_X1 U6914 ( .A1(n6626), .A2(n6627), .ZN(n5945) );
AND2_X1 U6915 ( .A1(n6623), .A2(n6624), .ZN(n5943) );
AND2_X1 U6916 ( .A1(n6620), .A2(n6621), .ZN(n5941) );
AND2_X1 U6917 ( .A1(n6617), .A2(n6618), .ZN(n5939) );
AND2_X1 U6918 ( .A1(n6614), .A2(n6615), .ZN(n5937) );
AND2_X1 U6919 ( .A1(n6611), .A2(n6612), .ZN(n5935) );
AND2_X1 U6920 ( .A1(n6608), .A2(n6609), .ZN(n5933) );
AND2_X1 U6921 ( .A1(n6602), .A2(n6603), .ZN(n5929) );
AND2_X1 U6922 ( .A1(n6599), .A2(n6600), .ZN(n5927) );
AND2_X1 U6923 ( .A1(n6596), .A2(n6597), .ZN(n5925) );
AND2_X1 U6924 ( .A1(n6593), .A2(n6594), .ZN(n5923) );
AND2_X1 U6925 ( .A1(n6590), .A2(n6591), .ZN(n5921) );
AND2_X1 U6926 ( .A1(n6587), .A2(n6588), .ZN(n5919) );
AND2_X1 U6927 ( .A1(n6584), .A2(n6585), .ZN(n5917) );
AND2_X1 U6928 ( .A1(n6581), .A2(n6582), .ZN(n5915) );
AND2_X1 U6929 ( .A1(n6578), .A2(n6579), .ZN(n5913) );
AND2_X1 U6930 ( .A1(n6575), .A2(n6576), .ZN(n5911) );
AND2_X1 U6931 ( .A1(n7046), .A2(n7047), .ZN(n6225) );
AND2_X1 U6932 ( .A1(n7043), .A2(n7044), .ZN(n6223) );
AND2_X1 U6933 ( .A1(n7040), .A2(n7041), .ZN(n6221) );
AND2_X1 U6934 ( .A1(n7037), .A2(n7038), .ZN(n6219) );
AND2_X1 U6935 ( .A1(n7034), .A2(n7035), .ZN(n6217) );
AND2_X1 U6936 ( .A1(n7031), .A2(n7032), .ZN(n6215) );
AND2_X1 U6937 ( .A1(n7028), .A2(n7029), .ZN(n6213) );
AND2_X1 U6938 ( .A1(n7025), .A2(n7026), .ZN(n6211) );
AND2_X1 U6939 ( .A1(n7022), .A2(n7023), .ZN(n6209) );
AND2_X1 U6940 ( .A1(n7019), .A2(n7020), .ZN(n6207) );
AND2_X1 U6941 ( .A1(n7013), .A2(n7014), .ZN(n6203) );
AND2_X1 U6942 ( .A1(n7010), .A2(n7011), .ZN(n6201) );
AND2_X1 U6943 ( .A1(n7007), .A2(n7008), .ZN(n6199) );
AND2_X1 U6944 ( .A1(n7004), .A2(n7005), .ZN(n6197) );
AND2_X1 U6945 ( .A1(n7001), .A2(n7002), .ZN(n6195) );
AND2_X1 U6946 ( .A1(n6998), .A2(n6999), .ZN(n6193) );
AND2_X1 U6947 ( .A1(n6995), .A2(n6996), .ZN(n6191) );
AND2_X1 U6948 ( .A1(n6992), .A2(n6993), .ZN(n6189) );
AND2_X1 U6949 ( .A1(n6989), .A2(n6990), .ZN(n6187) );
AND2_X1 U6950 ( .A1(n6986), .A2(n6987), .ZN(n6185) );
AND2_X1 U6951 ( .A1(n6980), .A2(n6981), .ZN(n6181) );
AND2_X1 U6952 ( .A1(n6977), .A2(n6978), .ZN(n6179) );
AND2_X1 U6953 ( .A1(n6974), .A2(n6975), .ZN(n6177) );
AND2_X1 U6954 ( .A1(n6971), .A2(n6972), .ZN(n6175) );
AND2_X1 U6955 ( .A1(n6968), .A2(n6969), .ZN(n6173) );
AND2_X1 U6956 ( .A1(n6965), .A2(n6966), .ZN(n6171) );
AND2_X1 U6957 ( .A1(n6962), .A2(n6963), .ZN(n6169) );
AND2_X1 U6958 ( .A1(n6959), .A2(n6960), .ZN(n6167) );
AND2_X1 U6959 ( .A1(n6956), .A2(n6957), .ZN(n6165) );
AND2_X1 U6960 ( .A1(n6953), .A2(n6954), .ZN(n6163) );
AND2_X1 U6961 ( .A1(n6947), .A2(n6948), .ZN(n6159) );
AND2_X1 U6962 ( .A1(n6944), .A2(n6945), .ZN(n6157) );
AND2_X1 U6963 ( .A1(n6941), .A2(n6942), .ZN(n6155) );
AND2_X1 U6964 ( .A1(n6938), .A2(n6939), .ZN(n6153) );
AND2_X1 U6965 ( .A1(n6935), .A2(n6936), .ZN(n6151) );
AND2_X1 U6966 ( .A1(n6932), .A2(n6933), .ZN(n6149) );
AND2_X1 U6967 ( .A1(n6929), .A2(n6930), .ZN(n6147) );
AND2_X1 U6968 ( .A1(n6926), .A2(n6927), .ZN(n6145) );
INV_X8 U6969 ( .A(n7287), .ZN(n7394) );
NAND2_X1 U6970 ( .A1(cv[138]), .A2(n7122), .ZN(n7286) );
NAND2_X1 U6971 ( .A1(n7286), .A2(n7285), .ZN(n7287) );
INV_X8 U6972 ( .A(n7291), .ZN(n7393) );
NAND2_X1 U6973 ( .A1(cv[139]), .A2(n7122), .ZN(n7290) );
NAND2_X1 U6974 ( .A1(n7290), .A2(n7289), .ZN(n7291) );
INV_X8 U6975 ( .A(n7295), .ZN(n7392) );
NAND2_X1 U6976 ( .A1(cv[140]), .A2(n7122), .ZN(n7294) );
NAND2_X1 U6977 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
INV_X8 U6978 ( .A(n7299), .ZN(n7391) );
NAND2_X1 U6979 ( .A1(cv[141]), .A2(n7122), .ZN(n7298) );
NAND2_X1 U6980 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
INV_X8 U6981 ( .A(n7303), .ZN(n7390) );
NAND2_X1 U6982 ( .A1(cv[142]), .A2(n7122), .ZN(n7302) );
NAND2_X1 U6983 ( .A1(n7302), .A2(n7301), .ZN(n7303) );
INV_X8 U6984 ( .A(n7307), .ZN(n7389) );
NAND2_X1 U6985 ( .A1(cv[143]), .A2(n7122), .ZN(n7306) );
NAND2_X1 U6986 ( .A1(n7306), .A2(n7305), .ZN(n7307) );
INV_X8 U6987 ( .A(n7311), .ZN(n7388) );
NAND2_X1 U6988 ( .A1(cv[144]), .A2(n7122), .ZN(n7310) );
NAND2_X1 U6989 ( .A1(n7310), .A2(n7309), .ZN(n7311) );
INV_X8 U6990 ( .A(n7315), .ZN(n7387) );
NAND2_X1 U6991 ( .A1(cv[145]), .A2(n7122), .ZN(n7314) );
NAND2_X1 U6992 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
INV_X8 U6993 ( .A(n7319), .ZN(n7386) );
NAND2_X1 U6994 ( .A1(cv[146]), .A2(n7122), .ZN(n7318) );
NAND2_X1 U6995 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
INV_X8 U6996 ( .A(n7323), .ZN(n7385) );
NAND2_X1 U6997 ( .A1(cv[147]), .A2(n7122), .ZN(n7322) );
NAND2_X1 U6998 ( .A1(n7322), .A2(n7321), .ZN(n7323) );
INV_X8 U6999 ( .A(n7327), .ZN(n7384) );
NAND2_X1 U7000 ( .A1(cv[148]), .A2(n7122), .ZN(n7326) );
NAND2_X1 U7001 ( .A1(n7326), .A2(n7325), .ZN(n7327) );
NAND2_X1 U7002 ( .A1(n7383), .A2(n6886), .ZN(cv_d[149]) );
NAND2_X1 U7003 ( .A1(cv[149]), .A2(n7123), .ZN(n7330) );
NAND2_X1 U7004 ( .A1(n7330), .A2(n7329), .ZN(n7331) );
INV_X8 U7005 ( .A(n7339), .ZN(n7381) );
NAND2_X1 U7006 ( .A1(cv[151]), .A2(n7123), .ZN(n7338) );
NAND2_X1 U7007 ( .A1(n7338), .A2(n7337), .ZN(n7339) );
INV_X8 U7008 ( .A(n7343), .ZN(n7380) );
NAND2_X1 U7009 ( .A1(cv[152]), .A2(n7123), .ZN(n7342) );
NAND2_X1 U7010 ( .A1(n7342), .A2(n7341), .ZN(n7343) );
NAND2_X1 U7011 ( .A1(n7379), .A2(n6871), .ZN(cv_d[153]) );
NAND2_X1 U7012 ( .A1(cv[153]), .A2(n7123), .ZN(n7346) );
NAND2_X1 U7013 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
NAND2_X1 U7014 ( .A1(n7378), .A2(n6868), .ZN(cv_d[154]) );
NAND2_X1 U7015 ( .A1(cv[154]), .A2(n7123), .ZN(n7350) );
NAND2_X1 U7016 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
INV_X1 U7017 ( .A(n7355), .ZN(n7377) );
NAND2_X1 U7018 ( .A1(cv[155]), .A2(n7123), .ZN(n7354) );
NAND2_X1 U7019 ( .A1(n7354), .A2(n7353), .ZN(n7355) );
INV_X8 U7020 ( .A(n7359), .ZN(n7376) );
NAND2_X1 U7021 ( .A1(cv[156]), .A2(n7123), .ZN(n7358) );
NAND2_X1 U7022 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
INV_X8 U7023 ( .A(n7363), .ZN(n7375) );
NAND2_X1 U7024 ( .A1(cv[157]), .A2(n7123), .ZN(n7362) );
NAND2_X1 U7025 ( .A1(n7362), .A2(n7361), .ZN(n7363) );
NAND2_X1 U7026 ( .A1(n7374), .A2(n6856), .ZN(cv_d[158]) );
NAND2_X1 U7027 ( .A1(cv[158]), .A2(n7123), .ZN(n7366) );
NAND2_X1 U7028 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
INV_X1 U7029 ( .A(n5906), .ZN(n7052) );
INV_X4 U7030 ( .A(n7052), .ZN(n7053) );
NAND2_X1 U7031 ( .A1(data_in[0]), .A2(n7228), .ZN(n5906) );
NAND3_X1 U7032 ( .A1(n7053), .A2(n5907), .A3(n5908), .ZN(w_d[0]) );
INV_X1 U7033 ( .A(n5673), .ZN(n7054) );
INV_X4 U7034 ( .A(n7054), .ZN(n7055) );
NAND2_X1 U7035 ( .A1(data_in[1]), .A2(n7228), .ZN(n5673) );
NAND3_X1 U7036 ( .A1(n7055), .A2(n5674), .A3(n5675), .ZN(w_d[1]) );
INV_X1 U7037 ( .A(n5440), .ZN(n7056) );
INV_X4 U7038 ( .A(n7056), .ZN(n7057) );
NAND2_X1 U7039 ( .A1(data_in[2]), .A2(n7229), .ZN(n5440) );
NAND3_X1 U7040 ( .A1(n7057), .A2(n5441), .A3(n5442), .ZN(w_d[2]) );
INV_X1 U7041 ( .A(n5215), .ZN(n7058) );
INV_X4 U7042 ( .A(n7058), .ZN(n7059) );
NAND2_X1 U7043 ( .A1(data_in[3]), .A2(n7229), .ZN(n5215) );
NAND3_X1 U7044 ( .A1(n7059), .A2(n5216), .A3(n5217), .ZN(w_d[3]) );
INV_X1 U7045 ( .A(n4829), .ZN(n7060) );
INV_X4 U7046 ( .A(n7060), .ZN(n7061) );
NAND2_X1 U7047 ( .A1(data_in[4]), .A2(n7229), .ZN(n4829) );
NAND3_X1 U7048 ( .A1(n7061), .A2(n4830), .A3(n4831), .ZN(w_d[4]) );
INV_X1 U7049 ( .A(n4686), .ZN(n7062) );
INV_X4 U7050 ( .A(n7062), .ZN(n7063) );
NAND2_X1 U7051 ( .A1(data_in[5]), .A2(n7229), .ZN(n4686) );
NAND3_X1 U7052 ( .A1(n7063), .A2(n4687), .A3(n4688), .ZN(w_d[5]) );
INV_X1 U7053 ( .A(n4675), .ZN(n7064) );
INV_X4 U7054 ( .A(n7064), .ZN(n7065) );
NAND2_X1 U7055 ( .A1(data_in[6]), .A2(n7229), .ZN(n4675) );
NAND3_X1 U7056 ( .A1(n7065), .A2(n4676), .A3(n4677), .ZN(w_d[6]) );
INV_X1 U7057 ( .A(n4672), .ZN(n7066) );
INV_X4 U7058 ( .A(n7066), .ZN(n7067) );
NAND2_X1 U7059 ( .A1(data_in[7]), .A2(n7229), .ZN(n4672) );
NAND3_X1 U7060 ( .A1(n7067), .A2(n4673), .A3(n4674), .ZN(w_d[7]) );
INV_X1 U7061 ( .A(n4669), .ZN(n7068) );
INV_X4 U7062 ( .A(n7068), .ZN(n7069) );
NAND2_X1 U7063 ( .A1(data_in[8]), .A2(n7229), .ZN(n4669) );
NAND3_X1 U7064 ( .A1(n7069), .A2(n4670), .A3(n4671), .ZN(w_d[8]) );
INV_X1 U7065 ( .A(n4654), .ZN(n7070) );
INV_X4 U7066 ( .A(n7070), .ZN(n7071) );
NAND2_X1 U7067 ( .A1(data_in[9]), .A2(n7227), .ZN(n4654) );
NAND3_X1 U7068 ( .A1(n7071), .A2(n4655), .A3(n4656), .ZN(w_d[9]) );
INV_X1 U7069 ( .A(n5883), .ZN(n7072) );
INV_X4 U7070 ( .A(n7072), .ZN(n7073) );
NAND2_X1 U7071 ( .A1(data_in[10]), .A2(n7227), .ZN(n5883) );
NAND3_X1 U7072 ( .A1(n7073), .A2(n5884), .A3(n5885), .ZN(w_d[10]) );
INV_X1 U7073 ( .A(n5860), .ZN(n7074) );
INV_X4 U7074 ( .A(n7074), .ZN(n7075) );
NAND2_X1 U7075 ( .A1(data_in[11]), .A2(n7227), .ZN(n5860) );
NAND3_X1 U7076 ( .A1(n7075), .A2(n5861), .A3(n5862), .ZN(w_d[11]) );
INV_X1 U7077 ( .A(n5837), .ZN(n7076) );
INV_X4 U7078 ( .A(n7076), .ZN(n7077) );
NAND2_X1 U7079 ( .A1(data_in[12]), .A2(n7227), .ZN(n5837) );
NAND3_X1 U7080 ( .A1(n7077), .A2(n5838), .A3(n5839), .ZN(w_d[12]) );
INV_X1 U7081 ( .A(n5814), .ZN(n7078) );
INV_X4 U7082 ( .A(n7078), .ZN(n7079) );
NAND2_X1 U7083 ( .A1(data_in[13]), .A2(n7227), .ZN(n5814) );
NAND3_X1 U7084 ( .A1(n7079), .A2(n5815), .A3(n5816), .ZN(w_d[13]) );
INV_X1 U7085 ( .A(n5791), .ZN(n7080) );
INV_X4 U7086 ( .A(n7080), .ZN(n7081) );
NAND2_X1 U7087 ( .A1(data_in[14]), .A2(n7227), .ZN(n5791) );
NAND3_X1 U7088 ( .A1(n7081), .A2(n5792), .A3(n5793), .ZN(w_d[14]) );
INV_X1 U7089 ( .A(n5768), .ZN(n7082) );
INV_X4 U7090 ( .A(n7082), .ZN(n7083) );
NAND2_X1 U7091 ( .A1(data_in[15]), .A2(n7227), .ZN(n5768) );
NAND3_X1 U7092 ( .A1(n7083), .A2(n5769), .A3(n5770), .ZN(w_d[15]) );
INV_X1 U7093 ( .A(n5745), .ZN(n7084) );
INV_X4 U7094 ( .A(n7084), .ZN(n7085) );
NAND2_X1 U7095 ( .A1(data_in[16]), .A2(n7227), .ZN(n5745) );
NAND3_X1 U7096 ( .A1(n7085), .A2(n5746), .A3(n5747), .ZN(w_d[16]) );
INV_X1 U7097 ( .A(n5722), .ZN(n7086) );
INV_X4 U7098 ( .A(n7086), .ZN(n7087) );
NAND2_X1 U7099 ( .A1(data_in[17]), .A2(n7227), .ZN(n5722) );
NAND3_X1 U7100 ( .A1(n7087), .A2(n5723), .A3(n5724), .ZN(w_d[17]) );
INV_X1 U7101 ( .A(n5699), .ZN(n7088) );
INV_X4 U7102 ( .A(n7088), .ZN(n7089) );
NAND2_X1 U7103 ( .A1(data_in[18]), .A2(n7227), .ZN(n5699) );
NAND3_X1 U7104 ( .A1(n7089), .A2(n5700), .A3(n5701), .ZN(w_d[18]) );
INV_X1 U7105 ( .A(n5676), .ZN(n7090) );
INV_X4 U7106 ( .A(n7090), .ZN(n7091) );
NAND2_X1 U7107 ( .A1(data_in[19]), .A2(n7227), .ZN(n5676) );
NAND3_X1 U7108 ( .A1(n7091), .A2(n5677), .A3(n5678), .ZN(w_d[19]) );
INV_X1 U7109 ( .A(n5650), .ZN(n7092) );
INV_X4 U7110 ( .A(n7092), .ZN(n7093) );
NAND2_X1 U7111 ( .A1(data_in[20]), .A2(n7228), .ZN(n5650) );
NAND3_X1 U7112 ( .A1(n7093), .A2(n5651), .A3(n5652), .ZN(w_d[20]) );
INV_X1 U7113 ( .A(n5627), .ZN(n7094) );
INV_X4 U7114 ( .A(n7094), .ZN(n7095) );
NAND2_X1 U7115 ( .A1(data_in[21]), .A2(n7228), .ZN(n5627) );
NAND3_X1 U7116 ( .A1(n7095), .A2(n5628), .A3(n5629), .ZN(w_d[21]) );
INV_X1 U7117 ( .A(n5604), .ZN(n7096) );
INV_X4 U7118 ( .A(n7096), .ZN(n7097) );
NAND2_X1 U7119 ( .A1(data_in[22]), .A2(n7228), .ZN(n5604) );
NAND3_X1 U7120 ( .A1(n7097), .A2(n5605), .A3(n5606), .ZN(w_d[22]) );
INV_X1 U7121 ( .A(n5581), .ZN(n7098) );
INV_X4 U7122 ( .A(n7098), .ZN(n7099) );
NAND2_X1 U7123 ( .A1(data_in[23]), .A2(n7228), .ZN(n5581) );
NAND3_X1 U7124 ( .A1(n7099), .A2(n5582), .A3(n5583), .ZN(w_d[23]) );
INV_X1 U7125 ( .A(n5558), .ZN(n7100) );
INV_X4 U7126 ( .A(n7100), .ZN(n7101) );
NAND2_X1 U7127 ( .A1(data_in[24]), .A2(n7228), .ZN(n5558) );
NAND3_X1 U7128 ( .A1(n7101), .A2(n5559), .A3(n5560), .ZN(w_d[24]) );
INV_X1 U7129 ( .A(n5535), .ZN(n7102) );
INV_X4 U7130 ( .A(n7102), .ZN(n7103) );
NAND2_X1 U7131 ( .A1(data_in[25]), .A2(n7228), .ZN(n5535) );
NAND3_X1 U7132 ( .A1(n7103), .A2(n5536), .A3(n5537), .ZN(w_d[25]) );
INV_X1 U7133 ( .A(n5512), .ZN(n7104) );
INV_X4 U7134 ( .A(n7104), .ZN(n7105) );
NAND2_X1 U7135 ( .A1(data_in[26]), .A2(n7228), .ZN(n5512) );
NAND3_X1 U7136 ( .A1(n7105), .A2(n5513), .A3(n5514), .ZN(w_d[26]) );
INV_X1 U7137 ( .A(n5489), .ZN(n7106) );
INV_X4 U7138 ( .A(n7106), .ZN(n7107) );
NAND2_X1 U7139 ( .A1(data_in[27]), .A2(n7228), .ZN(n5489) );
NAND3_X1 U7140 ( .A1(n7107), .A2(n5490), .A3(n5491), .ZN(w_d[27]) );
INV_X1 U7141 ( .A(n5466), .ZN(n7108) );
INV_X4 U7142 ( .A(n7108), .ZN(n7109) );
NAND2_X1 U7143 ( .A1(data_in[28]), .A2(n7228), .ZN(n5466) );
NAND3_X1 U7144 ( .A1(n7109), .A2(n5467), .A3(n5468), .ZN(w_d[28]) );
INV_X1 U7145 ( .A(n5443), .ZN(n7110) );
INV_X4 U7146 ( .A(n7110), .ZN(n7111) );
NAND2_X1 U7147 ( .A1(data_in[29]), .A2(n7229), .ZN(n5443) );
NAND3_X1 U7148 ( .A1(n7111), .A2(n5444), .A3(n5445), .ZN(w_d[29]) );
INV_X1 U7149 ( .A(n5417), .ZN(n7112) );
INV_X4 U7150 ( .A(n7112), .ZN(n7113) );
NAND2_X1 U7151 ( .A1(data_in[30]), .A2(n7229), .ZN(n5417) );
NAND3_X1 U7152 ( .A1(n7113), .A2(n5418), .A3(n5419), .ZN(w_d[30]) );
INV_X1 U7153 ( .A(n5394), .ZN(n7114) );
INV_X4 U7154 ( .A(n7114), .ZN(n7115) );
NAND2_X1 U7155 ( .A1(data_in[31]), .A2(n7229), .ZN(n5394) );
NAND3_X1 U7156 ( .A1(n7115), .A2(n5395), .A3(n5396), .ZN(w_d[31]) );
CLKBUF_X1 U7157 ( .A(start), .Z(n7116) );
CLKBUF_X1 U7158 ( .A(reset), .Z(n7117) );
NOR2_X1 U7159 ( .A1(n7116), .A2(n6243), .ZN(next_state[1]) );
INV_X1 U7160 ( .A(n7371), .ZN(n7373) );
NAND2_X1 U7161 ( .A1(cv[159]), .A2(n7123), .ZN(n7370) );
NAND2_X1 U7162 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
INV_X8 U7163 ( .A(n7335), .ZN(n7382) );
NAND2_X1 U7164 ( .A1(cv[150]), .A2(n7123), .ZN(n7334) );
NAND2_X1 U7165 ( .A1(n7334), .A2(n7333), .ZN(n7335) );
INV_X1 U7166 ( .A(rnd_cnt_q[5]), .ZN(n7398) );
XNOR2_X1 U7167 ( .A(rnd_cnt_q[6]), .B(n6231), .ZN(n6229) );
NAND4_X1 U7168 ( .A1(rnd_cnt_q[6]), .A2(n5038), .A3(n7399), .A4(n7398), .ZN(n6245) );
NAND2_X1 U7169 ( .A1(w[11]), .A2(n7238), .ZN(n4922) );
BUF_X4 U7170 ( .A(n4662), .Z(n7193) );
BUF_X4 U7171 ( .A(n4662), .Z(n7194) );
BUF_X4 U7172 ( .A(n4662), .Z(n7211) );
BUF_X4 U7173 ( .A(n4662), .Z(n7215) );
BUF_X4 U7174 ( .A(n7226), .Z(n7182) );
BUF_X4 U7175 ( .A(n7225), .Z(n7183) );
BUF_X4 U7176 ( .A(n7225), .Z(n7184) );
BUF_X4 U7177 ( .A(n7225), .Z(n7185) );
BUF_X4 U7178 ( .A(n7224), .Z(n7186) );
BUF_X4 U7179 ( .A(n7224), .Z(n7187) );
BUF_X4 U7180 ( .A(n7224), .Z(n7188) );
BUF_X4 U7181 ( .A(n7223), .Z(n7189) );
BUF_X4 U7182 ( .A(n7223), .Z(n7190) );
BUF_X4 U7183 ( .A(n7223), .Z(n7191) );
BUF_X4 U7184 ( .A(n4662), .Z(n7192) );
BUF_X4 U7185 ( .A(n4662), .Z(n7195) );
BUF_X4 U7186 ( .A(n7226), .Z(n7196) );
BUF_X4 U7187 ( .A(n7188), .Z(n7197) );
BUF_X4 U7188 ( .A(n7222), .Z(n7198) );
BUF_X4 U7189 ( .A(n7222), .Z(n7199) );
BUF_X4 U7190 ( .A(n7222), .Z(n7200) );
BUF_X4 U7191 ( .A(n7221), .Z(n7201) );
BUF_X4 U7192 ( .A(n7221), .Z(n7202) );
BUF_X4 U7193 ( .A(n7221), .Z(n7203) );
BUF_X4 U7194 ( .A(n7220), .Z(n7204) );
BUF_X4 U7195 ( .A(n7220), .Z(n7205) );
BUF_X4 U7196 ( .A(n7220), .Z(n7206) );
BUF_X4 U7197 ( .A(n7219), .Z(n7207) );
BUF_X4 U7198 ( .A(n7219), .Z(n7208) );
BUF_X4 U7199 ( .A(n7219), .Z(n7209) );
BUF_X4 U7200 ( .A(n4662), .Z(n7210) );
BUF_X4 U7201 ( .A(n7218), .Z(n7212) );
BUF_X4 U7202 ( .A(n7218), .Z(n7213) );
BUF_X4 U7203 ( .A(n7217), .Z(n7214) );
BUF_X4 U7204 ( .A(n7196), .Z(n7216) );
BUF_X4 U7205 ( .A(n4662), .Z(n7217) );
BUF_X4 U7206 ( .A(n4662), .Z(n7225) );
BUF_X4 U7207 ( .A(n4662), .Z(n7224) );
BUF_X4 U7208 ( .A(n4662), .Z(n7223) );
BUF_X4 U7209 ( .A(n4662), .Z(n7222) );
BUF_X4 U7210 ( .A(n4662), .Z(n7221) );
BUF_X4 U7211 ( .A(n4662), .Z(n7220) );
BUF_X4 U7212 ( .A(n4662), .Z(n7219) );
BUF_X4 U7213 ( .A(n4662), .Z(n7218) );
BUF_X4 U7214 ( .A(n4662), .Z(n7226) );
INV_X4 U7215 ( .A(n7395), .ZN(n7152) );
INV_X4 U7216 ( .A(n7166), .ZN(n7165) );
INV_X4 U7217 ( .A(n7166), .ZN(n7163) );
INV_X4 U7218 ( .A(n7166), .ZN(n7161) );
INV_X4 U7219 ( .A(n7166), .ZN(n7164) );
INV_X4 U7220 ( .A(n7166), .ZN(n7162) );
INV_X4 U7221 ( .A(n7166), .ZN(n7158) );
INV_X4 U7222 ( .A(n7166), .ZN(n7157) );
INV_X4 U7223 ( .A(n7166), .ZN(n7160) );
INV_X4 U7224 ( .A(n7166), .ZN(n7159) );
INV_X4 U7225 ( .A(n7166), .ZN(n7155) );
INV_X4 U7226 ( .A(n7166), .ZN(n7154) );
INV_X4 U7227 ( .A(n7166), .ZN(n7156) );
INV_X4 U7228 ( .A(n7395), .ZN(n7153) );
INV_X4 U7229 ( .A(n6248), .ZN(n7176) );
INV_X4 U7230 ( .A(n6248), .ZN(n7175) );
INV_X4 U7231 ( .A(n6248), .ZN(n7174) );
INV_X4 U7232 ( .A(n6248), .ZN(n7173) );
INV_X4 U7233 ( .A(n6248), .ZN(n7171) );
INV_X4 U7234 ( .A(n6248), .ZN(n7170) );
INV_X4 U7235 ( .A(n6248), .ZN(n7172) );
INV_X4 U7236 ( .A(n6248), .ZN(n7169) );
INV_X4 U7237 ( .A(n7153), .ZN(n7166) );
INV_X4 U7238 ( .A(n6248), .ZN(n7168) );
INV_X4 U7239 ( .A(n6248), .ZN(n7167) );
INV_X4 U7240 ( .A(n7283), .ZN(n7131) );
INV_X4 U7241 ( .A(n7284), .ZN(n7146) );
INV_X4 U7242 ( .A(n7283), .ZN(n7130) );
INV_X4 U7243 ( .A(n7284), .ZN(n7145) );
INV_X4 U7244 ( .A(n7283), .ZN(n7129) );
INV_X4 U7245 ( .A(n7284), .ZN(n7144) );
INV_X4 U7246 ( .A(n7283), .ZN(n7128) );
INV_X4 U7247 ( .A(n7284), .ZN(n7143) );
INV_X4 U7248 ( .A(n7283), .ZN(n7135) );
INV_X4 U7249 ( .A(n7284), .ZN(n7150) );
INV_X4 U7250 ( .A(n7283), .ZN(n7134) );
INV_X4 U7251 ( .A(n7284), .ZN(n7149) );
INV_X4 U7252 ( .A(n7283), .ZN(n7133) );
INV_X4 U7253 ( .A(n7284), .ZN(n7148) );
INV_X4 U7254 ( .A(n7283), .ZN(n7132) );
INV_X4 U7255 ( .A(n7284), .ZN(n7147) );
INV_X4 U7256 ( .A(n7284), .ZN(n7137) );
INV_X4 U7257 ( .A(n7283), .ZN(n7122) );
INV_X4 U7258 ( .A(n7284), .ZN(n7138) );
INV_X4 U7259 ( .A(n7283), .ZN(n7123) );
INV_X4 U7260 ( .A(n7283), .ZN(n7127) );
INV_X4 U7261 ( .A(n7284), .ZN(n7142) );
INV_X4 U7262 ( .A(n7283), .ZN(n7126) );
INV_X4 U7263 ( .A(n7284), .ZN(n7141) );
INV_X4 U7264 ( .A(n7283), .ZN(n7125) );
INV_X4 U7265 ( .A(n7284), .ZN(n7140) );
INV_X4 U7266 ( .A(n7283), .ZN(n7124) );
INV_X4 U7267 ( .A(n7284), .ZN(n7139) );
INV_X4 U7268 ( .A(n7283), .ZN(n7136) );
INV_X4 U7269 ( .A(n7284), .ZN(n7151) );
BUF_X4 U7270 ( .A(n7237), .Z(n7269) );
BUF_X4 U7271 ( .A(n4658), .Z(n7270) );
BUF_X4 U7272 ( .A(n7237), .Z(n7271) );
BUF_X4 U7273 ( .A(n7237), .Z(n7276) );
BUF_X4 U7274 ( .A(n7237), .Z(n7277) );
BUF_X4 U7275 ( .A(n7238), .Z(n7278) );
BUF_X4 U7276 ( .A(n7279), .Z(n7239) );
BUF_X4 U7277 ( .A(n7279), .Z(n7240) );
BUF_X4 U7278 ( .A(n7279), .Z(n7241) );
BUF_X4 U7279 ( .A(n7230), .Z(n7242) );
BUF_X4 U7280 ( .A(n7230), .Z(n7243) );
BUF_X4 U7281 ( .A(n7230), .Z(n7244) );
BUF_X4 U7282 ( .A(n7231), .Z(n7245) );
BUF_X4 U7283 ( .A(n7231), .Z(n7246) );
BUF_X4 U7284 ( .A(n7231), .Z(n7247) );
BUF_X4 U7285 ( .A(n7232), .Z(n7248) );
BUF_X4 U7286 ( .A(n7232), .Z(n7249) );
BUF_X4 U7287 ( .A(n7232), .Z(n7250) );
BUF_X4 U7288 ( .A(n4658), .Z(n7251) );
BUF_X4 U7289 ( .A(n7237), .Z(n7252) );
BUF_X4 U7290 ( .A(n7267), .Z(n7253) );
BUF_X4 U7291 ( .A(n7274), .Z(n7254) );
BUF_X4 U7292 ( .A(n7233), .Z(n7255) );
BUF_X4 U7293 ( .A(n7233), .Z(n7256) );
BUF_X4 U7294 ( .A(n7233), .Z(n7257) );
BUF_X4 U7295 ( .A(n7234), .Z(n7258) );
BUF_X4 U7296 ( .A(n7234), .Z(n7259) );
BUF_X4 U7297 ( .A(n7234), .Z(n7260) );
BUF_X4 U7298 ( .A(n7235), .Z(n7261) );
BUF_X4 U7299 ( .A(n7235), .Z(n7262) );
BUF_X4 U7300 ( .A(n7235), .Z(n7263) );
BUF_X4 U7301 ( .A(n7236), .Z(n7264) );
BUF_X4 U7302 ( .A(n7236), .Z(n7265) );
BUF_X4 U7303 ( .A(n7236), .Z(n7266) );
BUF_X4 U7304 ( .A(n7236), .Z(n7267) );
BUF_X4 U7305 ( .A(n4658), .Z(n7268) );
BUF_X4 U7306 ( .A(n7237), .Z(n7272) );
BUF_X4 U7307 ( .A(n7237), .Z(n7273) );
BUF_X4 U7308 ( .A(n7237), .Z(n7274) );
BUF_X4 U7309 ( .A(n7237), .Z(n7275) );
BUF_X4 U7310 ( .A(n7238), .Z(n7279) );
INV_X4 U7311 ( .A(n7120), .ZN(n7229) );
INV_X4 U7312 ( .A(n7120), .ZN(n7227) );
INV_X4 U7313 ( .A(n7120), .ZN(n7228) );
INV_X4 U7314 ( .A(n7181), .ZN(n7177) );
INV_X4 U7315 ( .A(n7181), .ZN(n7178) );
INV_X4 U7316 ( .A(n7181), .ZN(n7179) );
BUF_X4 U7317 ( .A(n4658), .Z(n7230) );
BUF_X4 U7318 ( .A(n4658), .Z(n7231) );
BUF_X4 U7319 ( .A(n4658), .Z(n7232) );
BUF_X4 U7320 ( .A(n4658), .Z(n7233) );
BUF_X4 U7321 ( .A(n4658), .Z(n7234) );
BUF_X4 U7322 ( .A(n4658), .Z(n7235) );
BUF_X4 U7323 ( .A(n4658), .Z(n7236) );
BUF_X4 U7324 ( .A(n4658), .Z(n7237) );
BUF_X4 U7325 ( .A(n4658), .Z(n7238) );
OR2_X2 U7326 ( .A1(n7403), .A2(n7152), .ZN(n7120) );
NAND3_X2 U7327 ( .A1(n6245), .A2(n7402), .A3(n7152), .ZN(n6230) );
INV_X4 U7328 ( .A(n7121), .ZN(n7180) );
NOR2_X2 U7329 ( .A1(n6233), .A2(n6230), .ZN(rnd_cnt_d[5]) );
NOR2_X2 U7330 ( .A1(n6234), .A2(n6230), .ZN(rnd_cnt_d[4]) );
INV_X4 U7331 ( .A(n7121), .ZN(n7181) );
NOR2_X2 U7332 ( .A1(n7152), .A2(load_in), .ZN(n4658) );
NOR2_X2 U7333 ( .A1(n6230), .A2(rnd_cnt_q[0]), .ZN(rnd_cnt_d[0]) );
AND2_X2 U7334 ( .A1(n5037), .A2(n7403), .ZN(n7121) );
NOR2_X2 U7335 ( .A1(n6244), .A2(n7167), .ZN(n6243) );
NOR2_X2 U7336 ( .A1(n7395), .A2(n6245), .ZN(n6244) );
NAND3_X2 U7337 ( .A1(n6246), .A2(n6230), .A3(n6247), .ZN(next_state[0]) );
NAND3_X2 U7338 ( .A1(n6248), .A2(n7395), .A3(n7116), .ZN(n6246) );
NAND3_X2 U7339 ( .A1(rnd_cnt_q[0]), .A2(n7401), .A3(n7396), .ZN(n6242) );
NOR2_X2 U7340 ( .A1(n6229), .A2(n6230), .ZN(rnd_cnt_d[6]) );
NOR2_X2 U7341 ( .A1(n6232), .A2(n7398), .ZN(n6231) );
NOR2_X2 U7342 ( .A1(n6235), .A2(n6230), .ZN(rnd_cnt_d[3]) );
XNOR2_X1 U7343 ( .A(n6236), .B(rnd_cnt_q[3]), .ZN(n6235) );
INV_X1 U7344 ( .A(n7119), .ZN(n7400) );
INV_X1 U7345 ( .A(rnd_cnt_q[4]), .ZN(n7399) );
NAND2_X1 U7346 ( .A1(n7119), .A2(n6239), .ZN(n6237) );
AND3_X4 U7347 ( .A1(rnd_cnt_q[1]), .A2(rnd_cnt_q[0]), .A3(n7119), .ZN(n6236));
XNOR2_X1 U7348 ( .A(rnd_cnt_q[4]), .B(n5038), .ZN(n6234) );
NAND2_X1 U7349 ( .A1(rnd_cnt_q[4]), .A2(n5038), .ZN(n6232) );
OR4_X1 U7350 ( .A1(n5038), .A2(rnd_cnt_q[4]), .A3(rnd_cnt_q[5]), .A4(rnd_cnt_q[6]), .ZN(n5037) );
OR2_X4 U7351 ( .A1(n7165), .A2(n7229), .ZN(n4662) );
INV_X4 U7352 ( .A(state[0]), .ZN(n7280) );
NAND2_X2 U7353 ( .A1(state[1]), .A2(n7280), .ZN(n6248) );
MUX2_X2 U7354 ( .A(cv_next[0]), .B(N157), .S(n7167), .Z(cv_next_d[0]) );
MUX2_X2 U7355 ( .A(cv_next[1]), .B(N158), .S(n7168), .Z(cv_next_d[1]) );
MUX2_X2 U7356 ( .A(cv_next[2]), .B(N159), .S(n7167), .Z(cv_next_d[2]) );
MUX2_X2 U7357 ( .A(cv_next[3]), .B(N160), .S(n7176), .Z(cv_next_d[3]) );
MUX2_X2 U7358 ( .A(cv_next[4]), .B(N161), .S(n7176), .Z(cv_next_d[4]) );
MUX2_X2 U7359 ( .A(cv_next[5]), .B(N162), .S(n7176), .Z(cv_next_d[5]) );
MUX2_X2 U7360 ( .A(cv_next[6]), .B(N163), .S(n7176), .Z(cv_next_d[6]) );
MUX2_X2 U7361 ( .A(cv_next[7]), .B(N164), .S(n7176), .Z(cv_next_d[7]) );
MUX2_X2 U7362 ( .A(cv_next[8]), .B(N165), .S(n7176), .Z(cv_next_d[8]) );
MUX2_X2 U7363 ( .A(cv_next[9]), .B(N166), .S(n7176), .Z(cv_next_d[9]) );
MUX2_X2 U7364 ( .A(cv_next[10]), .B(N167), .S(n7176), .Z(cv_next_d[10]) );
MUX2_X2 U7365 ( .A(cv_next[11]), .B(N168), .S(n7176), .Z(cv_next_d[11]) );
MUX2_X2 U7366 ( .A(cv_next[12]), .B(N169), .S(n7176), .Z(cv_next_d[12]) );
MUX2_X2 U7367 ( .A(cv_next[13]), .B(N170), .S(n7176), .Z(cv_next_d[13]) );
MUX2_X2 U7368 ( .A(cv_next[14]), .B(N171), .S(n7176), .Z(cv_next_d[14]) );
MUX2_X2 U7369 ( .A(cv_next[15]), .B(N172), .S(n7176), .Z(cv_next_d[15]) );
MUX2_X2 U7370 ( .A(cv_next[16]), .B(N173), .S(n7176), .Z(cv_next_d[16]) );
MUX2_X2 U7371 ( .A(cv_next[17]), .B(N174), .S(n7176), .Z(cv_next_d[17]) );
MUX2_X2 U7372 ( .A(cv_next[18]), .B(N175), .S(n7176), .Z(cv_next_d[18]) );
MUX2_X2 U7373 ( .A(cv_next[19]), .B(N176), .S(n7175), .Z(cv_next_d[19]) );
MUX2_X2 U7374 ( .A(cv_next[20]), .B(N177), .S(n7175), .Z(cv_next_d[20]) );
MUX2_X2 U7375 ( .A(cv_next[21]), .B(N178), .S(n7175), .Z(cv_next_d[21]) );
MUX2_X2 U7376 ( .A(cv_next[22]), .B(N179), .S(n7175), .Z(cv_next_d[22]) );
MUX2_X2 U7377 ( .A(cv_next[23]), .B(N180), .S(n7175), .Z(cv_next_d[23]) );
MUX2_X2 U7378 ( .A(cv_next[24]), .B(N181), .S(n7175), .Z(cv_next_d[24]) );
MUX2_X2 U7379 ( .A(cv_next[25]), .B(N182), .S(n7175), .Z(cv_next_d[25]) );
MUX2_X2 U7380 ( .A(cv_next[26]), .B(N183), .S(n7175), .Z(cv_next_d[26]) );
MUX2_X2 U7381 ( .A(cv_next[27]), .B(N184), .S(n7175), .Z(cv_next_d[27]) );
MUX2_X2 U7382 ( .A(cv_next[28]), .B(N185), .S(n7175), .Z(cv_next_d[28]) );
MUX2_X2 U7383 ( .A(cv_next[29]), .B(N186), .S(n7175), .Z(cv_next_d[29]) );
MUX2_X2 U7384 ( .A(cv_next[30]), .B(N187), .S(n7175), .Z(cv_next_d[30]) );
MUX2_X2 U7385 ( .A(cv_next[31]), .B(N188), .S(n7175), .Z(cv_next_d[31]) );
MUX2_X2 U7386 ( .A(cv_next[32]), .B(N125), .S(n7175), .Z(cv_next_d[32]) );
MUX2_X2 U7387 ( .A(cv_next[33]), .B(N126), .S(n7175), .Z(cv_next_d[33]) );
MUX2_X2 U7388 ( .A(cv_next[34]), .B(N127), .S(n7175), .Z(cv_next_d[34]) );
MUX2_X2 U7389 ( .A(cv_next[35]), .B(N128), .S(n7174), .Z(cv_next_d[35]) );
MUX2_X2 U7390 ( .A(cv_next[36]), .B(N129), .S(n7174), .Z(cv_next_d[36]) );
MUX2_X2 U7391 ( .A(cv_next[37]), .B(N130), .S(n7174), .Z(cv_next_d[37]) );
MUX2_X2 U7392 ( .A(cv_next[38]), .B(N131), .S(n7174), .Z(cv_next_d[38]) );
MUX2_X2 U7393 ( .A(cv_next[39]), .B(N132), .S(n7174), .Z(cv_next_d[39]) );
MUX2_X2 U7394 ( .A(cv_next[40]), .B(N133), .S(n7174), .Z(cv_next_d[40]) );
MUX2_X2 U7395 ( .A(cv_next[41]), .B(N134), .S(n7174), .Z(cv_next_d[41]) );
MUX2_X2 U7396 ( .A(cv_next[42]), .B(N135), .S(n7174), .Z(cv_next_d[42]) );
MUX2_X2 U7397 ( .A(cv_next[43]), .B(N136), .S(n7174), .Z(cv_next_d[43]) );
MUX2_X2 U7398 ( .A(cv_next[44]), .B(N137), .S(n7174), .Z(cv_next_d[44]) );
MUX2_X2 U7399 ( .A(cv_next[45]), .B(N138), .S(n7174), .Z(cv_next_d[45]) );
MUX2_X2 U7400 ( .A(cv_next[46]), .B(N139), .S(n7174), .Z(cv_next_d[46]) );
MUX2_X2 U7401 ( .A(cv_next[47]), .B(N140), .S(n7174), .Z(cv_next_d[47]) );
MUX2_X2 U7402 ( .A(cv_next[48]), .B(N141), .S(n7174), .Z(cv_next_d[48]) );
MUX2_X2 U7403 ( .A(cv_next[49]), .B(N142), .S(n7174), .Z(cv_next_d[49]) );
MUX2_X2 U7404 ( .A(cv_next[50]), .B(N143), .S(n7174), .Z(cv_next_d[50]) );
MUX2_X2 U7405 ( .A(cv_next[51]), .B(N144), .S(n7173), .Z(cv_next_d[51]) );
MUX2_X2 U7406 ( .A(cv_next[52]), .B(N145), .S(n7173), .Z(cv_next_d[52]) );
MUX2_X2 U7407 ( .A(cv_next[53]), .B(N146), .S(n7173), .Z(cv_next_d[53]) );
MUX2_X2 U7408 ( .A(cv_next[54]), .B(N147), .S(n7173), .Z(cv_next_d[54]) );
MUX2_X2 U7409 ( .A(cv_next[55]), .B(N148), .S(n7173), .Z(cv_next_d[55]) );
MUX2_X2 U7410 ( .A(cv_next[56]), .B(N149), .S(n7173), .Z(cv_next_d[56]) );
MUX2_X2 U7411 ( .A(cv_next[57]), .B(N150), .S(n7173), .Z(cv_next_d[57]) );
MUX2_X2 U7412 ( .A(cv_next[58]), .B(N151), .S(n7173), .Z(cv_next_d[58]) );
MUX2_X2 U7413 ( .A(cv_next[59]), .B(N152), .S(n7173), .Z(cv_next_d[59]) );
MUX2_X2 U7414 ( .A(cv_next[60]), .B(N153), .S(n7173), .Z(cv_next_d[60]) );
MUX2_X2 U7415 ( .A(cv_next[61]), .B(N154), .S(n7173), .Z(cv_next_d[61]) );
MUX2_X2 U7416 ( .A(cv_next[62]), .B(N155), .S(n7173), .Z(cv_next_d[62]) );
MUX2_X2 U7417 ( .A(cv_next[63]), .B(N156), .S(n7173), .Z(cv_next_d[63]) );
MUX2_X2 U7418 ( .A(cv_next[64]), .B(N93), .S(n7173), .Z(cv_next_d[64]) );
MUX2_X2 U7419 ( .A(cv_next[65]), .B(N94), .S(n7173), .Z(cv_next_d[65]) );
MUX2_X2 U7420 ( .A(cv_next[66]), .B(N95), .S(n7173), .Z(cv_next_d[66]) );
MUX2_X2 U7421 ( .A(cv_next[67]), .B(N96), .S(n7172), .Z(cv_next_d[67]) );
MUX2_X2 U7422 ( .A(cv_next[68]), .B(N97), .S(n7172), .Z(cv_next_d[68]) );
MUX2_X2 U7423 ( .A(cv_next[69]), .B(N98), .S(n7172), .Z(cv_next_d[69]) );
MUX2_X2 U7424 ( .A(cv_next[70]), .B(N99), .S(n7172), .Z(cv_next_d[70]) );
MUX2_X2 U7425 ( .A(cv_next[71]), .B(N100), .S(n7172), .Z(cv_next_d[71]) );
MUX2_X2 U7426 ( .A(cv_next[72]), .B(N101), .S(n7172), .Z(cv_next_d[72]) );
MUX2_X2 U7427 ( .A(cv_next[73]), .B(N102), .S(n7172), .Z(cv_next_d[73]) );
MUX2_X2 U7428 ( .A(cv_next[74]), .B(N103), .S(n7172), .Z(cv_next_d[74]) );
MUX2_X2 U7429 ( .A(cv_next[75]), .B(N104), .S(n7172), .Z(cv_next_d[75]) );
MUX2_X2 U7430 ( .A(cv_next[76]), .B(N105), .S(n7172), .Z(cv_next_d[76]) );
MUX2_X2 U7431 ( .A(cv_next[77]), .B(N106), .S(n7172), .Z(cv_next_d[77]) );
MUX2_X2 U7432 ( .A(cv_next[78]), .B(N107), .S(n7172), .Z(cv_next_d[78]) );
MUX2_X2 U7433 ( .A(cv_next[79]), .B(N108), .S(n7172), .Z(cv_next_d[79]) );
MUX2_X2 U7434 ( .A(cv_next[80]), .B(N109), .S(n7172), .Z(cv_next_d[80]) );
MUX2_X2 U7435 ( .A(cv_next[81]), .B(N110), .S(n7172), .Z(cv_next_d[81]) );
MUX2_X2 U7436 ( .A(cv_next[82]), .B(N111), .S(n7171), .Z(cv_next_d[82]) );
MUX2_X2 U7437 ( .A(cv_next[83]), .B(N112), .S(n7171), .Z(cv_next_d[83]) );
MUX2_X2 U7438 ( .A(cv_next[84]), .B(N113), .S(n7171), .Z(cv_next_d[84]) );
MUX2_X2 U7439 ( .A(cv_next[85]), .B(N114), .S(n7171), .Z(cv_next_d[85]) );
MUX2_X2 U7440 ( .A(cv_next[86]), .B(N115), .S(n7171), .Z(cv_next_d[86]) );
MUX2_X2 U7441 ( .A(cv_next[87]), .B(N116), .S(n7171), .Z(cv_next_d[87]) );
MUX2_X2 U7442 ( .A(cv_next[88]), .B(N117), .S(n7171), .Z(cv_next_d[88]) );
MUX2_X2 U7443 ( .A(cv_next[89]), .B(N118), .S(n7171), .Z(cv_next_d[89]) );
MUX2_X2 U7444 ( .A(cv_next[90]), .B(N119), .S(n7171), .Z(cv_next_d[90]) );
MUX2_X2 U7445 ( .A(cv_next[91]), .B(N120), .S(n7171), .Z(cv_next_d[91]) );
MUX2_X2 U7446 ( .A(cv_next[92]), .B(N121), .S(n7171), .Z(cv_next_d[92]) );
MUX2_X2 U7447 ( .A(cv_next[93]), .B(N122), .S(n7171), .Z(cv_next_d[93]) );
MUX2_X2 U7448 ( .A(cv_next[94]), .B(N123), .S(n7171), .Z(cv_next_d[94]) );
MUX2_X2 U7449 ( .A(cv_next[95]), .B(N124), .S(n7171), .Z(cv_next_d[95]) );
MUX2_X2 U7450 ( .A(cv_next[96]), .B(N61), .S(n7171), .Z(cv_next_d[96]) );
MUX2_X2 U7451 ( .A(cv_next[97]), .B(N62), .S(n7171), .Z(cv_next_d[97]) );
MUX2_X2 U7452 ( .A(cv_next[98]), .B(N63), .S(n7170), .Z(cv_next_d[98]) );
MUX2_X2 U7453 ( .A(cv_next[99]), .B(N64), .S(n7170), .Z(cv_next_d[99]) );
MUX2_X2 U7454 ( .A(cv_next[100]), .B(N65), .S(n7170), .Z(cv_next_d[100]) );
MUX2_X2 U7455 ( .A(cv_next[101]), .B(N66), .S(n7170), .Z(cv_next_d[101]) );
MUX2_X2 U7456 ( .A(cv_next[102]), .B(N67), .S(n7170), .Z(cv_next_d[102]) );
MUX2_X2 U7457 ( .A(cv_next[103]), .B(N68), .S(n7170), .Z(cv_next_d[103]) );
MUX2_X2 U7458 ( .A(cv_next[104]), .B(N69), .S(n7170), .Z(cv_next_d[104]) );
MUX2_X2 U7459 ( .A(cv_next[105]), .B(N70), .S(n7170), .Z(cv_next_d[105]) );
MUX2_X2 U7460 ( .A(cv_next[106]), .B(N71), .S(n7170), .Z(cv_next_d[106]) );
MUX2_X2 U7461 ( .A(cv_next[107]), .B(N72), .S(n7170), .Z(cv_next_d[107]) );
MUX2_X2 U7462 ( .A(cv_next[108]), .B(N73), .S(n7170), .Z(cv_next_d[108]) );
MUX2_X2 U7463 ( .A(cv_next[109]), .B(N74), .S(n7170), .Z(cv_next_d[109]) );
MUX2_X2 U7464 ( .A(cv_next[110]), .B(N75), .S(n7170), .Z(cv_next_d[110]) );
MUX2_X2 U7465 ( .A(cv_next[111]), .B(N76), .S(n7170), .Z(cv_next_d[111]) );
MUX2_X2 U7466 ( .A(cv_next[112]), .B(N77), .S(n7170), .Z(cv_next_d[112]) );
MUX2_X2 U7467 ( .A(cv_next[113]), .B(N78), .S(n7170), .Z(cv_next_d[113]) );
MUX2_X2 U7468 ( .A(cv_next[114]), .B(N79), .S(n7169), .Z(cv_next_d[114]) );
MUX2_X2 U7469 ( .A(cv_next[115]), .B(N80), .S(n7169), .Z(cv_next_d[115]) );
MUX2_X2 U7470 ( .A(cv_next[116]), .B(N81), .S(n7169), .Z(cv_next_d[116]) );
MUX2_X2 U7471 ( .A(cv_next[117]), .B(N82), .S(n7169), .Z(cv_next_d[117]) );
MUX2_X2 U7472 ( .A(cv_next[118]), .B(N83), .S(n7169), .Z(cv_next_d[118]) );
MUX2_X2 U7473 ( .A(cv_next[119]), .B(N84), .S(n7169), .Z(cv_next_d[119]) );
MUX2_X2 U7474 ( .A(cv_next[120]), .B(N85), .S(n7169), .Z(cv_next_d[120]) );
MUX2_X2 U7475 ( .A(cv_next[121]), .B(N86), .S(n7172), .Z(cv_next_d[121]) );
MUX2_X2 U7476 ( .A(cv_next[122]), .B(N87), .S(n7169), .Z(cv_next_d[122]) );
MUX2_X2 U7477 ( .A(cv_next[123]), .B(N88), .S(n7169), .Z(cv_next_d[123]) );
MUX2_X2 U7478 ( .A(cv_next[124]), .B(N89), .S(n7169), .Z(cv_next_d[124]) );
MUX2_X2 U7479 ( .A(cv_next[125]), .B(N90), .S(n7169), .Z(cv_next_d[125]) );
MUX2_X2 U7480 ( .A(cv_next[126]), .B(N91), .S(n7169), .Z(cv_next_d[126]) );
MUX2_X2 U7481 ( .A(cv_next[127]), .B(N92), .S(n7169), .Z(cv_next_d[127]) );
MUX2_X2 U7482 ( .A(cv_next[128]), .B(N29), .S(n7169), .Z(cv_next_d[128]) );
MUX2_X2 U7483 ( .A(cv_next[129]), .B(N30), .S(n7169), .Z(cv_next_d[129]) );
MUX2_X2 U7484 ( .A(cv_next[130]), .B(N31), .S(n7169), .Z(cv_next_d[130]) );
MUX2_X2 U7485 ( .A(cv_next[131]), .B(N32), .S(n7168), .Z(cv_next_d[131]) );
MUX2_X2 U7486 ( .A(cv_next[132]), .B(N33), .S(n7168), .Z(cv_next_d[132]) );
MUX2_X2 U7487 ( .A(cv_next[133]), .B(N34), .S(n7168), .Z(cv_next_d[133]) );
MUX2_X2 U7488 ( .A(cv_next[134]), .B(N35), .S(n7168), .Z(cv_next_d[134]) );
MUX2_X2 U7489 ( .A(cv_next[135]), .B(N36), .S(n7168), .Z(cv_next_d[135]) );
MUX2_X2 U7490 ( .A(cv_next[136]), .B(N37), .S(n7168), .Z(cv_next_d[136]) );
MUX2_X2 U7491 ( .A(cv_next[137]), .B(N38), .S(n7168), .Z(cv_next_d[137]) );
MUX2_X2 U7492 ( .A(cv_next[138]), .B(N39), .S(n7168), .Z(cv_next_d[138]) );
MUX2_X2 U7493 ( .A(cv_next[139]), .B(N40), .S(n7168), .Z(cv_next_d[139]) );
MUX2_X2 U7494 ( .A(cv_next[140]), .B(N41), .S(n7168), .Z(cv_next_d[140]) );
MUX2_X2 U7495 ( .A(cv_next[141]), .B(N42), .S(n7168), .Z(cv_next_d[141]) );
MUX2_X2 U7496 ( .A(cv_next[142]), .B(N43), .S(n7168), .Z(cv_next_d[142]) );
MUX2_X2 U7497 ( .A(cv_next[143]), .B(N44), .S(n7168), .Z(cv_next_d[143]) );
MUX2_X2 U7498 ( .A(cv_next[144]), .B(N45), .S(n7168), .Z(cv_next_d[144]) );
MUX2_X2 U7499 ( .A(cv_next[145]), .B(N46), .S(n7168), .Z(cv_next_d[145]) );
MUX2_X2 U7500 ( .A(cv_next[146]), .B(N47), .S(n7168), .Z(cv_next_d[146]) );
MUX2_X2 U7501 ( .A(cv_next[147]), .B(N48), .S(n7167), .Z(cv_next_d[147]) );
MUX2_X2 U7502 ( .A(cv_next[148]), .B(N49), .S(n7167), .Z(cv_next_d[148]) );
MUX2_X2 U7503 ( .A(cv_next[149]), .B(N50), .S(n7167), .Z(cv_next_d[149]) );
MUX2_X2 U7504 ( .A(cv_next[150]), .B(N51), .S(n7167), .Z(cv_next_d[150]) );
MUX2_X2 U7505 ( .A(cv_next[151]), .B(N52), .S(n7167), .Z(cv_next_d[151]) );
MUX2_X2 U7506 ( .A(cv_next[152]), .B(N53), .S(n7167), .Z(cv_next_d[152]) );
MUX2_X2 U7507 ( .A(cv_next[153]), .B(N54), .S(n7167), .Z(cv_next_d[153]) );
MUX2_X2 U7508 ( .A(cv_next[154]), .B(N55), .S(n7167), .Z(cv_next_d[154]) );
MUX2_X2 U7509 ( .A(cv_next[155]), .B(N56), .S(n7167), .Z(cv_next_d[155]) );
MUX2_X2 U7510 ( .A(cv_next[156]), .B(N57), .S(n7167), .Z(cv_next_d[156]) );
MUX2_X2 U7511 ( .A(cv_next[157]), .B(N58), .S(n7167), .Z(cv_next_d[157]) );
MUX2_X2 U7512 ( .A(cv_next[158]), .B(N59), .S(n7167), .Z(cv_next_d[158]) );
MUX2_X2 U7513 ( .A(cv_next[159]), .B(N60), .S(n7167), .Z(cv_next_d[159]) );
INV_X4 U7514 ( .A(state[1]), .ZN(n7281) );
NAND2_X2 U7515 ( .A1(state[0]), .A2(n7281), .ZN(n7395) );
INV_X4 U7516 ( .A(use_prev_cv), .ZN(n7282) );
NAND2_X2 U7517 ( .A1(n7395), .A2(n7282), .ZN(n7283) );
NAND2_X2 U7518 ( .A1(use_prev_cv), .A2(n7395), .ZN(n7284) );
NAND2_X2 U7519 ( .A1(cv_next[138]), .A2(n7137), .ZN(n7285) );
NAND2_X2 U7520 ( .A1(sha1_round_wire[138]), .A2(n7152), .ZN(n7288) );
NAND2_X2 U7521 ( .A1(n7394), .A2(n7288), .ZN(rnd_d[138]) );
NAND2_X2 U7522 ( .A1(cv_next[139]), .A2(n7137), .ZN(n7289) );
NAND2_X2 U7523 ( .A1(sha1_round_wire[139]), .A2(n7162), .ZN(n7292) );
NAND2_X2 U7524 ( .A1(n7393), .A2(n7292), .ZN(rnd_d[139]) );
NAND2_X2 U7525 ( .A1(cv_next[140]), .A2(n7137), .ZN(n7293) );
NAND2_X2 U7526 ( .A1(sha1_round_wire[140]), .A2(n7158), .ZN(n7296) );
NAND2_X2 U7527 ( .A1(n7392), .A2(n7296), .ZN(rnd_d[140]) );
NAND2_X2 U7528 ( .A1(cv_next[141]), .A2(n7137), .ZN(n7297) );
NAND2_X2 U7529 ( .A1(sha1_round_wire[141]), .A2(n7158), .ZN(n7300) );
NAND2_X2 U7530 ( .A1(n7391), .A2(n7300), .ZN(rnd_d[141]) );
NAND2_X2 U7531 ( .A1(cv_next[142]), .A2(n7137), .ZN(n7301) );
NAND2_X2 U7532 ( .A1(sha1_round_wire[142]), .A2(n7158), .ZN(n7304) );
NAND2_X2 U7533 ( .A1(n7390), .A2(n7304), .ZN(rnd_d[142]) );
NAND2_X2 U7534 ( .A1(cv_next[143]), .A2(n7137), .ZN(n7305) );
NAND2_X2 U7535 ( .A1(sha1_round_wire[143]), .A2(n7158), .ZN(n7308) );
NAND2_X2 U7536 ( .A1(n7389), .A2(n7308), .ZN(rnd_d[143]) );
NAND2_X2 U7537 ( .A1(cv_next[144]), .A2(n7137), .ZN(n7309) );
NAND2_X2 U7538 ( .A1(sha1_round_wire[144]), .A2(n7158), .ZN(n7312) );
NAND2_X2 U7539 ( .A1(n7388), .A2(n7312), .ZN(rnd_d[144]) );
NAND2_X2 U7540 ( .A1(cv_next[145]), .A2(n7137), .ZN(n7313) );
NAND2_X2 U7541 ( .A1(sha1_round_wire[145]), .A2(n7158), .ZN(n7316) );
NAND2_X2 U7542 ( .A1(n7387), .A2(n7316), .ZN(rnd_d[145]) );
NAND2_X2 U7543 ( .A1(cv_next[146]), .A2(n7137), .ZN(n7317) );
NAND2_X2 U7544 ( .A1(sha1_round_wire[146]), .A2(n7159), .ZN(n7320) );
NAND2_X2 U7545 ( .A1(n7386), .A2(n7320), .ZN(rnd_d[146]) );
NAND2_X2 U7546 ( .A1(cv_next[147]), .A2(n7137), .ZN(n7321) );
NAND2_X2 U7547 ( .A1(sha1_round_wire[147]), .A2(n7159), .ZN(n7324) );
NAND2_X2 U7548 ( .A1(n7385), .A2(n7324), .ZN(rnd_d[147]) );
NAND2_X2 U7549 ( .A1(cv_next[148]), .A2(n7137), .ZN(n7325) );
NAND2_X2 U7550 ( .A1(sha1_round_wire[148]), .A2(n7159), .ZN(n7328) );
NAND2_X2 U7551 ( .A1(n7384), .A2(n7328), .ZN(rnd_d[148]) );
NAND2_X2 U7552 ( .A1(cv_next[149]), .A2(n7138), .ZN(n7329) );
NAND2_X2 U7553 ( .A1(sha1_round_wire[149]), .A2(n7159), .ZN(n7332) );
NAND2_X2 U7554 ( .A1(n7332), .A2(n7383), .ZN(rnd_d[149]) );
NAND2_X2 U7555 ( .A1(cv_next[150]), .A2(n7138), .ZN(n7333) );
NAND2_X2 U7556 ( .A1(sha1_round_wire[150]), .A2(n7159), .ZN(n7336) );
NAND2_X2 U7557 ( .A1(n7382), .A2(n7336), .ZN(rnd_d[150]) );
NAND2_X2 U7558 ( .A1(cv_next[151]), .A2(n7138), .ZN(n7337) );
NAND2_X2 U7559 ( .A1(cv_next[152]), .A2(n7138), .ZN(n7341) );
NAND2_X2 U7560 ( .A1(sha1_round_wire[152]), .A2(n7159), .ZN(n7344) );
NAND2_X2 U7561 ( .A1(n7380), .A2(n7344), .ZN(rnd_d[152]) );
NAND2_X2 U7562 ( .A1(cv_next[153]), .A2(n7138), .ZN(n7345) );
NAND2_X2 U7563 ( .A1(sha1_round_wire[153]), .A2(n7159), .ZN(n7348) );
NAND2_X2 U7564 ( .A1(n7348), .A2(n7379), .ZN(rnd_d[153]) );
NAND2_X2 U7565 ( .A1(cv_next[154]), .A2(n7138), .ZN(n7349) );
NAND2_X2 U7566 ( .A1(sha1_round_wire[154]), .A2(n7159), .ZN(n7352) );
NAND2_X2 U7567 ( .A1(n7352), .A2(n7378), .ZN(rnd_d[154]) );
NAND2_X2 U7568 ( .A1(cv_next[155]), .A2(n7138), .ZN(n7353) );
NAND2_X2 U7569 ( .A1(sha1_round_wire[155]), .A2(n7159), .ZN(n7356) );
NAND2_X2 U7570 ( .A1(cv_next[156]), .A2(n7138), .ZN(n7357) );
NAND2_X2 U7571 ( .A1(sha1_round_wire[156]), .A2(n7159), .ZN(n7360) );
NAND2_X2 U7572 ( .A1(n7376), .A2(n7360), .ZN(rnd_d[156]) );
NAND2_X2 U7573 ( .A1(cv_next[157]), .A2(n7138), .ZN(n7361) );
NAND2_X2 U7574 ( .A1(n7375), .A2(n7364), .ZN(rnd_d[157]) );
NAND2_X2 U7575 ( .A1(cv_next[158]), .A2(n7138), .ZN(n7365) );
NAND2_X2 U7576 ( .A1(sha1_round_wire[158]), .A2(n7159), .ZN(n7368) );
NAND2_X2 U7577 ( .A1(n7368), .A2(n7374), .ZN(rnd_d[158]) );
NAND2_X2 U7578 ( .A1(cv_next[159]), .A2(n7138), .ZN(n7369) );
INV_X4 U7579 ( .A(n6230), .ZN(n7396) );
INV_X4 U7580 ( .A(rnd_cnt_d[0]), .ZN(n7397) );
INV_X4 U7581 ( .A(rnd_cnt_q[1]), .ZN(n7401) );
INV_X4 U7582 ( .A(n7116), .ZN(n7402) );
INV_X4 U7583 ( .A(load_in), .ZN(n7403) );
NAND2_X2 _sha1_round_U575  ( .A1(_sha1_round_n3200 ), .A2(_sha1_round_n821 ),.ZN(_sha1_round_k[13] ) );
INV_X4 _sha1_round_U574  ( .A(_sha1_round_k_23 ), .ZN(_sha1_round_n821 ) );
NAND2_X2 _sha1_round_U573  ( .A1(_sha1_round_n819 ), .A2(_sha1_round_n510 ),.ZN(_sha1_round_k_23 ) );
INV_X4 _sha1_round_U572  ( .A(_sha1_round_n2 ), .ZN(_sha1_round_n818 ) );
NAND2_X2 _sha1_round_U571  ( .A1(rnd_q[32]), .A2(_sha1_round_n812 ), .ZN(_sha1_round_n813 ) );
NAND2_X2 _sha1_round_U570  ( .A1(_sha1_round_n811 ), .A2(_sha1_round_n810 ),.ZN(_sha1_round_n812 ) );
NAND2_X2 _sha1_round_U569  ( .A1(_sha1_round_n808 ), .A2(_sha1_round_n807 ),.ZN(_sha1_round_n809 ) );
INV_X4 _sha1_round_U568  ( .A(rnd_q[64]), .ZN(_sha1_round_n807 ) );
NAND2_X2 _sha1_round_U567  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n808 ),.ZN(_sha1_round_n811 ) );
INV_X4 _sha1_round_U566  ( .A(rnd_q[32]), .ZN(_sha1_round_n804 ) );
INV_X4 _sha1_round_U565  ( .A(_sha1_round_n806 ), .ZN(_sha1_round_n805 ) );
XOR2_X2 _sha1_round_U564  ( .A(_sha1_round_n808 ), .B(rnd_q[64]), .Z(_sha1_round_n806 ) );
INV_X4 _sha1_round_U563  ( .A(rnd_q[96]), .ZN(_sha1_round_n808 ) );
NAND2_X2 _sha1_round_U562  ( .A1(_sha1_round_n798 ), .A2(_sha1_round_n797 ),.ZN(_sha1_round_n799 ) );
NAND2_X2 _sha1_round_U561  ( .A1(_sha1_round_n795 ), .A2(_sha1_round_n794 ),.ZN(_sha1_round_n796 ) );
INV_X4 _sha1_round_U560  ( .A(rnd_q[65]), .ZN(_sha1_round_n794 ) );
NAND2_X2 _sha1_round_U559  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n795 ),.ZN(_sha1_round_n798 ) );
INV_X4 _sha1_round_U558  ( .A(_sha1_round_n793 ), .ZN(_sha1_round_n792 ) );
XOR2_X2 _sha1_round_U557  ( .A(_sha1_round_n795 ), .B(rnd_q[65]), .Z(_sha1_round_n793 ) );
INV_X4 _sha1_round_U556  ( .A(rnd_q[97]), .ZN(_sha1_round_n795 ) );
NAND2_X2 _sha1_round_U555  ( .A1(rnd_q[34]), .A2(_sha1_round_n786 ), .ZN(_sha1_round_n787 ) );
NAND2_X2 _sha1_round_U554  ( .A1(_sha1_round_n785 ), .A2(_sha1_round_n784 ),.ZN(_sha1_round_n786 ) );
NAND2_X2 _sha1_round_U553  ( .A1(_sha1_round_n782 ), .A2(_sha1_round_n781 ),.ZN(_sha1_round_n783 ) );
INV_X4 _sha1_round_U552  ( .A(rnd_q[66]), .ZN(_sha1_round_n781 ) );
NAND2_X2 _sha1_round_U551  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n782 ),.ZN(_sha1_round_n785 ) );
INV_X4 _sha1_round_U550  ( .A(rnd_q[34]), .ZN(_sha1_round_n778 ) );
INV_X4 _sha1_round_U549  ( .A(_sha1_round_n780 ), .ZN(_sha1_round_n779 ) );
XOR2_X2 _sha1_round_U548  ( .A(_sha1_round_n782 ), .B(rnd_q[66]), .Z(_sha1_round_n780 ) );
INV_X4 _sha1_round_U547  ( .A(rnd_q[98]), .ZN(_sha1_round_n782 ) );
NAND2_X2 _sha1_round_U546  ( .A1(_sha1_round_n772 ), .A2(_sha1_round_n771 ),.ZN(_sha1_round_n773 ) );
NAND2_X2 _sha1_round_U545  ( .A1(_sha1_round_n769 ), .A2(_sha1_round_n768 ),.ZN(_sha1_round_n770 ) );
INV_X4 _sha1_round_U544  ( .A(rnd_q[67]), .ZN(_sha1_round_n768 ) );
NAND2_X2 _sha1_round_U543  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n769 ),.ZN(_sha1_round_n772 ) );
INV_X4 _sha1_round_U542  ( .A(rnd_q[35]), .ZN(_sha1_round_n764 ) );
INV_X4 _sha1_round_U541  ( .A(_sha1_round_n766 ), .ZN(_sha1_round_n765 ) );
XOR2_X2 _sha1_round_U540  ( .A(_sha1_round_n769 ), .B(rnd_q[67]), .Z(_sha1_round_n766 ) );
INV_X4 _sha1_round_U539  ( .A(rnd_q[99]), .ZN(_sha1_round_n769 ) );
MUX2_X2 _sha1_round_U538  ( .A(_sha1_round_n761 ), .B(_sha1_round_n760 ),.S(rnd_q[36]), .Z(_sha1_round_n762 ) );
NOR3_X2 _sha1_round_U537  ( .A1(_sha1_round_n759 ), .A2(_sha1_round_n758 ),.A3(_sha1_round_n757 ), .ZN(_sha1_round_n760 ) );
NOR2_X2 _sha1_round_U536  ( .A1(_sha1_round_n755 ), .A2(_sha1_round_n3180 ),.ZN(_sha1_round_n758 ) );
NOR2_X2 _sha1_round_U535  ( .A1(rnd_q[68]), .A2(rnd_q[100]), .ZN(_sha1_round_n755 ) );
NOR2_X2 _sha1_round_U534  ( .A1(rnd_q[100]), .A2(_sha1_round_n510 ), .ZN(_sha1_round_n759 ) );
NAND2_X2 _sha1_round_U533  ( .A1(_sha1_round_n374 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n761 ) );
NAND3_X2 _sha1_round_U532  ( .A1(rnd_q[68]), .A2(rnd_q[100]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n763 ) );
NOR2_X2 _sha1_round_U531  ( .A1(rnd_q[69]), .A2(rnd_q[101]), .ZN(_sha1_round_n750 ) );
NAND3_X2 _sha1_round_U530  ( .A1(rnd_q[69]), .A2(rnd_q[101]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n754 ) );
NOR2_X2 _sha1_round_U529  ( .A1(rnd_q[70]), .A2(rnd_q[102]), .ZN(_sha1_round_n745 ) );
NAND3_X2 _sha1_round_U528  ( .A1(rnd_q[70]), .A2(rnd_q[102]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n749 ) );
NOR3_X2 _sha1_round_U527  ( .A1(_sha1_round_n740 ), .A2(_sha1_round_n739 ),.A3(_sha1_round_n738 ), .ZN(_sha1_round_n741 ) );
NOR2_X2 _sha1_round_U526  ( .A1(_sha1_round_n737 ), .A2(_sha1_round_n514 ),.ZN(_sha1_round_n739 ) );
NOR2_X2 _sha1_round_U525  ( .A1(rnd_q[71]), .A2(rnd_q[103]), .ZN(_sha1_round_n737 ) );
NOR2_X2 _sha1_round_U524  ( .A1(rnd_q[103]), .A2(_sha1_round_n510 ), .ZN(_sha1_round_n740 ) );
NAND3_X2 _sha1_round_U523  ( .A1(rnd_q[71]), .A2(rnd_q[103]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n744 ) );
NOR2_X2 _sha1_round_U522  ( .A1(_sha1_round_n729 ), .A2(_sha1_round_n514 ),.ZN(_sha1_round_n731 ) );
NOR2_X2 _sha1_round_U521  ( .A1(rnd_q[72]), .A2(rnd_q[104]), .ZN(_sha1_round_n729 ) );
NAND3_X2 _sha1_round_U520  ( .A1(rnd_q[72]), .A2(rnd_q[104]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n736 ) );
NAND3_X2 _sha1_round_U519  ( .A1(rnd_q[73]), .A2(rnd_q[105]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n728 ) );
NOR2_X2 _sha1_round_U518  ( .A1(_sha1_round_n714 ), .A2(_sha1_round_n3180 ),.ZN(_sha1_round_n716 ) );
NOR2_X2 _sha1_round_U517  ( .A1(rnd_q[74]), .A2(rnd_q[106]), .ZN(_sha1_round_n714 ) );
NOR2_X2 _sha1_round_U516  ( .A1(rnd_q[106]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n717 ) );
NAND3_X2 _sha1_round_U515  ( .A1(rnd_q[74]), .A2(rnd_q[106]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n721 ) );
NOR2_X2 _sha1_round_U514  ( .A1(rnd_q[75]), .A2(rnd_q[107]), .ZN(_sha1_round_n706 ) );
NAND3_X2 _sha1_round_U513  ( .A1(rnd_q[75]), .A2(rnd_q[107]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n713 ) );
MUX2_X2 _sha1_round_U512  ( .A(_sha1_round_n703 ), .B(_sha1_round_n702 ),.S(rnd_q[44]), .Z(_sha1_round_n704 ) );
NOR3_X2 _sha1_round_U511  ( .A1(_sha1_round_n701 ), .A2(_sha1_round_n700 ),.A3(_sha1_round_n699 ), .ZN(_sha1_round_n702 ) );
NOR2_X2 _sha1_round_U510  ( .A1(_sha1_round_n698 ), .A2(_sha1_round_n3190 ),.ZN(_sha1_round_n700 ) );
NOR2_X2 _sha1_round_U509  ( .A1(rnd_q[76]), .A2(rnd_q[108]), .ZN(_sha1_round_n698 ) );
NAND3_X2 _sha1_round_U508  ( .A1(rnd_q[76]), .A2(rnd_q[108]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n705 ) );
MUX2_X2 _sha1_round_U507  ( .A(_sha1_round_n695 ), .B(_sha1_round_n694 ),.S(rnd_q[45]), .Z(_sha1_round_n696 ) );
NOR3_X2 _sha1_round_U506  ( .A1(_sha1_round_n693 ), .A2(_sha1_round_n692 ),.A3(_sha1_round_n691 ), .ZN(_sha1_round_n694 ) );
NOR2_X2 _sha1_round_U505  ( .A1(_sha1_round_n690 ), .A2(_sha1_round_n3160 ),.ZN(_sha1_round_n692 ) );
NOR2_X2 _sha1_round_U504  ( .A1(rnd_q[77]), .A2(rnd_q[109]), .ZN(_sha1_round_n690 ) );
NAND3_X2 _sha1_round_U503  ( .A1(rnd_q[77]), .A2(rnd_q[109]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n697 ) );
MUX2_X2 _sha1_round_U502  ( .A(_sha1_round_n687 ), .B(_sha1_round_n686 ),.S(rnd_q[46]), .Z(_sha1_round_n688 ) );
NOR3_X2 _sha1_round_U501  ( .A1(_sha1_round_n685 ), .A2(_sha1_round_n684 ),.A3(_sha1_round_n683 ), .ZN(_sha1_round_n686 ) );
NOR2_X2 _sha1_round_U500  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n368 ),.ZN(_sha1_round_n683 ) );
NOR2_X2 _sha1_round_U499  ( .A1(_sha1_round_n682 ), .A2(_sha1_round_n3160 ),.ZN(_sha1_round_n684 ) );
NOR2_X2 _sha1_round_U498  ( .A1(rnd_q[78]), .A2(rnd_q[110]), .ZN(_sha1_round_n682 ) );
NAND3_X2 _sha1_round_U497  ( .A1(rnd_q[78]), .A2(rnd_q[110]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n689 ) );
NAND2_X2 _sha1_round_U496  ( .A1(_sha1_round_n681 ), .A2(_sha1_round_n680 ),.ZN(_sha1_round_f [15]) );
MUX2_X2 _sha1_round_U495  ( .A(_sha1_round_n679 ), .B(_sha1_round_n678 ),.S(rnd_q[47]), .Z(_sha1_round_n680 ) );
NOR3_X2 _sha1_round_U494  ( .A1(_sha1_round_n677 ), .A2(_sha1_round_n676 ),.A3(_sha1_round_n675 ), .ZN(_sha1_round_n678 ) );
NOR2_X2 _sha1_round_U493  ( .A1(_sha1_round_n674 ), .A2(_sha1_round_n3120 ),.ZN(_sha1_round_n676 ) );
NOR2_X2 _sha1_round_U492  ( .A1(rnd_q[79]), .A2(rnd_q[111]), .ZN(_sha1_round_n674 ) );
NAND3_X2 _sha1_round_U491  ( .A1(rnd_q[79]), .A2(rnd_q[111]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n681 ) );
NAND2_X2 _sha1_round_U490  ( .A1(_sha1_round_n673 ), .A2(_sha1_round_n672 ),.ZN(_sha1_round_f [16]) );
MUX2_X2 _sha1_round_U489  ( .A(_sha1_round_n671 ), .B(_sha1_round_n670 ),.S(rnd_q[48]), .Z(_sha1_round_n672 ) );
NOR3_X2 _sha1_round_U488  ( .A1(_sha1_round_n669 ), .A2(_sha1_round_n668 ),.A3(_sha1_round_n667 ), .ZN(_sha1_round_n670 ) );
NOR2_X2 _sha1_round_U487  ( .A1(_sha1_round_n666 ), .A2(_sha1_round_n3160 ),.ZN(_sha1_round_n668 ) );
NOR2_X2 _sha1_round_U486  ( .A1(rnd_q[80]), .A2(rnd_q[112]), .ZN(_sha1_round_n666 ) );
NAND3_X2 _sha1_round_U485  ( .A1(rnd_q[80]), .A2(rnd_q[112]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n673 ) );
NAND2_X2 _sha1_round_U484  ( .A1(_sha1_round_n665 ), .A2(_sha1_round_n664 ),.ZN(_sha1_round_f [17]) );
MUX2_X2 _sha1_round_U483  ( .A(_sha1_round_n663 ), .B(_sha1_round_n662 ),.S(rnd_q[49]), .Z(_sha1_round_n664 ) );
NOR3_X2 _sha1_round_U482  ( .A1(_sha1_round_n661 ), .A2(_sha1_round_n660 ),.A3(_sha1_round_n659 ), .ZN(_sha1_round_n662 ) );
NOR2_X2 _sha1_round_U481  ( .A1(_sha1_round_n658 ), .A2(_sha1_round_n3200 ),.ZN(_sha1_round_n660 ) );
NOR2_X2 _sha1_round_U480  ( .A1(rnd_q[81]), .A2(rnd_q[113]), .ZN(_sha1_round_n658 ) );
NAND3_X2 _sha1_round_U479  ( .A1(rnd_q[81]), .A2(rnd_q[113]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n665 ) );
NAND2_X2 _sha1_round_U478  ( .A1(_sha1_round_n657 ), .A2(_sha1_round_n656 ),.ZN(_sha1_round_f [18]) );
MUX2_X2 _sha1_round_U477  ( .A(_sha1_round_n655 ), .B(_sha1_round_n654 ),.S(rnd_q[50]), .Z(_sha1_round_n656 ) );
NOR3_X2 _sha1_round_U476  ( .A1(_sha1_round_n653 ), .A2(_sha1_round_n652 ),.A3(_sha1_round_n651 ), .ZN(_sha1_round_n654 ) );
NOR2_X2 _sha1_round_U475  ( .A1(_sha1_round_n650 ), .A2(_sha1_round_n513 ),.ZN(_sha1_round_n652 ) );
NOR2_X2 _sha1_round_U474  ( .A1(rnd_q[82]), .A2(rnd_q[114]), .ZN(_sha1_round_n650 ) );
NAND3_X2 _sha1_round_U473  ( .A1(rnd_q[82]), .A2(rnd_q[114]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n657 ) );
NAND2_X2 _sha1_round_U472  ( .A1(_sha1_round_n649 ), .A2(_sha1_round_n648 ),.ZN(_sha1_round_f [19]) );
MUX2_X2 _sha1_round_U471  ( .A(_sha1_round_n647 ), .B(_sha1_round_n646 ),.S(rnd_q[51]), .Z(_sha1_round_n648 ) );
NOR3_X2 _sha1_round_U470  ( .A1(_sha1_round_n645 ), .A2(_sha1_round_n644 ),.A3(_sha1_round_n643 ), .ZN(_sha1_round_n646 ) );
NOR2_X2 _sha1_round_U469  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n371 ),.ZN(_sha1_round_n643 ) );
NOR2_X2 _sha1_round_U468  ( .A1(_sha1_round_n642 ), .A2(_sha1_round_n3180 ),.ZN(_sha1_round_n644 ) );
NOR2_X2 _sha1_round_U467  ( .A1(rnd_q[83]), .A2(rnd_q[115]), .ZN(_sha1_round_n642 ) );
NAND3_X2 _sha1_round_U466  ( .A1(rnd_q[83]), .A2(rnd_q[115]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n649 ) );
MUX2_X2 _sha1_round_U465  ( .A(_sha1_round_n639 ), .B(_sha1_round_n638 ),.S(rnd_q[52]), .Z(_sha1_round_n640 ) );
NOR3_X2 _sha1_round_U464  ( .A1(_sha1_round_n637 ), .A2(_sha1_round_n636 ),.A3(_sha1_round_n635 ), .ZN(_sha1_round_n638 ) );
NOR2_X2 _sha1_round_U463  ( .A1(_sha1_round_n634 ), .A2(_sha1_round_n3180 ),.ZN(_sha1_round_n636 ) );
NOR2_X2 _sha1_round_U462  ( .A1(rnd_q[84]), .A2(rnd_q[116]), .ZN(_sha1_round_n634 ) );
NAND3_X2 _sha1_round_U461  ( .A1(rnd_q[84]), .A2(rnd_q[116]), .A3(_sha1_round_n517 ), .ZN(_sha1_round_n641 ) );
NAND2_X2 _sha1_round_U460  ( .A1(_sha1_round_n633 ), .A2(_sha1_round_n632 ),.ZN(_sha1_round_f [21]) );
MUX2_X2 _sha1_round_U459  ( .A(_sha1_round_n631 ), .B(_sha1_round_n630 ),.S(rnd_q[53]), .Z(_sha1_round_n632 ) );
NOR3_X2 _sha1_round_U458  ( .A1(_sha1_round_n629 ), .A2(_sha1_round_n628 ),.A3(_sha1_round_n627 ), .ZN(_sha1_round_n630 ) );
NOR2_X2 _sha1_round_U457  ( .A1(_sha1_round_n626 ), .A2(_sha1_round_n514 ),.ZN(_sha1_round_n628 ) );
NOR2_X2 _sha1_round_U456  ( .A1(rnd_q[85]), .A2(rnd_q[117]), .ZN(_sha1_round_n626 ) );
NAND3_X2 _sha1_round_U455  ( .A1(rnd_q[85]), .A2(rnd_q[117]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n633 ) );
NAND2_X2 _sha1_round_U454  ( .A1(_sha1_round_n625 ), .A2(_sha1_round_n624 ),.ZN(_sha1_round_f [22]) );
MUX2_X2 _sha1_round_U453  ( .A(_sha1_round_n623 ), .B(_sha1_round_n622 ),.S(rnd_q[54]), .Z(_sha1_round_n624 ) );
NOR3_X2 _sha1_round_U452  ( .A1(_sha1_round_n621 ), .A2(_sha1_round_n620 ),.A3(_sha1_round_n619 ), .ZN(_sha1_round_n622 ) );
NOR2_X2 _sha1_round_U451  ( .A1(_sha1_round_n618 ), .A2(_sha1_round_n514 ),.ZN(_sha1_round_n620 ) );
NOR2_X2 _sha1_round_U450  ( .A1(rnd_q[86]), .A2(rnd_q[118]), .ZN(_sha1_round_n618 ) );
NAND3_X2 _sha1_round_U449  ( .A1(rnd_q[86]), .A2(rnd_q[118]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n625 ) );
NAND2_X2 _sha1_round_U448  ( .A1(_sha1_round_n617 ), .A2(_sha1_round_n616 ),.ZN(_sha1_round_f [23]) );
MUX2_X2 _sha1_round_U447  ( .A(_sha1_round_n615 ), .B(_sha1_round_n614 ),.S(rnd_q[55]), .Z(_sha1_round_n616 ) );
AND3_X2 _sha1_round_U446  ( .A1(_sha1_round_n613 ), .A2(_sha1_round_n612 ),.A3(_sha1_round_n611 ), .ZN(_sha1_round_n614 ) );
NAND2_X2 _sha1_round_U445  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n610 ),.ZN(_sha1_round_n611 ) );
INV_X4 _sha1_round_U444  ( .A(rnd_q[119]), .ZN(_sha1_round_n610 ) );
NAND2_X2 _sha1_round_U443  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n609 ),.ZN(_sha1_round_n615 ) );
INV_X4 _sha1_round_U442  ( .A(_sha1_round_n168 ), .ZN(_sha1_round_n609 ) );
NAND3_X2 _sha1_round_U441  ( .A1(rnd_q[87]), .A2(rnd_q[119]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n617 ) );
NAND2_X2 _sha1_round_U440  ( .A1(_sha1_round_n608 ), .A2(_sha1_round_n607 ),.ZN(_sha1_round_f [24]) );
MUX2_X2 _sha1_round_U439  ( .A(_sha1_round_n606 ), .B(_sha1_round_n605 ),.S(rnd_q[56]), .Z(_sha1_round_n607 ) );
AND3_X2 _sha1_round_U438  ( .A1(_sha1_round_n604 ), .A2(_sha1_round_n603 ),.A3(_sha1_round_n602 ), .ZN(_sha1_round_n605 ) );
NAND2_X2 _sha1_round_U437  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n601 ),.ZN(_sha1_round_n602 ) );
INV_X4 _sha1_round_U436  ( .A(rnd_q[120]), .ZN(_sha1_round_n601 ) );
NAND2_X2 _sha1_round_U435  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n600 ),.ZN(_sha1_round_n606 ) );
INV_X4 _sha1_round_U434  ( .A(_sha1_round_n159 ), .ZN(_sha1_round_n600 ) );
NAND3_X2 _sha1_round_U433  ( .A1(rnd_q[88]), .A2(rnd_q[120]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n608 ) );
NAND2_X2 _sha1_round_U432  ( .A1(_sha1_round_n599 ), .A2(_sha1_round_n598 ),.ZN(_sha1_round_f [25]) );
MUX2_X2 _sha1_round_U431  ( .A(_sha1_round_n597 ), .B(_sha1_round_n596 ),.S(rnd_q[57]), .Z(_sha1_round_n598 ) );
AND3_X2 _sha1_round_U430  ( .A1(_sha1_round_n595 ), .A2(_sha1_round_n594 ),.A3(_sha1_round_n593 ), .ZN(_sha1_round_n596 ) );
NAND2_X2 _sha1_round_U429  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n592 ),.ZN(_sha1_round_n593 ) );
INV_X4 _sha1_round_U428  ( .A(rnd_q[121]), .ZN(_sha1_round_n592 ) );
NAND2_X2 _sha1_round_U427  ( .A1(_sha1_round_n150 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n594 ) );
NAND2_X2 _sha1_round_U426  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n591 ),.ZN(_sha1_round_n597 ) );
INV_X4 _sha1_round_U425  ( .A(_sha1_round_n150 ), .ZN(_sha1_round_n591 ) );
NAND3_X2 _sha1_round_U424  ( .A1(rnd_q[89]), .A2(rnd_q[121]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n599 ) );
NAND2_X2 _sha1_round_U423  ( .A1(_sha1_round_n590 ), .A2(_sha1_round_n589 ),.ZN(_sha1_round_f [26]) );
MUX2_X2 _sha1_round_U422  ( .A(_sha1_round_n588 ), .B(_sha1_round_n587 ),.S(rnd_q[58]), .Z(_sha1_round_n589 ) );
AND3_X2 _sha1_round_U421  ( .A1(_sha1_round_n586 ), .A2(_sha1_round_n585 ),.A3(_sha1_round_n584 ), .ZN(_sha1_round_n587 ) );
NAND2_X2 _sha1_round_U420  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n583 ),.ZN(_sha1_round_n584 ) );
INV_X4 _sha1_round_U419  ( .A(rnd_q[122]), .ZN(_sha1_round_n583 ) );
NAND2_X2 _sha1_round_U418  ( .A1(_sha1_round_n141 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n585 ) );
NAND2_X2 _sha1_round_U417  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n582 ),.ZN(_sha1_round_n588 ) );
INV_X4 _sha1_round_U416  ( .A(_sha1_round_n141 ), .ZN(_sha1_round_n582 ) );
NAND3_X2 _sha1_round_U415  ( .A1(rnd_q[90]), .A2(rnd_q[122]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n590 ) );
NAND2_X2 _sha1_round_U414  ( .A1(_sha1_round_n581 ), .A2(_sha1_round_n580 ),.ZN(_sha1_round_f [27]) );
MUX2_X2 _sha1_round_U413  ( .A(_sha1_round_n579 ), .B(_sha1_round_n578 ),.S(rnd_q[59]), .Z(_sha1_round_n580 ) );
AND3_X2 _sha1_round_U412  ( .A1(_sha1_round_n577 ), .A2(_sha1_round_n576 ),.A3(_sha1_round_n575 ), .ZN(_sha1_round_n578 ) );
NAND2_X2 _sha1_round_U411  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n574 ),.ZN(_sha1_round_n575 ) );
INV_X4 _sha1_round_U410  ( .A(rnd_q[123]), .ZN(_sha1_round_n574 ) );
NAND2_X2 _sha1_round_U409  ( .A1(_sha1_round_n132 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n576 ) );
NAND2_X2 _sha1_round_U408  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n573 ),.ZN(_sha1_round_n579 ) );
INV_X4 _sha1_round_U407  ( .A(_sha1_round_n132 ), .ZN(_sha1_round_n573 ) );
NAND3_X2 _sha1_round_U406  ( .A1(rnd_q[91]), .A2(rnd_q[123]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n581 ) );
NAND2_X2 _sha1_round_U405  ( .A1(_sha1_round_n572 ), .A2(_sha1_round_n571 ),.ZN(_sha1_round_f [28]) );
MUX2_X2 _sha1_round_U404  ( .A(_sha1_round_n570 ), .B(_sha1_round_n569 ),.S(rnd_q[60]), .Z(_sha1_round_n571 ) );
AND3_X2 _sha1_round_U403  ( .A1(_sha1_round_n568 ), .A2(_sha1_round_n567 ),.A3(_sha1_round_n566 ), .ZN(_sha1_round_n569 ) );
NAND2_X2 _sha1_round_U402  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n565 ),.ZN(_sha1_round_n566 ) );
INV_X4 _sha1_round_U401  ( .A(rnd_q[124]), .ZN(_sha1_round_n565 ) );
NAND2_X2 _sha1_round_U400  ( .A1(_sha1_round_n123 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n567 ) );
NAND2_X2 _sha1_round_U399  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n564 ),.ZN(_sha1_round_n570 ) );
INV_X4 _sha1_round_U398  ( .A(_sha1_round_n123 ), .ZN(_sha1_round_n564 ) );
NAND3_X2 _sha1_round_U397  ( .A1(rnd_q[92]), .A2(rnd_q[124]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n572 ) );
NAND2_X2 _sha1_round_U396  ( .A1(_sha1_round_n563 ), .A2(_sha1_round_n562 ),.ZN(_sha1_round_f [29]) );
MUX2_X2 _sha1_round_U395  ( .A(_sha1_round_n561 ), .B(_sha1_round_n560 ),.S(rnd_q[61]), .Z(_sha1_round_n562 ) );
AND3_X2 _sha1_round_U394  ( .A1(_sha1_round_n559 ), .A2(_sha1_round_n558 ),.A3(_sha1_round_n557 ), .ZN(_sha1_round_n560 ) );
NAND2_X2 _sha1_round_U393  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n556 ),.ZN(_sha1_round_n557 ) );
INV_X4 _sha1_round_U392  ( .A(rnd_q[125]), .ZN(_sha1_round_n556 ) );
NAND2_X2 _sha1_round_U391  ( .A1(_sha1_round_n114 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n558 ) );
NAND2_X2 _sha1_round_U390  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n555 ),.ZN(_sha1_round_n561 ) );
INV_X4 _sha1_round_U389  ( .A(_sha1_round_n114 ), .ZN(_sha1_round_n555 ) );
NAND3_X2 _sha1_round_U388  ( .A1(rnd_q[93]), .A2(rnd_q[125]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n563 ) );
NAND2_X2 _sha1_round_U387  ( .A1(_sha1_round_n554 ), .A2(_sha1_round_n553 ),.ZN(_sha1_round_f [30]) );
MUX2_X2 _sha1_round_U386  ( .A(_sha1_round_n552 ), .B(_sha1_round_n551 ),.S(rnd_q[62]), .Z(_sha1_round_n553 ) );
AND3_X2 _sha1_round_U385  ( .A1(_sha1_round_n550 ), .A2(_sha1_round_n549 ),.A3(_sha1_round_n548 ), .ZN(_sha1_round_n551 ) );
NAND2_X2 _sha1_round_U384  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n547 ),.ZN(_sha1_round_n548 ) );
INV_X4 _sha1_round_U383  ( .A(rnd_q[126]), .ZN(_sha1_round_n547 ) );
NAND2_X2 _sha1_round_U382  ( .A1(_sha1_round_n96 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n549 ) );
NAND2_X2 _sha1_round_U381  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n546 ),.ZN(_sha1_round_n552 ) );
INV_X4 _sha1_round_U380  ( .A(_sha1_round_n96 ), .ZN(_sha1_round_n546 ) );
NAND3_X2 _sha1_round_U379  ( .A1(rnd_q[94]), .A2(rnd_q[126]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n554 ) );
NAND2_X2 _sha1_round_U378  ( .A1(_sha1_round_n545 ), .A2(_sha1_round_n544 ),.ZN(_sha1_round_f [31]) );
MUX2_X2 _sha1_round_U377  ( .A(_sha1_round_n543 ), .B(_sha1_round_n542 ),.S(rnd_q[63]), .Z(_sha1_round_n544 ) );
AND3_X2 _sha1_round_U376  ( .A1(_sha1_round_n541 ), .A2(_sha1_round_n540 ),.A3(_sha1_round_n539 ), .ZN(_sha1_round_n542 ) );
NAND2_X2 _sha1_round_U375  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_n538 ),.ZN(_sha1_round_n539 ) );
INV_X4 _sha1_round_U374  ( .A(rnd_q[127]), .ZN(_sha1_round_n538 ) );
NAND2_X2 _sha1_round_U373  ( .A1(_sha1_round_n87 ), .A2(_sha1_round_n3370 ),.ZN(_sha1_round_n540 ) );
NAND2_X2 _sha1_round_U372  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_n537 ),.ZN(_sha1_round_n543 ) );
INV_X4 _sha1_round_U371  ( .A(_sha1_round_n87 ), .ZN(_sha1_round_n537 ) );
NAND3_X2 _sha1_round_U370  ( .A1(rnd_q[95]), .A2(rnd_q[127]), .A3(_sha1_round_n3300 ), .ZN(_sha1_round_n545 ) );
NAND2_X2 _sha1_round_U369  ( .A1(_sha1_round_n533 ), .A2(_sha1_round_n534 ),.ZN(_sha1_round_n536 ) );
INV_X4 _sha1_round_U368  ( .A(_sha1_round_n520 ), .ZN(_sha1_round_n532 ) );
INV_X32 _sha1_round_U367  ( .A(_sha1_round_n516 ), .ZN(_sha1_round_n515 ) );
NAND2_X4 _sha1_round_U366  ( .A1(_sha1_round_n510 ), .A2(_sha1_round_n3120 ),.ZN(_sha1_round_k[3] ) );
NAND2_X4 _sha1_round_U365  ( .A1(_sha1_round_n530 ), .A2(_sha1_round_n529 ),.ZN(_sha1_round_n819 ) );
NAND2_X4 _sha1_round_U364  ( .A1(_sha1_round_n819 ), .A2(_sha1_round_n820 ),.ZN(_sha1_round_n823 ) );
NAND2_X4 _sha1_round_U363  ( .A1(_sha1_round_n748 ), .A2(_sha1_round_n749 ),.ZN(_sha1_round_f [6]) );
NAND2_X1 _sha1_round_U362  ( .A1(rnd_cnt_q[6]), .A2(_sha1_round_n531 ), .ZN(_sha1_round_n534 ) );
NAND2_X4 _sha1_round_U361  ( .A1(_sha1_round_n536 ), .A2(_sha1_round_n535 ),.ZN(_sha1_round_n820 ) );
NAND3_X1 _sha1_round_U360  ( .A1(rnd_q[35]), .A2(_sha1_round_n767 ), .A3(_sha1_round_n766 ), .ZN(_sha1_round_n775 ) );
INV_X16 _sha1_round_U359  ( .A(_sha1_round_n823 ), .ZN(_sha1_round_n516 ) );
NAND2_X1 _sha1_round_U358  ( .A1(_sha1_round_n819 ), .A2(_sha1_round_n514 ),.ZN(_sha1_round_k_26 ) );
NAND2_X2 _sha1_round_U357  ( .A1(_sha1_round_n818 ), .A2(_sha1_round_n819 ),.ZN(_sha1_round_k_27 ) );
NAND2_X4 _sha1_round_U356  ( .A1(_sha1_round_n727 ), .A2(_sha1_round_n728 ),.ZN(_sha1_round_f [9]) );
INV_X1 _sha1_round_U355  ( .A(_sha1_round_n820 ), .ZN(_sha1_round_n824 ) );
INV_X4 _sha1_round_U354  ( .A(_sha1_round_N332 ), .ZN(_sha1_round_n508 ) );
NOR2_X1 _sha1_round_U353  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n378 ),.ZN(_sha1_round_n699 ) );
NOR2_X1 _sha1_round_U352  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n376 ),.ZN(_sha1_round_n659 ) );
NOR2_X1 _sha1_round_U351  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n380 ),.ZN(_sha1_round_n619 ) );
NAND2_X1 _sha1_round_U350  ( .A1(_sha1_round_n510 ), .A2(_sha1_round_n516 ),.ZN(_sha1_round_k_30 ) );
NAND2_X1 _sha1_round_U349  ( .A1(_sha1_round_n363 ), .A2(_sha1_round_n516 ),.ZN(_sha1_round_k[15] ) );
NAND3_X1 _sha1_round_U348  ( .A1(_sha1_round_n765 ), .A2(_sha1_round_n764 ),.A3(_sha1_round_n767 ), .ZN(_sha1_round_n777 ) );
NAND2_X1 _sha1_round_U347  ( .A1(_sha1_round_n3150 ), .A2(_sha1_round_n783 ),.ZN(_sha1_round_n784 ) );
NAND2_X1 _sha1_round_U346  ( .A1(_sha1_round_n3150 ), .A2(_sha1_round_n809 ),.ZN(_sha1_round_n810 ) );
NAND2_X1 _sha1_round_U345  ( .A1(_sha1_round_n167 ), .A2(_sha1_round_n360 ),.ZN(_sha1_round_n613 ) );
NAND2_X1 _sha1_round_U344  ( .A1(_sha1_round_n149 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n595 ) );
NAND2_X1 _sha1_round_U343  ( .A1(_sha1_round_n158 ), .A2(_sha1_round_n360 ),.ZN(_sha1_round_n604 ) );
NAND2_X1 _sha1_round_U342  ( .A1(_sha1_round_n140 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n586 ) );
NAND2_X1 _sha1_round_U341  ( .A1(_sha1_round_n131 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n577 ) );
NAND2_X1 _sha1_round_U340  ( .A1(_sha1_round_n122 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n568 ) );
NAND2_X1 _sha1_round_U339  ( .A1(_sha1_round_n113 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n559 ) );
NAND2_X1 _sha1_round_U338  ( .A1(_sha1_round_n95 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n550 ) );
NAND2_X1 _sha1_round_U337  ( .A1(_sha1_round_n86 ), .A2(_sha1_round_n364 ),.ZN(_sha1_round_n541 ) );
BUF_X4 _sha1_round_U336  ( .A(rnd_q[137]), .Z(sha1_round_wire[105]) );
BUF_X4 _sha1_round_U335  ( .A(rnd_q[138]), .Z(sha1_round_wire[106]) );
BUF_X4 _sha1_round_U334  ( .A(rnd_q[139]), .Z(sha1_round_wire[107]) );
BUF_X4 _sha1_round_U333  ( .A(rnd_q[140]), .Z(sha1_round_wire[108]) );
BUF_X4 _sha1_round_U332  ( .A(rnd_q[141]), .Z(sha1_round_wire[109]) );
BUF_X4 _sha1_round_U331  ( .A(rnd_q[142]), .Z(sha1_round_wire[110]) );
BUF_X4 _sha1_round_U330  ( .A(rnd_q[143]), .Z(sha1_round_wire[111]) );
BUF_X4 _sha1_round_U329  ( .A(rnd_q[144]), .Z(sha1_round_wire[112]) );
BUF_X4 _sha1_round_U328  ( .A(rnd_q[145]), .Z(sha1_round_wire[113]) );
BUF_X4 _sha1_round_U327  ( .A(rnd_q[146]), .Z(sha1_round_wire[114]) );
BUF_X4 _sha1_round_U326  ( .A(rnd_q[147]), .Z(sha1_round_wire[115]) );
BUF_X4 _sha1_round_U325  ( .A(rnd_q[148]), .Z(sha1_round_wire[116]) );
BUF_X4 _sha1_round_U324  ( .A(rnd_q[149]), .Z(sha1_round_wire[117]) );
BUF_X4 _sha1_round_U323  ( .A(rnd_q[150]), .Z(sha1_round_wire[118]) );
BUF_X4 _sha1_round_U322  ( .A(rnd_q[151]), .Z(sha1_round_wire[119]) );
BUF_X4 _sha1_round_U321  ( .A(rnd_q[152]), .Z(sha1_round_wire[120]) );
BUF_X4 _sha1_round_U320  ( .A(rnd_q[153]), .Z(sha1_round_wire[121]) );
BUF_X4 _sha1_round_U319  ( .A(rnd_q[154]), .Z(sha1_round_wire[122]) );
BUF_X4 _sha1_round_U318  ( .A(rnd_q[155]), .Z(sha1_round_wire[123]) );
BUF_X4 _sha1_round_U317  ( .A(rnd_q[156]), .Z(sha1_round_wire[124]) );
BUF_X4 _sha1_round_U316  ( .A(rnd_q[157]), .Z(sha1_round_wire[125]) );
BUF_X4 _sha1_round_U315  ( .A(rnd_q[158]), .Z(sha1_round_wire[126]) );
BUF_X4 _sha1_round_U314  ( .A(rnd_q[159]), .Z(sha1_round_wire[127]) );
INV_X4 _sha1_round_U313  ( .A(rnd_cnt_q[3]), .ZN(_sha1_round_n524 ) );
BUF_X4 _sha1_round_U312  ( .A(rnd_q[134]), .Z(sha1_round_wire[102]) );
BUF_X4 _sha1_round_U311  ( .A(rnd_q[133]), .Z(sha1_round_wire[101]) );
BUF_X4 _sha1_round_U310  ( .A(rnd_q[131]), .Z(sha1_round_wire[99]) );
BUF_X4 _sha1_round_U309  ( .A(rnd_q[130]), .Z(sha1_round_wire[98]) );
BUF_X4 _sha1_round_U308  ( .A(rnd_q[129]), .Z(sha1_round_wire[97]) );
BUF_X4 _sha1_round_U307  ( .A(rnd_q[128]), .Z(sha1_round_wire[96]) );
BUF_X4 _sha1_round_U306  ( .A(rnd_q[96]), .Z(sha1_round_wire[94]) );
BUF_X4 _sha1_round_U305  ( .A(rnd_q[117]), .Z(sha1_round_wire[83]) );
BUF_X4 _sha1_round_U304  ( .A(rnd_q[116]), .Z(sha1_round_wire[82]) );
BUF_X4 _sha1_round_U303  ( .A(rnd_q[113]), .Z(sha1_round_wire[79]) );
BUF_X4 _sha1_round_U302  ( .A(rnd_q[112]), .Z(sha1_round_wire[78]) );
BUF_X4 _sha1_round_U301  ( .A(rnd_q[110]), .Z(sha1_round_wire[76]) );
BUF_X4 _sha1_round_U300  ( .A(rnd_q[109]), .Z(sha1_round_wire[75]) );
BUF_X4 _sha1_round_U299  ( .A(rnd_q[106]), .Z(sha1_round_wire[72]) );
BUF_X4 _sha1_round_U298  ( .A(rnd_q[105]), .Z(sha1_round_wire[71]) );
BUF_X4 _sha1_round_U297  ( .A(rnd_q[104]), .Z(sha1_round_wire[70]) );
BUF_X4 _sha1_round_U296  ( .A(rnd_q[103]), .Z(sha1_round_wire[69]) );
BUF_X4 _sha1_round_U295  ( .A(rnd_q[99]), .Z(sha1_round_wire[65]) );
BUF_X4 _sha1_round_U294  ( .A(rnd_q[95]), .Z(sha1_round_wire[63]) );
BUF_X4 _sha1_round_U293  ( .A(rnd_q[91]), .Z(sha1_round_wire[59]) );
BUF_X4 _sha1_round_U292  ( .A(rnd_q[90]), .Z(sha1_round_wire[58]) );
BUF_X4 _sha1_round_U291  ( .A(rnd_q[89]), .Z(sha1_round_wire[57]) );
BUF_X4 _sha1_round_U290  ( .A(rnd_q[88]), .Z(sha1_round_wire[56]) );
BUF_X4 _sha1_round_U289  ( .A(rnd_q[87]), .Z(sha1_round_wire[55]) );
BUF_X4 _sha1_round_U288  ( .A(rnd_q[85]), .Z(sha1_round_wire[53]) );
BUF_X4 _sha1_round_U287  ( .A(rnd_q[81]), .Z(sha1_round_wire[49]) );
BUF_X4 _sha1_round_U286  ( .A(rnd_q[80]), .Z(sha1_round_wire[48]) );
BUF_X4 _sha1_round_U285  ( .A(rnd_q[78]), .Z(sha1_round_wire[46]) );
BUF_X4 _sha1_round_U284  ( .A(rnd_q[76]), .Z(sha1_round_wire[44]) );
BUF_X4 _sha1_round_U283  ( .A(rnd_q[74]), .Z(sha1_round_wire[42]) );
BUF_X4 _sha1_round_U282  ( .A(rnd_q[72]), .Z(sha1_round_wire[40]) );
BUF_X4 _sha1_round_U281  ( .A(rnd_q[71]), .Z(sha1_round_wire[39]) );
BUF_X4 _sha1_round_U280  ( .A(rnd_q[67]), .Z(sha1_round_wire[35]) );
BUF_X4 _sha1_round_U279  ( .A(rnd_q[66]), .Z(sha1_round_wire[34]) );
BUF_X4 _sha1_round_U278  ( .A(rnd_q[65]), .Z(sha1_round_wire[33]) );
BUF_X4 _sha1_round_U277  ( .A(rnd_q[62]), .Z(sha1_round_wire[30]) );
BUF_X4 _sha1_round_U276  ( .A(rnd_q[61]), .Z(sha1_round_wire[29]) );
BUF_X4 _sha1_round_U275  ( .A(rnd_q[60]), .Z(sha1_round_wire[28]) );
BUF_X4 _sha1_round_U274  ( .A(rnd_q[59]), .Z(sha1_round_wire[27]) );
BUF_X4 _sha1_round_U273  ( .A(rnd_q[58]), .Z(sha1_round_wire[26]) );
BUF_X4 _sha1_round_U272  ( .A(rnd_q[57]), .Z(sha1_round_wire[25]) );
BUF_X4 _sha1_round_U271  ( .A(rnd_q[55]), .Z(sha1_round_wire[23]) );
BUF_X4 _sha1_round_U270  ( .A(rnd_q[54]), .Z(sha1_round_wire[22]) );
BUF_X4 _sha1_round_U269  ( .A(rnd_q[53]), .Z(sha1_round_wire[21]) );
BUF_X4 _sha1_round_U268  ( .A(rnd_q[51]), .Z(sha1_round_wire[19]) );
BUF_X4 _sha1_round_U267  ( .A(rnd_q[50]), .Z(sha1_round_wire[18]) );
BUF_X4 _sha1_round_U266  ( .A(rnd_q[49]), .Z(sha1_round_wire[17]) );
BUF_X4 _sha1_round_U265  ( .A(rnd_q[47]), .Z(sha1_round_wire[15]) );
BUF_X4 _sha1_round_U264  ( .A(rnd_q[46]), .Z(sha1_round_wire[14]) );
BUF_X4 _sha1_round_U263  ( .A(rnd_q[43]), .Z(sha1_round_wire[11]) );
BUF_X4 _sha1_round_U262  ( .A(rnd_q[42]), .Z(sha1_round_wire[10]) );
BUF_X4 _sha1_round_U261  ( .A(rnd_q[41]), .Z(sha1_round_wire[9]) );
BUF_X4 _sha1_round_U260  ( .A(rnd_q[38]), .Z(sha1_round_wire[6]) );
BUF_X4 _sha1_round_U259  ( .A(rnd_q[37]), .Z(sha1_round_wire[5]) );
BUF_X4 _sha1_round_U258  ( .A(rnd_q[36]), .Z(sha1_round_wire[4]) );
BUF_X4 _sha1_round_U257  ( .A(rnd_q[35]), .Z(sha1_round_wire[3]) );
BUF_X4 _sha1_round_U256  ( .A(rnd_q[34]), .Z(sha1_round_wire[2]) );
BUF_X4 _sha1_round_U255  ( .A(rnd_q[33]), .Z(sha1_round_wire[1]) );
BUF_X4 _sha1_round_U254  ( .A(rnd_q[32]), .Z(sha1_round_wire[0]) );
BUF_X4 _sha1_round_U253  ( .A(rnd_q[136]), .Z(sha1_round_wire[104]) );
BUF_X4 _sha1_round_U252  ( .A(rnd_q[135]), .Z(sha1_round_wire[103]) );
BUF_X4 _sha1_round_U251  ( .A(rnd_q[132]), .Z(sha1_round_wire[100]) );
BUF_X4 _sha1_round_U250  ( .A(rnd_q[127]), .Z(sha1_round_wire[93]) );
BUF_X4 _sha1_round_U249  ( .A(rnd_q[126]), .Z(sha1_round_wire[92]) );
BUF_X4 _sha1_round_U248  ( .A(rnd_q[125]), .Z(sha1_round_wire[91]) );
BUF_X4 _sha1_round_U247  ( .A(rnd_q[124]), .Z(sha1_round_wire[90]) );
BUF_X4 _sha1_round_U246  ( .A(rnd_q[123]), .Z(sha1_round_wire[89]) );
BUF_X4 _sha1_round_U245  ( .A(rnd_q[122]), .Z(sha1_round_wire[88]) );
BUF_X4 _sha1_round_U244  ( .A(rnd_q[121]), .Z(sha1_round_wire[87]) );
BUF_X4 _sha1_round_U243  ( .A(rnd_q[119]), .Z(sha1_round_wire[85]) );
BUF_X4 _sha1_round_U242  ( .A(rnd_q[118]), .Z(sha1_round_wire[84]) );
BUF_X4 _sha1_round_U241  ( .A(rnd_q[115]), .Z(sha1_round_wire[81]) );
BUF_X4 _sha1_round_U240  ( .A(rnd_q[114]), .Z(sha1_round_wire[80]) );
BUF_X4 _sha1_round_U239  ( .A(rnd_q[111]), .Z(sha1_round_wire[77]) );
BUF_X4 _sha1_round_U238  ( .A(rnd_q[107]), .Z(sha1_round_wire[73]) );
BUF_X4 _sha1_round_U237  ( .A(rnd_q[100]), .Z(sha1_round_wire[66]) );
BUF_X4 _sha1_round_U236  ( .A(rnd_q[94]), .Z(sha1_round_wire[62]) );
BUF_X4 _sha1_round_U235  ( .A(rnd_q[93]), .Z(sha1_round_wire[61]) );
BUF_X4 _sha1_round_U234  ( .A(rnd_q[92]), .Z(sha1_round_wire[60]) );
BUF_X4 _sha1_round_U233  ( .A(rnd_q[86]), .Z(sha1_round_wire[54]) );
BUF_X4 _sha1_round_U232  ( .A(rnd_q[83]), .Z(sha1_round_wire[51]) );
BUF_X4 _sha1_round_U231  ( .A(rnd_q[82]), .Z(sha1_round_wire[50]) );
BUF_X4 _sha1_round_U230  ( .A(rnd_q[79]), .Z(sha1_round_wire[47]) );
BUF_X4 _sha1_round_U229  ( .A(rnd_q[75]), .Z(sha1_round_wire[43]) );
BUF_X4 _sha1_round_U228  ( .A(rnd_q[68]), .Z(sha1_round_wire[36]) );
BUF_X4 _sha1_round_U227  ( .A(rnd_q[64]), .Z(sha1_round_wire[32]) );
BUF_X4 _sha1_round_U226  ( .A(rnd_q[63]), .Z(sha1_round_wire[31]) );
BUF_X4 _sha1_round_U225  ( .A(rnd_q[56]), .Z(sha1_round_wire[24]) );
BUF_X4 _sha1_round_U224  ( .A(rnd_q[48]), .Z(sha1_round_wire[16]) );
BUF_X4 _sha1_round_U223  ( .A(rnd_q[45]), .Z(sha1_round_wire[13]) );
BUF_X4 _sha1_round_U222  ( .A(rnd_q[44]), .Z(sha1_round_wire[12]) );
BUF_X4 _sha1_round_U221  ( .A(rnd_q[40]), .Z(sha1_round_wire[8]) );
BUF_X4 _sha1_round_U220  ( .A(rnd_q[120]), .Z(sha1_round_wire[86]) );
BUF_X4 _sha1_round_U219  ( .A(rnd_q[108]), .Z(sha1_round_wire[74]) );
BUF_X4 _sha1_round_U218  ( .A(rnd_q[98]), .Z(sha1_round_wire[64]) );
BUF_X4 _sha1_round_U217  ( .A(rnd_q[52]), .Z(sha1_round_wire[20]) );
BUF_X4 _sha1_round_U216  ( .A(rnd_q[97]), .Z(sha1_round_wire[95]) );
BUF_X4 _sha1_round_U215  ( .A(rnd_q[77]), .Z(sha1_round_wire[45]) );
BUF_X4 _sha1_round_U214  ( .A(rnd_q[73]), .Z(sha1_round_wire[41]) );
BUF_X4 _sha1_round_U213  ( .A(rnd_q[84]), .Z(sha1_round_wire[52]) );
BUF_X4 _sha1_round_U212  ( .A(rnd_q[70]), .Z(sha1_round_wire[38]) );
BUF_X4 _sha1_round_U211  ( .A(rnd_q[102]), .Z(sha1_round_wire[68]) );
BUF_X4 _sha1_round_U210  ( .A(rnd_q[69]), .Z(sha1_round_wire[37]) );
BUF_X4 _sha1_round_U209  ( .A(rnd_q[101]), .Z(sha1_round_wire[67]) );
XOR2_X2 _sha1_round_U208  ( .A(rnd_q[118]), .B(rnd_q[86]), .Z(_sha1_round_n380 ) );
XOR2_X2 _sha1_round_U207  ( .A(rnd_q[112]), .B(rnd_q[80]), .Z(_sha1_round_n379 ) );
XOR2_X2 _sha1_round_U206  ( .A(rnd_q[108]), .B(rnd_q[76]), .Z(_sha1_round_n378 ) );
XOR2_X2 _sha1_round_U205  ( .A(rnd_q[109]), .B(rnd_q[77]), .Z(_sha1_round_n377 ) );
XOR2_X2 _sha1_round_U204  ( .A(rnd_q[113]), .B(rnd_q[81]), .Z(_sha1_round_n376 ) );
XOR2_X2 _sha1_round_U203  ( .A(rnd_q[111]), .B(rnd_q[79]), .Z(_sha1_round_n375 ) );
XOR2_X2 _sha1_round_U202  ( .A(rnd_q[100]), .B(rnd_q[68]), .Z(_sha1_round_n374 ) );
XOR2_X2 _sha1_round_U201  ( .A(rnd_q[114]), .B(rnd_q[82]), .Z(_sha1_round_n373 ) );
XOR2_X2 _sha1_round_U200  ( .A(rnd_q[107]), .B(rnd_q[75]), .Z(_sha1_round_n372 ) );
XOR2_X2 _sha1_round_U199  ( .A(rnd_q[115]), .B(rnd_q[83]), .Z(_sha1_round_n371 ) );
XOR2_X2 _sha1_round_U198  ( .A(rnd_q[104]), .B(rnd_q[72]), .Z(_sha1_round_n370 ) );
XOR2_X2 _sha1_round_U197  ( .A(rnd_q[117]), .B(rnd_q[85]), .Z(_sha1_round_n369 ) );
XOR2_X2 _sha1_round_U196  ( .A(rnd_q[110]), .B(rnd_q[78]), .Z(_sha1_round_n368 ) );
XOR2_X2 _sha1_round_U195  ( .A(rnd_q[106]), .B(rnd_q[74]), .Z(_sha1_round_n367 ) );
XOR2_X2 _sha1_round_U194  ( .A(rnd_q[116]), .B(rnd_q[84]), .Z(_sha1_round_n366 ) );
XOR2_X2 _sha1_round_U193  ( .A(rnd_q[101]), .B(rnd_q[69]), .Z(_sha1_round_n365 ) );
NAND2_X1 _sha1_round_U192  ( .A1(_sha1_round_n365 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n752 ) );
NAND2_X4 _sha1_round_U191  ( .A1(_sha1_round_n819 ), .A2(_sha1_round_n820 ),.ZN(_sha1_round_n767 ) );
NAND2_X1 _sha1_round_U190  ( .A1(_sha1_round_n3120 ), .A2(_sha1_round_n820 ),.ZN(_sha1_round_n3170 ) );
INV_X2 _sha1_round_U189  ( .A(_sha1_round_n360 ), .ZN(_sha1_round_n363 ) );
INV_X4 _sha1_round_U188  ( .A(_sha1_round_n3140 ), .ZN(_sha1_round_n510 ) );
INV_X4 _sha1_round_U187  ( .A(_sha1_round_n363 ), .ZN(_sha1_round_n364 ) );
NAND3_X1 _sha1_round_U186  ( .A1(rnd_q[64]), .A2(rnd_q[96]), .A3(_sha1_round_k[3] ), .ZN(_sha1_round_n815 ) );
OR2_X4 _sha1_round_U185  ( .A1(rnd_q[73]), .A2(rnd_q[105]), .ZN(_sha1_round_n362 ) );
NAND2_X4 _sha1_round_U184  ( .A1(_sha1_round_n712 ), .A2(_sha1_round_n713 ),.ZN(_sha1_round_f [11]) );
NAND2_X4 _sha1_round_U183  ( .A1(_sha1_round_n721 ), .A2(_sha1_round_n720 ),.ZN(_sha1_round_f [10]) );
NAND2_X4 _sha1_round_U182  ( .A1(_sha1_round_n753 ), .A2(_sha1_round_n754 ),.ZN(_sha1_round_f [5]) );
NOR2_X1 _sha1_round_U180  ( .A1(_sha1_round_n706 ), .A2(_sha1_round_n3120 ),.ZN(_sha1_round_n708 ) );
NOR2_X1 _sha1_round_U179  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n3210 ),.ZN(_sha1_round_n722 ) );
NOR2_X1 _sha1_round_U177  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n3240 ),.ZN(_sha1_round_n738 ) );
NAND2_X1 _sha1_round_U176  ( .A1(_sha1_round_n372 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n711 ) );
INV_X4 _sha1_round_U175  ( .A(rnd_q[43]), .ZN(_sha1_round_n357 ) );
NAND2_X2 _sha1_round_U174  ( .A1(_sha1_round_n711 ), .A2(_sha1_round_n357 ),.ZN(_sha1_round_n358 ) );
NAND2_X2 _sha1_round_U173  ( .A1(_sha1_round_n3230 ), .A2(_sha1_round_n532 ),.ZN(_sha1_round_n533 ) );
NAND2_X2 _sha1_round_U172  ( .A1(_sha1_round_n367 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n719 ) );
INV_X1 _sha1_round_U170  ( .A(rnd_q[42]), .ZN(_sha1_round_n354 ) );
NAND2_X2 _sha1_round_U169  ( .A1(_sha1_round_n719 ), .A2(_sha1_round_n354 ),.ZN(_sha1_round_n355 ) );
NAND2_X1 _sha1_round_U167  ( .A1(_sha1_round_n3220 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n747 ) );
INV_X1 _sha1_round_U166  ( .A(rnd_q[38]), .ZN(_sha1_round_n351 ) );
NAND2_X2 _sha1_round_U165  ( .A1(_sha1_round_n747 ), .A2(_sha1_round_n351 ),.ZN(_sha1_round_n352 ) );
INV_X1 _sha1_round_U164  ( .A(rnd_q[41]), .ZN(_sha1_round_n348 ) );
NAND2_X2 _sha1_round_U163  ( .A1(_sha1_round_n726 ), .A2(_sha1_round_n348 ),.ZN(_sha1_round_n349 ) );
INV_X1 _sha1_round_U162  ( .A(rnd_q[37]), .ZN(_sha1_round_n3450 ) );
NAND2_X2 _sha1_round_U160  ( .A1(_sha1_round_n752 ), .A2(_sha1_round_n3450 ),.ZN(_sha1_round_n3460 ) );
NAND3_X1 _sha1_round_U159  ( .A1(rnd_q[65]), .A2(rnd_q[97]), .A3(_sha1_round_k[3] ), .ZN(_sha1_round_n802 ) );
NAND2_X4 _sha1_round_U157  ( .A1(_sha1_round_n3250 ), .A2(_sha1_round_n800 ),.ZN(_sha1_round_f [1]) );
NOR2_X1 _sha1_round_U156  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n369 ),.ZN(_sha1_round_n627 ) );
NOR2_X1 _sha1_round_U155  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n373 ),.ZN(_sha1_round_n651 ) );
NAND3_X1 _sha1_round_U154  ( .A1(rnd_q[67]), .A2(rnd_q[99]), .A3(_sha1_round_k[3] ), .ZN(_sha1_round_n776 ) );
NAND3_X1 _sha1_round_U153  ( .A1(rnd_q[66]), .A2(rnd_q[98]), .A3(_sha1_round_k[3] ), .ZN(_sha1_round_n789 ) );
AND2_X2 _sha1_round_U152  ( .A1(_sha1_round_n3150 ), .A2(_sha1_round_n362 ),.ZN(_sha1_round_n723 ) );
NAND2_X1 _sha1_round_U150  ( .A1(_sha1_round_n3150 ), .A2(_sha1_round_n796 ),.ZN(_sha1_round_n797 ) );
NOR2_X2 _sha1_round_U149  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n367 ),.ZN(_sha1_round_n715 ) );
NOR2_X2 _sha1_round_U147  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n372 ),.ZN(_sha1_round_n707 ) );
INV_X2 _sha1_round_U146  ( .A(_sha1_round_n3170 ), .ZN(_sha1_round_n817 ) );
NAND2_X4 _sha1_round_U145  ( .A1(_sha1_round_n736 ), .A2(_sha1_round_n735 ),.ZN(_sha1_round_f [8]) );
OR2_X2 _sha1_round_U144  ( .A1(_sha1_round_n750 ), .A2(_sha1_round_n3120 ),.ZN(_sha1_round_n3420 ) );
OR2_X4 _sha1_round_U143  ( .A1(rnd_q[101]), .A2(_sha1_round_n510 ), .ZN(_sha1_round_n3410 ) );
AND3_X4 _sha1_round_U142  ( .A1(_sha1_round_n3410 ), .A2(_sha1_round_n3420 ),.A3(_sha1_round_n3430 ), .ZN(_sha1_round_n751 ) );
NAND2_X4 _sha1_round_U140  ( .A1(_sha1_round_n697 ), .A2(_sha1_round_n696 ),.ZN(_sha1_round_f [13]) );
NAND2_X2 _sha1_round_U139  ( .A1(_sha1_round_n531 ), .A2(_sha1_round_n524 ),.ZN(_sha1_round_n522 ) );
NAND2_X2 _sha1_round_U137  ( .A1(_sha1_round_n524 ), .A2(_sha1_round_n523 ),.ZN(_sha1_round_n526 ) );
OR2_X1 _sha1_round_U136  ( .A1(_sha1_round_n745 ), .A2(_sha1_round_n3160 ),.ZN(_sha1_round_n3390 ) );
OR2_X1 _sha1_round_U135  ( .A1(rnd_q[102]), .A2(_sha1_round_n510 ), .ZN(_sha1_round_n3380 ) );
AND3_X4 _sha1_round_U134  ( .A1(_sha1_round_n3380 ), .A2(_sha1_round_n3390 ),.A3(_sha1_round_n3400 ), .ZN(_sha1_round_n746 ) );
NAND2_X2 _sha1_round_U133  ( .A1(_sha1_round_n3150 ), .A2(_sha1_round_n770 ),.ZN(_sha1_round_n771 ) );
INV_X2 _sha1_round_U132  ( .A(rnd_q[33]), .ZN(_sha1_round_n791 ) );
NOR2_X2 _sha1_round_U130  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n374 ),.ZN(_sha1_round_n757 ) );
NOR2_X2 _sha1_round_U129  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n379 ),.ZN(_sha1_round_n667 ) );
NOR2_X2 _sha1_round_U127  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n375 ),.ZN(_sha1_round_n675 ) );
INV_X1 _sha1_round_U126  ( .A(_sha1_round_n819 ), .ZN(_sha1_round_n825 ) );
OR2_X2 _sha1_round_U125  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n3220 ),.ZN(_sha1_round_n3400 ) );
OR2_X2 _sha1_round_U124  ( .A1(_sha1_round_n756 ), .A2(_sha1_round_n365 ),.ZN(_sha1_round_n3430 ) );
NAND2_X1 _sha1_round_U123  ( .A1(rnd_cnt_q[6]), .A2(rnd_cnt_q[5]), .ZN(_sha1_round_n535 ) );
NAND3_X2 _sha1_round_U122  ( .A1(rnd_cnt_q[5]), .A2(_sha1_round_n531 ), .A3(_sha1_round_n524 ), .ZN(_sha1_round_n528 ) );
NAND2_X1 _sha1_round_U120  ( .A1(_sha1_round_n370 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n734 ) );
NAND2_X1 _sha1_round_U119  ( .A1(_sha1_round_n366 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n639 ) );
NAND2_X2 _sha1_round_U117  ( .A1(_sha1_round_n3210 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n726 ) );
NAND2_X1 _sha1_round_U116  ( .A1(_sha1_round_n368 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n687 ) );
NAND2_X1 _sha1_round_U115  ( .A1(_sha1_round_n371 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n647 ) );
NAND2_X1 _sha1_round_U114  ( .A1(_sha1_round_n379 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n671 ) );
NAND2_X1 _sha1_round_U113  ( .A1(_sha1_round_n375 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n679 ) );
NAND2_X1 _sha1_round_U112  ( .A1(_sha1_round_n378 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n703 ) );
NAND3_X1 _sha1_round_U111  ( .A1(rnd_q[34]), .A2(_sha1_round_n515 ), .A3(_sha1_round_n780 ), .ZN(_sha1_round_n788 ) );
NAND2_X1 _sha1_round_U110  ( .A1(_sha1_round_n377 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n695 ) );
NAND3_X1 _sha1_round_U109  ( .A1(_sha1_round_n779 ), .A2(_sha1_round_n778 ),.A3(_sha1_round_n515 ), .ZN(_sha1_round_n790 ) );
NAND2_X1 _sha1_round_U108  ( .A1(_sha1_round_n369 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n631 ) );
NAND2_X1 _sha1_round_U107  ( .A1(_sha1_round_n168 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n612 ) );
NAND2_X1 _sha1_round_U106  ( .A1(_sha1_round_n373 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n655 ) );
NAND2_X1 _sha1_round_U105  ( .A1(_sha1_round_n159 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n603 ) );
NAND2_X1 _sha1_round_U104  ( .A1(_sha1_round_n376 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n663 ) );
NAND2_X1 _sha1_round_U103  ( .A1(_sha1_round_n380 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n623 ) );
INV_X1 _sha1_round_U102  ( .A(rnd_q[40]), .ZN(_sha1_round_n3340 ) );
NAND2_X2 _sha1_round_U100  ( .A1(_sha1_round_n734 ), .A2(_sha1_round_n3340 ),.ZN(_sha1_round_n3350 ) );
NAND2_X4 _sha1_round_U99  ( .A1(_sha1_round_n705 ), .A2(_sha1_round_n704 ),.ZN(_sha1_round_f [12]) );
NOR2_X2 _sha1_round_U97  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n377 ),.ZN(_sha1_round_n691 ) );
NAND2_X2 _sha1_round_U96  ( .A1(_sha1_round_n3270 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n814 ) );
INV_X4 _sha1_round_U95  ( .A(rnd_q[39]), .ZN(_sha1_round_n3440 ) );
NAND2_X1 _sha1_round_U94  ( .A1(_sha1_round_n3240 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n742 ) );
INV_X4 _sha1_round_U93  ( .A(_sha1_round_n3440 ), .ZN(sha1_round_wire[7]) );
NAND2_X2 _sha1_round_U92  ( .A1(_sha1_round_n742 ), .A2(_sha1_round_n3440 ),.ZN(_sha1_round_n3330 ) );
NAND2_X2 _sha1_round_U90  ( .A1(_sha1_round_n741 ), .A2(sha1_round_wire[7]),.ZN(_sha1_round_n3320 ) );
INV_X4 _sha1_round_U89  ( .A(_sha1_round_k[3] ), .ZN(_sha1_round_n518 ) );
INV_X2 _sha1_round_U87  ( .A(_sha1_round_n518 ), .ZN(_sha1_round_n3300 ) );
INV_X4 _sha1_round_U86  ( .A(rnd_cnt_q[5]), .ZN(_sha1_round_n525 ) );
AND2_X4 _sha1_round_U85  ( .A1(_sha1_round_n804 ), .A2(_sha1_round_n805 ),.ZN(_sha1_round_n3290 ) );
AND2_X4 _sha1_round_U84  ( .A1(_sha1_round_n791 ), .A2(_sha1_round_n792 ),.ZN(_sha1_round_n3280 ) );
AND2_X4 _sha1_round_U83  ( .A1(rnd_q[32]), .A2(_sha1_round_n806 ), .ZN(_sha1_round_n3270 ) );
OR2_X2 _sha1_round_U82  ( .A1(_sha1_round_n723 ), .A2(_sha1_round_n724 ),.ZN(_sha1_round_n3260 ) );
XOR2_X2 _sha1_round_U81  ( .A(rnd_q[103]), .B(rnd_q[71]), .Z(_sha1_round_n3240 ) );
AND2_X4 _sha1_round_U80  ( .A1(n7119), .A2(rnd_cnt_q[5]), .ZN(_sha1_round_n3230 ) );
XOR2_X2 _sha1_round_U79  ( .A(rnd_q[102]), .B(rnd_q[70]), .Z(_sha1_round_n3220 ) );
XOR2_X2 _sha1_round_U78  ( .A(rnd_q[105]), .B(rnd_q[73]), .Z(_sha1_round_n3210 ) );
BUF_X4 _sha1_round_U77  ( .A(_sha1_round_n515 ), .Z(_sha1_round_n3370 ) );
NAND2_X1 _sha1_round_U76  ( .A1(n7119), .A2(rnd_cnt_q[4]), .ZN(_sha1_round_n519 ) );
NAND2_X4 _sha1_round_U75  ( .A1(_sha1_round_n358 ), .A2(_sha1_round_n359 ),.ZN(_sha1_round_n712 ) );
NAND2_X2 _sha1_round_U74  ( .A1(_sha1_round_n532 ), .A2(n7119), .ZN(_sha1_round_n521 ) );
NAND3_X2 _sha1_round_U73  ( .A1(rnd_q[33]), .A2(_sha1_round_n515 ), .A3(_sha1_round_n793 ), .ZN(_sha1_round_n801 ) );
NAND2_X2 _sha1_round_U72  ( .A1(_sha1_round_n641 ), .A2(_sha1_round_n640 ),.ZN(_sha1_round_f [20]) );
NAND2_X2 _sha1_round_U71  ( .A1(_sha1_round_n689 ), .A2(_sha1_round_n688 ),.ZN(_sha1_round_f [14]) );
NAND2_X2 _sha1_round_U70  ( .A1(_sha1_round_n510 ), .A2(_sha1_round_n817 ),.ZN(_sha1_round_n2 ) );
NAND2_X2 _sha1_round_U69  ( .A1(rnd_q[33]), .A2(_sha1_round_n799 ), .ZN(_sha1_round_n800 ) );
NAND2_X2 _sha1_round_U68  ( .A1(rnd_q[35]), .A2(_sha1_round_n773 ), .ZN(_sha1_round_n774 ) );
NAND2_X2 _sha1_round_U67  ( .A1(_sha1_round_n718 ), .A2(rnd_q[42]), .ZN(_sha1_round_n356 ) );
NAND2_X2 _sha1_round_U66  ( .A1(_sha1_round_n733 ), .A2(rnd_q[40]), .ZN(_sha1_round_n3360 ) );
NOR2_X2 _sha1_round_U65  ( .A1(_sha1_round_n722 ), .A2(_sha1_round_n3260 ),.ZN(_sha1_round_n725 ) );
NAND2_X2 _sha1_round_U64  ( .A1(_sha1_round_n725 ), .A2(rnd_q[41]), .ZN(_sha1_round_n350 ) );
NAND2_X2 _sha1_round_U63  ( .A1(_sha1_round_n746 ), .A2(rnd_q[38]), .ZN(_sha1_round_n353 ) );
NOR3_X2 _sha1_round_U62  ( .A1(_sha1_round_n709 ), .A2(_sha1_round_n708 ),.A3(_sha1_round_n707 ), .ZN(_sha1_round_n710 ) );
NAND2_X2 _sha1_round_U61  ( .A1(_sha1_round_n349 ), .A2(_sha1_round_n350 ),.ZN(_sha1_round_n727 ) );
NOR2_X2 _sha1_round_U60  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n366 ),.ZN(_sha1_round_n635 ) );
INV_X1 _sha1_round_U59  ( .A(_sha1_round_n514 ), .ZN(_sha1_round_n360 ) );
INV_X8 _sha1_round_U58  ( .A(_sha1_round_n512 ), .ZN(_sha1_round_n514 ) );
NAND4_X4 _sha1_round_U57  ( .A1(_sha1_round_n777 ), .A2(_sha1_round_n776 ),.A3(_sha1_round_n775 ), .A4(_sha1_round_n774 ), .ZN(_sha1_round_f [3]));
NOR2_X1 _sha1_round_U56  ( .A1(rnd_q[107]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n709 ) );
NOR2_X1 _sha1_round_U55  ( .A1(rnd_q[116]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n637 ) );
NOR2_X1 _sha1_round_U54  ( .A1(rnd_q[104]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n732 ) );
NOR2_X1 _sha1_round_U53  ( .A1(rnd_q[115]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n645 ) );
NOR2_X1 _sha1_round_U52  ( .A1(rnd_q[108]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n701 ) );
NOR2_X1 _sha1_round_U51  ( .A1(rnd_q[117]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n629 ) );
NOR2_X1 _sha1_round_U50  ( .A1(rnd_q[113]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n661 ) );
NOR2_X1 _sha1_round_U49  ( .A1(rnd_q[118]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n621 ) );
NOR2_X1 _sha1_round_U48  ( .A1(rnd_q[114]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n653 ) );
NAND2_X4 _sha1_round_U47  ( .A1(_sha1_round_n352 ), .A2(_sha1_round_n353 ),.ZN(_sha1_round_n748 ) );
INV_X8 _sha1_round_U46  ( .A(_sha1_round_n767 ), .ZN(_sha1_round_n756 ) );
INV_X4 _sha1_round_U45  ( .A(n7119), .ZN(_sha1_round_n523 ) );
NAND4_X2 _sha1_round_U44  ( .A1(_sha1_round_n521 ), .A2(_sha1_round_n529 ),.A3(_sha1_round_n522 ), .A4(rnd_cnt_q[5]), .ZN(_sha1_round_n822 ) );
NAND3_X2 _sha1_round_U43  ( .A1(_sha1_round_n525 ), .A2(_sha1_round_n526 ),.A3(rnd_cnt_q[4]), .ZN(_sha1_round_n527 ) );
NAND2_X2 _sha1_round_U42  ( .A1(_sha1_round_n528 ), .A2(_sha1_round_n527 ),.ZN(_sha1_round_n530 ) );
AND4_X4 _sha1_round_U41  ( .A1(_sha1_round_n520 ), .A2(_sha1_round_n529 ),.A3(_sha1_round_n519 ), .A4(_sha1_round_n525 ), .ZN(_sha1_round_n3140 ) );
INV_X4 _sha1_round_U40  ( .A(_sha1_round_n508 ), .ZN(_sha1_round_n509 ) );
NAND3_X2 _sha1_round_U39  ( .A1(_sha1_round_n3130 ), .A2(_sha1_round_n815 ),.A3(_sha1_round_n813 ), .ZN(_sha1_round_f [0]) );
INV_X4 _sha1_round_U38  ( .A(rnd_cnt_q[6]), .ZN(_sha1_round_n529 ) );
INV_X4 _sha1_round_U37  ( .A(_sha1_round_n3150 ), .ZN(_sha1_round_n3160 ) );
INV_X8 _sha1_round_U36  ( .A(_sha1_round_n3160 ), .ZN(_sha1_round_n512 ) );
INV_X8 _sha1_round_U35  ( .A(_sha1_round_n518 ), .ZN(_sha1_round_n517 ) );
NAND2_X2 _sha1_round_U34  ( .A1(_sha1_round_n762 ), .A2(_sha1_round_n763 ),.ZN(_sha1_round_f [4]) );
NAND4_X2 _sha1_round_U33  ( .A1(_sha1_round_n790 ), .A2(_sha1_round_n788 ),.A3(_sha1_round_n789 ), .A4(_sha1_round_n787 ), .ZN(_sha1_round_f [2]));
NAND2_X2 _sha1_round_U32  ( .A1(_sha1_round_n355 ), .A2(_sha1_round_n356 ),.ZN(_sha1_round_n720 ) );
NAND2_X2 _sha1_round_U31  ( .A1(_sha1_round_n3320 ), .A2(_sha1_round_n3330 ),.ZN(_sha1_round_n743 ) );
NAND2_X2 _sha1_round_U30  ( .A1(_sha1_round_n744 ), .A2(_sha1_round_n743 ),.ZN(_sha1_round_f [7]) );
NAND2_X2 _sha1_round_U29  ( .A1(_sha1_round_n710 ), .A2(rnd_q[43]), .ZN(_sha1_round_n359 ) );
NOR2_X2 _sha1_round_U28  ( .A1(_sha1_round_n516 ), .A2(_sha1_round_n370 ),.ZN(_sha1_round_n730 ) );
INV_X8 _sha1_round_U27  ( .A(_sha1_round_n3140 ), .ZN(_sha1_round_n361 ) );
NOR2_X2 _sha1_round_U26  ( .A1(rnd_q[109]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n693 ) );
NOR2_X2 _sha1_round_U25  ( .A1(rnd_q[110]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n685 ) );
NOR2_X2 _sha1_round_U24  ( .A1(rnd_q[111]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n677 ) );
NOR2_X1 _sha1_round_U23  ( .A1(rnd_q[105]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n724 ) );
NOR2_X2 _sha1_round_U22  ( .A1(rnd_q[112]), .A2(_sha1_round_n361 ), .ZN(_sha1_round_n669 ) );
INV_X16 _sha1_round_U21  ( .A(_sha1_round_n361 ), .ZN(_sha1_round_n511 ) );
INV_X8 _sha1_round_U20  ( .A(_sha1_round_n822 ), .ZN(_sha1_round_n3150 ) );
INV_X2 _sha1_round_U19  ( .A(_sha1_round_n512 ), .ZN(_sha1_round_n3200 ) );
INV_X2 _sha1_round_U18  ( .A(_sha1_round_n512 ), .ZN(_sha1_round_n513 ) );
INV_X2 _sha1_round_U17  ( .A(_sha1_round_n512 ), .ZN(_sha1_round_n3190 ) );
INV_X4 _sha1_round_U16  ( .A(_sha1_round_n3150 ), .ZN(_sha1_round_n3180 ) );
NAND4_X2 _sha1_round_U15  ( .A1(_sha1_round_n521 ), .A2(_sha1_round_n529 ),.A3(_sha1_round_n522 ), .A4(rnd_cnt_q[5]), .ZN(_sha1_round_n3120 ) );
INV_X8 _sha1_round_U14  ( .A(rnd_cnt_q[4]), .ZN(_sha1_round_n531 ) );
NAND2_X4 _sha1_round_U13  ( .A1(rnd_cnt_q[3]), .A2(rnd_cnt_q[4]), .ZN(_sha1_round_n520 ) );
NOR3_X4 _sha1_round_U12  ( .A1(_sha1_round_n717 ), .A2(_sha1_round_n716 ),.A3(_sha1_round_n715 ), .ZN(_sha1_round_n718 ) );
NAND2_X2 _sha1_round_U11  ( .A1(_sha1_round_n3280 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n803 ) );
NOR3_X4 _sha1_round_U10  ( .A1(_sha1_round_n732 ), .A2(_sha1_round_n731 ),.A3(_sha1_round_n730 ), .ZN(_sha1_round_n733 ) );
NAND2_X2 _sha1_round_U9  ( .A1(_sha1_round_n3350 ), .A2(_sha1_round_n3360 ),.ZN(_sha1_round_n735 ) );
AND3_X4 _sha1_round_U8  ( .A1(_sha1_round_n801 ), .A2(_sha1_round_n803 ),.A3(_sha1_round_n802 ), .ZN(_sha1_round_n3250 ) );
NAND2_X2 _sha1_round_U7  ( .A1(_sha1_round_n3290 ), .A2(_sha1_round_n515 ),.ZN(_sha1_round_n816 ) );
AND2_X2 _sha1_round_U6  ( .A1(_sha1_round_n816 ), .A2(_sha1_round_n814 ),.ZN(_sha1_round_n3130 ) );
NAND2_X4 _sha1_round_U5  ( .A1(_sha1_round_n751 ), .A2(rnd_q[37]), .ZN(_sha1_round_n3470 ) );
NAND2_X4 _sha1_round_U3  ( .A1(_sha1_round_n3470 ), .A2(_sha1_round_n3460 ),.ZN(_sha1_round_n753 ) );
XNOR2_X2 _sha1_round_U181  ( .A(rnd_q[87]), .B(rnd_q[119]), .ZN(_sha1_round_n168 ) );
OR2_X2 _sha1_round_U178  ( .A1(rnd_q[87]), .A2(rnd_q[119]), .ZN(_sha1_round_n167 ) );
XNOR2_X2 _sha1_round_U171  ( .A(rnd_q[88]), .B(rnd_q[120]), .ZN(_sha1_round_n159 ) );
OR2_X2 _sha1_round_U168  ( .A1(rnd_q[88]), .A2(rnd_q[120]), .ZN(_sha1_round_n158 ) );
XNOR2_X2 _sha1_round_U161  ( .A(rnd_q[89]), .B(rnd_q[121]), .ZN(_sha1_round_n150 ) );
OR2_X2 _sha1_round_U158  ( .A1(rnd_q[89]), .A2(rnd_q[121]), .ZN(_sha1_round_n149 ) );
XNOR2_X2 _sha1_round_U151  ( .A(rnd_q[90]), .B(rnd_q[122]), .ZN(_sha1_round_n141 ) );
OR2_X2 _sha1_round_U148  ( .A1(rnd_q[90]), .A2(rnd_q[122]), .ZN(_sha1_round_n140 ) );
XNOR2_X2 _sha1_round_U141  ( .A(rnd_q[91]), .B(rnd_q[123]), .ZN(_sha1_round_n132 ) );
OR2_X2 _sha1_round_U138  ( .A1(rnd_q[91]), .A2(rnd_q[123]), .ZN(_sha1_round_n131 ) );
XNOR2_X2 _sha1_round_U131  ( .A(rnd_q[92]), .B(rnd_q[124]), .ZN(_sha1_round_n123 ) );
OR2_X2 _sha1_round_U128  ( .A1(rnd_q[92]), .A2(rnd_q[124]), .ZN(_sha1_round_n122 ) );
XNOR2_X2 _sha1_round_U121  ( .A(rnd_q[93]), .B(rnd_q[125]), .ZN(_sha1_round_n114 ) );
OR2_X2 _sha1_round_U118  ( .A1(rnd_q[93]), .A2(rnd_q[125]), .ZN(_sha1_round_n113 ) );
XNOR2_X2 _sha1_round_U101  ( .A(rnd_q[94]), .B(rnd_q[126]), .ZN(_sha1_round_n96 ) );
OR2_X2 _sha1_round_U98  ( .A1(rnd_q[94]), .A2(rnd_q[126]), .ZN(_sha1_round_n95 ) );
XNOR2_X2 _sha1_round_U91  ( .A(rnd_q[95]), .B(rnd_q[127]), .ZN(_sha1_round_n87 ) );
OR2_X2 _sha1_round_U88  ( .A1(rnd_q[95]), .A2(rnd_q[127]), .ZN(_sha1_round_n86 ) );
NAND2_X2 _sha1_round_add_79_4_U377  ( .A1(_sha1_round_N316 ), .A2(rnd_q[155]), .ZN(_sha1_round_add_79_4_n243 ) );
INV_X4 _sha1_round_add_79_4_U376  ( .A(_sha1_round_add_79_4_n56 ), .ZN(_sha1_round_add_79_4_n311 ) );
NAND4_X2 _sha1_round_add_79_4_U375  ( .A1(_sha1_round_N320 ), .A2(rnd_q[159]), .A3(_sha1_round_add_79_4_n336 ), .A4(_sha1_round_add_79_4_n72 ), .ZN(_sha1_round_add_79_4_n341 ) );
NAND2_X2 _sha1_round_add_79_4_U374  ( .A1(_sha1_round_N322 ), .A2(rnd_q[129]), .ZN(_sha1_round_add_79_4_n70 ) );
INV_X4 _sha1_round_add_79_4_U373  ( .A(_sha1_round_add_79_4_n70 ), .ZN(_sha1_round_add_79_4_n344 ) );
INV_X4 _sha1_round_add_79_4_U372  ( .A(_sha1_round_add_79_4_n67 ), .ZN(_sha1_round_add_79_4_n345 ) );
NAND2_X2 _sha1_round_add_79_4_U371  ( .A1(_sha1_round_add_79_4_n316 ), .A2(_sha1_round_add_79_4_n68 ), .ZN(_sha1_round_add_79_4_n280 ) );
INV_X4 _sha1_round_add_79_4_U370  ( .A(_sha1_round_add_79_4_n280 ), .ZN(_sha1_round_add_79_4_n62 ) );
INV_X4 _sha1_round_add_79_4_U369  ( .A(_sha1_round_add_79_4_n60 ), .ZN(_sha1_round_add_79_4_n318 ) );
NAND2_X2 _sha1_round_add_79_4_U368  ( .A1(_sha1_round_add_79_4_n62 ), .A2(_sha1_round_add_79_4_n318 ), .ZN(_sha1_round_add_79_4_n329 ) );
INV_X4 _sha1_round_add_79_4_U367  ( .A(_sha1_round_add_79_4_n75 ), .ZN(_sha1_round_add_79_4_n336 ) );
INV_X4 _sha1_round_add_79_4_U366  ( .A(_sha1_round_add_79_4_n80 ), .ZN(_sha1_round_add_79_4_n337 ) );
INV_X4 _sha1_round_add_79_4_U365  ( .A(_sha1_round_add_79_4_n72 ), .ZN(_sha1_round_add_79_4_n339 ) );
INV_X4 _sha1_round_add_79_4_U364  ( .A(_sha1_round_add_79_4_n64 ), .ZN(_sha1_round_add_79_4_n314 ) );
NAND2_X2 _sha1_round_add_79_4_U363  ( .A1(_sha1_round_N319 ), .A2(rnd_q[158]), .ZN(_sha1_round_add_79_4_n86 ) );
INV_X4 _sha1_round_add_79_4_U362  ( .A(_sha1_round_add_79_4_n90 ), .ZN(_sha1_round_add_79_4_n335 ) );
NAND2_X2 _sha1_round_add_79_4_U361  ( .A1(_sha1_round_add_79_4_n243 ), .A2(_sha1_round_add_79_4_n139 ), .ZN(_sha1_round_add_79_4_n333 ) );
INV_X4 _sha1_round_add_79_4_U360  ( .A(_sha1_round_add_79_4_n85 ), .ZN(_sha1_round_add_79_4_n332 ) );
NAND2_X2 _sha1_round_add_79_4_U359  ( .A1(_sha1_round_N318 ), .A2(rnd_q[157]), .ZN(_sha1_round_add_79_4_n87 ) );
NAND2_X2 _sha1_round_add_79_4_U358  ( .A1(_sha1_round_add_79_4_n311 ), .A2(_sha1_round_add_79_4_n54 ), .ZN(_sha1_round_add_79_4_n328 ) );
NAND2_X2 _sha1_round_add_79_4_U357  ( .A1(_sha1_round_N325 ), .A2(rnd_q[132]), .ZN(_sha1_round_add_79_4_n55 ) );
NAND2_X2 _sha1_round_add_79_4_U356  ( .A1(_sha1_round_add_79_4_n328 ), .A2(_sha1_round_add_79_4_n55 ), .ZN(_sha1_round_add_79_4_n324 ) );
INV_X4 _sha1_round_add_79_4_U355  ( .A(_sha1_round_N326 ), .ZN(_sha1_round_add_79_4_n326 ) );
INV_X4 _sha1_round_add_79_4_U354  ( .A(rnd_q[133]), .ZN(_sha1_round_add_79_4_n327 ) );
NAND2_X2 _sha1_round_add_79_4_U353  ( .A1(_sha1_round_N326 ), .A2(rnd_q[133]), .ZN(_sha1_round_add_79_4_n308 ) );
NAND2_X2 _sha1_round_add_79_4_U352  ( .A1(_sha1_round_add_79_4_n313 ), .A2(_sha1_round_add_79_4_n308 ), .ZN(_sha1_round_add_79_4_n325 ) );
XNOR2_X2 _sha1_round_add_79_4_U351  ( .A(_sha1_round_add_79_4_n324 ), .B(_sha1_round_add_79_4_n325 ), .ZN(sha1_round_wire[138]) );
NAND2_X2 _sha1_round_add_79_4_U350  ( .A1(_sha1_round_add_79_4_n324 ), .A2(_sha1_round_add_79_4_n313 ), .ZN(_sha1_round_add_79_4_n323 ) );
NAND2_X2 _sha1_round_add_79_4_U349  ( .A1(_sha1_round_add_79_4_n308 ), .A2(_sha1_round_add_79_4_n323 ), .ZN(_sha1_round_add_79_4_n319 ) );
INV_X4 _sha1_round_add_79_4_U348  ( .A(rnd_q[134]), .ZN(_sha1_round_add_79_4_n322 ) );
XNOR2_X2 _sha1_round_add_79_4_U347  ( .A(_sha1_round_add_79_4_n319 ), .B(_sha1_round_add_79_4_n320 ), .ZN(sha1_round_wire[139]) );
NAND2_X2 _sha1_round_add_79_4_U346  ( .A1(_sha1_round_add_79_4_n312 ), .A2(_sha1_round_add_79_4_n55 ), .ZN(_sha1_round_add_79_4_n310 ) );
INV_X4 _sha1_round_add_79_4_U345  ( .A(_sha1_round_add_79_4_n308 ), .ZN(_sha1_round_add_79_4_n306 ) );
NAND2_X2 _sha1_round_add_79_4_U344  ( .A1(_sha1_round_N328 ), .A2(rnd_q[135]), .ZN(_sha1_round_add_79_4_n296 ) );
INV_X4 _sha1_round_add_79_4_U343  ( .A(_sha1_round_add_79_4_n296 ), .ZN(_sha1_round_add_79_4_n275 ) );
XNOR2_X2 _sha1_round_add_79_4_U342  ( .A(_sha1_round_add_79_4_n297 ), .B(_sha1_round_add_79_4_n301 ), .ZN(sha1_round_wire[140]) );
NAND2_X2 _sha1_round_add_79_4_U341  ( .A1(_sha1_round_N329 ), .A2(rnd_q[136]), .ZN(_sha1_round_add_79_4_n271 ) );
XNOR2_X2 _sha1_round_add_79_4_U340  ( .A(_sha1_round_add_79_4_n299 ), .B(_sha1_round_add_79_4_n45 ), .ZN(sha1_round_wire[141]) );
INV_X4 _sha1_round_add_79_4_U339  ( .A(_sha1_round_add_79_4_n298 ), .ZN(_sha1_round_add_79_4_n278 ) );
INV_X4 _sha1_round_add_79_4_U338  ( .A(rnd_q[138]), .ZN(_sha1_round_add_79_4_n289 ) );
INV_X4 _sha1_round_add_79_4_U337  ( .A(_sha1_round_add_79_4_n233 ), .ZN(_sha1_round_add_79_4_n269 ) );
XNOR2_X2 _sha1_round_add_79_4_U336  ( .A(_sha1_round_add_79_4_n286 ), .B(_sha1_round_add_79_4_n287 ), .ZN(sha1_round_wire[143]) );
NOR2_X4 _sha1_round_add_79_4_U335  ( .A1(rnd_q[139]), .A2(_sha1_round_n509 ),.ZN(_sha1_round_add_79_4_n254 ) );
INV_X4 _sha1_round_add_79_4_U334  ( .A(_sha1_round_add_79_4_n86 ), .ZN(_sha1_round_add_79_4_n284 ) );
INV_X4 _sha1_round_add_79_4_U333  ( .A(_sha1_round_add_79_4_n149 ), .ZN(_sha1_round_add_79_4_n272 ) );
NOR2_X4 _sha1_round_add_79_4_U332  ( .A1(_sha1_round_add_79_4_n269 ), .A2(_sha1_round_add_79_4_n49 ), .ZN(_sha1_round_add_79_4_n277 ) );
INV_X4 _sha1_round_add_79_4_U331  ( .A(_sha1_round_N333 ), .ZN(_sha1_round_add_79_4_n263 ) );
INV_X4 _sha1_round_add_79_4_U330  ( .A(rnd_q[140]), .ZN(_sha1_round_add_79_4_n264 ) );
XNOR2_X2 _sha1_round_add_79_4_U329  ( .A(_sha1_round_add_79_4_n262 ), .B(_sha1_round_add_79_4_n39 ), .ZN(sha1_round_wire[145]) );
INV_X4 _sha1_round_add_79_4_U328  ( .A(_sha1_round_add_79_4_n247 ), .ZN(_sha1_round_add_79_4_n257 ) );
XNOR2_X2 _sha1_round_add_79_4_U327  ( .A(_sha1_round_add_79_4_n255 ), .B(_sha1_round_add_79_4_n256 ), .ZN(sha1_round_wire[146]) );
XNOR2_X2 _sha1_round_add_79_4_U326  ( .A(_sha1_round_add_79_4_n244 ), .B(_sha1_round_add_79_4_n38 ), .ZN(sha1_round_wire[147]) );
NAND2_X2 _sha1_round_add_79_4_U325  ( .A1(_sha1_round_N317 ), .A2(rnd_q[156]), .ZN(_sha1_round_add_79_4_n139 ) );
INV_X4 _sha1_round_add_79_4_U324  ( .A(_sha1_round_add_79_4_n139 ), .ZN(_sha1_round_add_79_4_n242 ) );
XNOR2_X2 _sha1_round_add_79_4_U323  ( .A(_sha1_round_add_79_4_n243 ), .B(_sha1_round_add_79_4_n241 ), .ZN(sha1_round_wire[129]) );
NOR2_X4 _sha1_round_add_79_4_U322  ( .A1(_sha1_round_add_79_4_n231 ), .A2(_sha1_round_add_79_4_n232 ), .ZN(_sha1_round_add_79_4_n216 ) );
INV_X4 _sha1_round_add_79_4_U321  ( .A(_sha1_round_N337 ), .ZN(_sha1_round_add_79_4_n227 ) );
INV_X4 _sha1_round_add_79_4_U320  ( .A(rnd_q[144]), .ZN(_sha1_round_add_79_4_n228 ) );
XNOR2_X2 _sha1_round_add_79_4_U319  ( .A(_sha1_round_add_79_4_n226 ), .B(_sha1_round_add_79_4_n40 ), .ZN(sha1_round_wire[149]) );
NAND2_X2 _sha1_round_add_79_4_U318  ( .A1(rnd_q[143]), .A2(_sha1_round_N336 ), .ZN(_sha1_round_add_79_4_n224 ) );
NAND2_X2 _sha1_round_add_79_4_U317  ( .A1(_sha1_round_add_79_4_n220 ), .A2(_sha1_round_add_79_4_n204 ), .ZN(_sha1_round_add_79_4_n223 ) );
NAND2_X2 _sha1_round_add_79_4_U316  ( .A1(_sha1_round_N338 ), .A2(rnd_q[145]), .ZN(_sha1_round_add_79_4_n201 ) );
XNOR2_X2 _sha1_round_add_79_4_U315  ( .A(_sha1_round_add_79_4_n221 ), .B(_sha1_round_add_79_4_n46 ), .ZN(sha1_round_wire[150]) );
NAND2_X2 _sha1_round_add_79_4_U314  ( .A1(_sha1_round_add_79_4_n223 ), .A2(_sha1_round_add_79_4_n203 ), .ZN(_sha1_round_add_79_4_n215 ) );
NAND2_X2 _sha1_round_add_79_4_U313  ( .A1(_sha1_round_add_79_4_n217 ), .A2(_sha1_round_add_79_4_n203 ), .ZN(_sha1_round_add_79_4_n212 ) );
NAND2_X2 _sha1_round_add_79_4_U312  ( .A1(_sha1_round_N339 ), .A2(rnd_q[146]), .ZN(_sha1_round_add_79_4_n155 ) );
NAND2_X2 _sha1_round_add_79_4_U311  ( .A1(_sha1_round_add_79_4_n155 ), .A2(_sha1_round_add_79_4_n154 ), .ZN(_sha1_round_add_79_4_n214 ) );
INV_X4 _sha1_round_add_79_4_U310  ( .A(_sha1_round_add_79_4_n212 ), .ZN(_sha1_round_add_79_4_n211 ) );
NAND3_X2 _sha1_round_add_79_4_U309  ( .A1(_sha1_round_add_79_4_n209 ), .A2(_sha1_round_add_79_4_n210 ), .A3(_sha1_round_add_79_4_n136 ), .ZN(_sha1_round_add_79_4_n206 ) );
NAND2_X2 _sha1_round_add_79_4_U308  ( .A1(_sha1_round_add_79_4_n220 ), .A2(_sha1_round_add_79_4_n204 ), .ZN(_sha1_round_add_79_4_n202 ) );
NAND2_X2 _sha1_round_add_79_4_U307  ( .A1(_sha1_round_add_79_4_n202 ), .A2(_sha1_round_add_79_4_n203 ), .ZN(_sha1_round_add_79_4_n200 ) );
NAND2_X2 _sha1_round_add_79_4_U306  ( .A1(_sha1_round_add_79_4_n199 ), .A2(_sha1_round_add_79_4_n155 ), .ZN(_sha1_round_add_79_4_n198 ) );
NAND2_X2 _sha1_round_add_79_4_U305  ( .A1(_sha1_round_add_79_4_n149 ), .A2(_sha1_round_add_79_4_n196 ), .ZN(_sha1_round_add_79_4_n195 ) );
NAND2_X2 _sha1_round_add_79_4_U304  ( .A1(_sha1_round_N340 ), .A2(rnd_q[147]), .ZN(_sha1_round_add_79_4_n185 ) );
INV_X4 _sha1_round_add_79_4_U303  ( .A(rnd_q[147]), .ZN(_sha1_round_add_79_4_n193 ) );
NAND2_X2 _sha1_round_add_79_4_U302  ( .A1(_sha1_round_add_79_4_n185 ), .A2(_sha1_round_add_79_4_n178 ), .ZN(_sha1_round_add_79_4_n191 ) );
NAND2_X2 _sha1_round_add_79_4_U301  ( .A1(_sha1_round_add_79_4_n190 ), .A2(_sha1_round_add_79_4_n185 ), .ZN(_sha1_round_add_79_4_n186 ) );
INV_X4 _sha1_round_add_79_4_U300  ( .A(_sha1_round_N341 ), .ZN(_sha1_round_add_79_4_n188 ) );
INV_X4 _sha1_round_add_79_4_U299  ( .A(rnd_q[148]), .ZN(_sha1_round_add_79_4_n189 ) );
XNOR2_X2 _sha1_round_add_79_4_U298  ( .A(_sha1_round_add_79_4_n186 ), .B(_sha1_round_add_79_4_n187 ), .ZN(sha1_round_wire[153]) );
NAND2_X2 _sha1_round_add_79_4_U297  ( .A1(_sha1_round_add_79_4_n184 ), .A2(_sha1_round_add_79_4_n185 ), .ZN(_sha1_round_add_79_4_n183 ) );
NAND2_X2 _sha1_round_add_79_4_U296  ( .A1(_sha1_round_add_79_4_n174 ), .A2(_sha1_round_add_79_4_n172 ), .ZN(_sha1_round_add_79_4_n181 ) );
XNOR2_X2 _sha1_round_add_79_4_U295  ( .A(_sha1_round_add_79_4_n180 ), .B(_sha1_round_add_79_4_n181 ), .ZN(sha1_round_wire[154]) );
INV_X4 _sha1_round_add_79_4_U294  ( .A(_sha1_round_add_79_4_n179 ), .ZN(_sha1_round_add_79_4_n175 ) );
INV_X4 _sha1_round_add_79_4_U293  ( .A(_sha1_round_add_79_4_n178 ), .ZN(_sha1_round_add_79_4_n177 ) );
NOR3_X4 _sha1_round_add_79_4_U292  ( .A1(_sha1_round_add_79_4_n175 ), .A2(_sha1_round_add_79_4_n176 ), .A3(_sha1_round_add_79_4_n177 ), .ZN(_sha1_round_add_79_4_n156 ) );
NAND2_X2 _sha1_round_add_79_4_U291  ( .A1(_sha1_round_add_79_4_n173 ), .A2(_sha1_round_add_79_4_n174 ), .ZN(_sha1_round_add_79_4_n171 ) );
INV_X4 _sha1_round_add_79_4_U290  ( .A(rnd_q[150]), .ZN(_sha1_round_add_79_4_n169 ) );
XNOR2_X2 _sha1_round_add_79_4_U289  ( .A(_sha1_round_add_79_4_n166 ), .B(_sha1_round_add_79_4_n167 ), .ZN(sha1_round_wire[155]) );
XNOR2_X2 _sha1_round_add_79_4_U288  ( .A(_sha1_round_add_79_4_n159 ), .B(_sha1_round_add_79_4_n160 ), .ZN(sha1_round_wire[156]) );
NOR3_X4 _sha1_round_add_79_4_U287  ( .A1(_sha1_round_add_79_4_n272 ), .A2(_sha1_round_add_79_4_n147 ), .A3(_sha1_round_add_79_4_n148 ), .ZN(_sha1_round_add_79_4_n99 ) );
NAND2_X2 _sha1_round_add_79_4_U286  ( .A1(_sha1_round_add_79_4_n42 ), .A2(_sha1_round_add_79_4_n139 ), .ZN(_sha1_round_add_79_4_n89 ) );
NAND2_X2 _sha1_round_add_79_4_U285  ( .A1(_sha1_round_add_79_4_n90 ), .A2(_sha1_round_add_79_4_n87 ), .ZN(_sha1_round_add_79_4_n138 ) );
XNOR2_X2 _sha1_round_add_79_4_U284  ( .A(_sha1_round_add_79_4_n89 ), .B(_sha1_round_add_79_4_n138 ), .ZN(sha1_round_wire[130]) );
INV_X4 _sha1_round_add_79_4_U283  ( .A(_sha1_round_add_79_4_n131 ), .ZN(_sha1_round_add_79_4_n129 ) );
INV_X4 _sha1_round_add_79_4_U282  ( .A(_sha1_round_add_79_4_n106 ), .ZN(_sha1_round_add_79_4_n128 ) );
INV_X4 _sha1_round_add_79_4_U281  ( .A(_sha1_round_add_79_4_n105 ), .ZN(_sha1_round_add_79_4_n126 ) );
NAND3_X2 _sha1_round_add_79_4_U280  ( .A1(_sha1_round_add_79_4_n123 ), .A2(_sha1_round_add_79_4_n124 ), .A3(_sha1_round_add_79_4_n125 ), .ZN(_sha1_round_add_79_4_n122 ) );
INV_X4 _sha1_round_add_79_4_U279  ( .A(_sha1_round_add_79_4_n116 ), .ZN(_sha1_round_add_79_4_n120 ) );
XNOR2_X2 _sha1_round_add_79_4_U278  ( .A(_sha1_round_add_79_4_n118 ), .B(_sha1_round_add_79_4_n119 ), .ZN(sha1_round_wire[158]) );
NAND2_X2 _sha1_round_add_79_4_U277  ( .A1(_sha1_round_add_79_4_n116 ), .A2(_sha1_round_add_79_4_n117 ), .ZN(_sha1_round_add_79_4_n114 ) );
NAND2_X2 _sha1_round_add_79_4_U276  ( .A1(_sha1_round_add_79_4_n108 ), .A2(_sha1_round_add_79_4_n109 ), .ZN(_sha1_round_add_79_4_n102 ) );
INV_X4 _sha1_round_add_79_4_U275  ( .A(_sha1_round_add_79_4_n99 ), .ZN(_sha1_round_add_79_4_n98 ) );
XNOR2_X2 _sha1_round_add_79_4_U274  ( .A(rnd_q[154]), .B(_sha1_round_N347 ),.ZN(_sha1_round_add_79_4_n92 ) );
NAND2_X2 _sha1_round_add_79_4_U273  ( .A1(_sha1_round_add_79_4_n89 ), .A2(_sha1_round_add_79_4_n90 ), .ZN(_sha1_round_add_79_4_n88 ) );
NAND2_X2 _sha1_round_add_79_4_U272  ( .A1(_sha1_round_add_79_4_n87 ), .A2(_sha1_round_add_79_4_n88 ), .ZN(_sha1_round_add_79_4_n83 ) );
NAND2_X2 _sha1_round_add_79_4_U271  ( .A1(_sha1_round_add_79_4_n85 ), .A2(_sha1_round_add_79_4_n86 ), .ZN(_sha1_round_add_79_4_n84 ) );
XNOR2_X2 _sha1_round_add_79_4_U270  ( .A(_sha1_round_add_79_4_n83 ), .B(_sha1_round_add_79_4_n84 ), .ZN(sha1_round_wire[131]) );
NAND2_X2 _sha1_round_add_79_4_U269  ( .A1(_sha1_round_N320 ), .A2(rnd_q[159]), .ZN(_sha1_round_add_79_4_n79 ) );
NAND2_X2 _sha1_round_add_79_4_U268  ( .A1(_sha1_round_add_79_4_n337 ), .A2(_sha1_round_add_79_4_n79 ), .ZN(_sha1_round_add_79_4_n82 ) );
XNOR2_X2 _sha1_round_add_79_4_U267  ( .A(_sha1_round_add_79_4_n82 ), .B(_sha1_round_add_79_4_n81 ), .ZN(sha1_round_wire[132]) );
INV_X4 _sha1_round_add_79_4_U266  ( .A(_sha1_round_add_79_4_n81 ), .ZN(_sha1_round_add_79_4_n63 ) );
NAND2_X2 _sha1_round_add_79_4_U265  ( .A1(_sha1_round_N321 ), .A2(rnd_q[128]), .ZN(_sha1_round_add_79_4_n74 ) );
INV_X4 _sha1_round_add_79_4_U264  ( .A(_sha1_round_add_79_4_n74 ), .ZN(_sha1_round_add_79_4_n78 ) );
XNOR2_X2 _sha1_round_add_79_4_U263  ( .A(_sha1_round_add_79_4_n76 ), .B(_sha1_round_add_79_4_n77 ), .ZN(sha1_round_wire[133]) );
NAND2_X2 _sha1_round_add_79_4_U262  ( .A1(_sha1_round_add_79_4_n72 ), .A2(_sha1_round_add_79_4_n70 ), .ZN(_sha1_round_add_79_4_n73 ) );
NAND2_X2 _sha1_round_add_79_4_U261  ( .A1(_sha1_round_add_79_4_n41 ), .A2(_sha1_round_add_79_4_n74 ), .ZN(_sha1_round_add_79_4_n71 ) );
XNOR2_X2 _sha1_round_add_79_4_U260  ( .A(_sha1_round_add_79_4_n73 ), .B(_sha1_round_add_79_4_n71 ), .ZN(sha1_round_wire[134]) );
NAND2_X2 _sha1_round_add_79_4_U259  ( .A1(_sha1_round_add_79_4_n71 ), .A2(_sha1_round_add_79_4_n72 ), .ZN(_sha1_round_add_79_4_n69 ) );
NAND2_X2 _sha1_round_add_79_4_U258  ( .A1(_sha1_round_add_79_4_n69 ), .A2(_sha1_round_add_79_4_n70 ), .ZN(_sha1_round_add_79_4_n65 ) );
NAND2_X2 _sha1_round_add_79_4_U257  ( .A1(_sha1_round_add_79_4_n67 ), .A2(_sha1_round_add_79_4_n68 ), .ZN(_sha1_round_add_79_4_n66 ) );
XNOR2_X2 _sha1_round_add_79_4_U256  ( .A(_sha1_round_add_79_4_n65 ), .B(_sha1_round_add_79_4_n66 ), .ZN(sha1_round_wire[135]) );
INV_X4 _sha1_round_add_79_4_U255  ( .A(_sha1_round_add_79_4_n312 ), .ZN(_sha1_round_add_79_4_n59 ) );
XNOR2_X2 _sha1_round_add_79_4_U254  ( .A(_sha1_round_add_79_4_n57 ), .B(_sha1_round_add_79_4_n58 ), .ZN(sha1_round_wire[136]) );
NAND2_X2 _sha1_round_add_79_4_U253  ( .A1(_sha1_round_add_79_4_n55 ), .A2(_sha1_round_add_79_4_n311 ), .ZN(_sha1_round_add_79_4_n53 ) );
XNOR2_X2 _sha1_round_add_79_4_U252  ( .A(_sha1_round_add_79_4_n53 ), .B(_sha1_round_add_79_4_n54 ), .ZN(sha1_round_wire[137]) );
NAND2_X4 _sha1_round_add_79_4_U251  ( .A1(_sha1_round_add_79_4_n251 ), .A2(_sha1_round_add_79_4_n252 ), .ZN(_sha1_round_add_79_4_n236 ) );
NAND2_X1 _sha1_round_add_79_4_U250  ( .A1(_sha1_round_N333 ), .A2(rnd_q[140]), .ZN(_sha1_round_add_79_4_n260 ) );
NOR2_X1 _sha1_round_add_79_4_U249  ( .A1(_sha1_round_add_79_4_n250 ), .A2(_sha1_round_add_79_4_n236 ), .ZN(_sha1_round_add_79_4_n245 ) );
NAND2_X4 _sha1_round_add_79_4_U248  ( .A1(_sha1_round_add_79_4_n263 ), .A2(_sha1_round_add_79_4_n264 ), .ZN(_sha1_round_add_79_4_n252 ) );
NAND2_X4 _sha1_round_add_79_4_U247  ( .A1(_sha1_round_add_79_4_n163 ), .A2(_sha1_round_add_79_4_n164 ), .ZN(_sha1_round_add_79_4_n111 ) );
NAND3_X4 _sha1_round_add_79_4_U246  ( .A1(_sha1_round_add_79_4_n252 ), .A2(_sha1_round_n509 ), .A3(rnd_q[139]), .ZN(_sha1_round_add_79_4_n259 ));
NOR3_X2 _sha1_round_add_79_4_U245  ( .A1(_sha1_round_add_79_4_n147 ), .A2(_sha1_round_add_79_4_n148 ), .A3(_sha1_round_add_79_4_n100 ), .ZN(_sha1_round_add_79_4_n196 ) );
NOR3_X2 _sha1_round_add_79_4_U244  ( .A1(_sha1_round_add_79_4_n272 ), .A2(_sha1_round_add_79_4_n240 ), .A3(_sha1_round_add_79_4_n148 ), .ZN(_sha1_round_add_79_4_n267 ) );
NAND2_X1 _sha1_round_add_79_4_U243  ( .A1(_sha1_round_add_79_4_n307 ), .A2(_sha1_round_add_79_4_n303 ), .ZN(_sha1_round_add_79_4_n320 ) );
NAND2_X4 _sha1_round_add_79_4_U242  ( .A1(_sha1_round_add_79_4_n194 ), .A2(_sha1_round_add_79_4_n195 ), .ZN(_sha1_round_add_79_4_n165 ) );
NAND2_X1 _sha1_round_add_79_4_U241  ( .A1(_sha1_round_N343 ), .A2(rnd_q[150]), .ZN(_sha1_round_add_79_4_n164 ) );
NAND2_X4 _sha1_round_add_79_4_U240  ( .A1(_sha1_round_add_79_4_n168 ), .A2(_sha1_round_add_79_4_n169 ), .ZN(_sha1_round_add_79_4_n157 ) );
NAND2_X1 _sha1_round_add_79_4_U239  ( .A1(_sha1_round_add_79_4_n164 ), .A2(_sha1_round_add_79_4_n157 ), .ZN(_sha1_round_add_79_4_n167 ) );
NAND2_X1 _sha1_round_add_79_4_U238  ( .A1(_sha1_round_N346 ), .A2(rnd_q[153]), .ZN(_sha1_round_add_79_4_n116 ) );
NAND2_X1 _sha1_round_add_79_4_U237  ( .A1(_sha1_round_N344 ), .A2(rnd_q[151]), .ZN(_sha1_round_add_79_4_n131 ) );
NAND2_X1 _sha1_round_add_79_4_U236  ( .A1(rnd_q[144]), .A2(_sha1_round_N337 ), .ZN(_sha1_round_add_79_4_n204 ) );
INV_X1 _sha1_round_add_79_4_U235  ( .A(_sha1_round_add_79_4_n252 ), .ZN(_sha1_round_add_79_4_n261 ) );
NAND2_X1 _sha1_round_add_79_4_U234  ( .A1(_sha1_round_add_79_4_n117 ), .A2(_sha1_round_add_79_4_n127 ), .ZN(_sha1_round_add_79_4_n142 ) );
NAND2_X1 _sha1_round_add_79_4_U233  ( .A1(_sha1_round_add_79_4_n136 ), .A2(_sha1_round_add_79_4_n127 ), .ZN(_sha1_round_add_79_4_n135 ) );
NAND2_X1 _sha1_round_add_79_4_U232  ( .A1(_sha1_round_N334 ), .A2(rnd_q[141]), .ZN(_sha1_round_add_79_4_n247 ) );
NAND2_X1 _sha1_round_add_79_4_U231  ( .A1(_sha1_round_add_79_4_n131 ), .A2(_sha1_round_add_79_4_n158 ), .ZN(_sha1_round_add_79_4_n160 ) );
NAND2_X4 _sha1_round_add_79_4_U230  ( .A1(_sha1_round_add_79_4_n188 ), .A2(_sha1_round_add_79_4_n189 ), .ZN(_sha1_round_add_79_4_n179 ) );
NAND2_X1 _sha1_round_add_79_4_U229  ( .A1(_sha1_round_add_79_4_n179 ), .A2(_sha1_round_add_79_4_n184 ), .ZN(_sha1_round_add_79_4_n187 ) );
NOR2_X1 _sha1_round_add_79_4_U228  ( .A1(_sha1_round_add_79_4_n254 ), .A2(_sha1_round_add_79_4_n52 ), .ZN(_sha1_round_add_79_4_n266 ) );
NOR2_X1 _sha1_round_add_79_4_U227  ( .A1(_sha1_round_add_79_4_n254 ), .A2(_sha1_round_add_79_4_n250 ), .ZN(_sha1_round_add_79_4_n265 ) );
NOR3_X1 _sha1_round_add_79_4_U226  ( .A1(_sha1_round_add_79_4_n250 ), .A2(_sha1_round_add_79_4_n261 ), .A3(_sha1_round_add_79_4_n254 ), .ZN(_sha1_round_add_79_4_n258 ) );
NAND3_X2 _sha1_round_add_79_4_U225  ( .A1(_sha1_round_add_79_4_n95 ), .A2(_sha1_round_add_79_4_n146 ), .A3(_sha1_round_add_79_4_n145 ), .ZN(_sha1_round_add_79_4_n94 ) );
INV_X4 _sha1_round_add_79_4_U224  ( .A(_sha1_round_add_79_4_n273 ), .ZN(_sha1_round_add_79_4_n281 ) );
NAND2_X2 _sha1_round_add_79_4_U223  ( .A1(_sha1_round_add_79_4_n86 ), .A2(_sha1_round_add_79_4_n331 ), .ZN(_sha1_round_add_79_4_n81 ) );
AND2_X2 _sha1_round_add_79_4_U222  ( .A1(_sha1_round_n509 ), .A2(rnd_q[139]),.ZN(_sha1_round_add_79_4_n52 ) );
AND2_X2 _sha1_round_add_79_4_U221  ( .A1(_sha1_round_N336 ), .A2(rnd_q[143]),.ZN(_sha1_round_add_79_4_n51 ) );
NOR2_X2 _sha1_round_add_79_4_U220  ( .A1(_sha1_round_add_79_4_n344 ), .A2(_sha1_round_add_79_4_n345 ), .ZN(_sha1_round_add_79_4_n343 ) );
NAND3_X1 _sha1_round_add_79_4_U219  ( .A1(rnd_q[128]), .A2(_sha1_round_N321 ), .A3(_sha1_round_add_79_4_n72 ), .ZN(_sha1_round_add_79_4_n342 ) );
NAND3_X2 _sha1_round_add_79_4_U218  ( .A1(_sha1_round_add_79_4_n341 ), .A2(_sha1_round_add_79_4_n342 ), .A3(_sha1_round_add_79_4_n343 ), .ZN(_sha1_round_add_79_4_n316 ) );
OR2_X2 _sha1_round_add_79_4_U217  ( .A1(rnd_q[155]), .A2(_sha1_round_N316 ),.ZN(_sha1_round_add_79_4_n50 ) );
OR2_X2 _sha1_round_add_79_4_U216  ( .A1(_sha1_round_N318 ), .A2(rnd_q[157]),.ZN(_sha1_round_add_79_4_n90 ) );
NOR2_X2 _sha1_round_add_79_4_U215  ( .A1(rnd_q[159]), .A2(_sha1_round_N320 ),.ZN(_sha1_round_add_79_4_n80 ) );
NOR2_X2 _sha1_round_add_79_4_U214  ( .A1(rnd_q[156]), .A2(_sha1_round_N317 ),.ZN(_sha1_round_add_79_4_n140 ) );
NOR2_X2 _sha1_round_add_79_4_U213  ( .A1(rnd_q[128]), .A2(_sha1_round_N321 ),.ZN(_sha1_round_add_79_4_n75 ) );
OR2_X2 _sha1_round_add_79_4_U212  ( .A1(_sha1_round_N319 ), .A2(rnd_q[158]),.ZN(_sha1_round_add_79_4_n85 ) );
AND2_X2 _sha1_round_add_79_4_U211  ( .A1(_sha1_round_add_79_4_n203 ), .A2(_sha1_round_add_79_4_n201 ), .ZN(_sha1_round_add_79_4_n46 ) );
AND2_X2 _sha1_round_add_79_4_U210  ( .A1(_sha1_round_add_79_4_n271 ), .A2(_sha1_round_add_79_4_n298 ), .ZN(_sha1_round_add_79_4_n45 ) );
NOR2_X1 _sha1_round_add_79_4_U209  ( .A1(_sha1_round_add_79_4_n112 ), .A2(_sha1_round_add_79_4_n120 ), .ZN(_sha1_round_add_79_4_n119 ) );
NOR2_X1 _sha1_round_add_79_4_U208  ( .A1(_sha1_round_add_79_4_n269 ), .A2(_sha1_round_add_79_4_n5 ), .ZN(_sha1_round_add_79_4_n287 ) );
NOR2_X1 _sha1_round_add_79_4_U207  ( .A1(_sha1_round_add_79_4_n3 ), .A2(_sha1_round_add_79_4_n49 ), .ZN(_sha1_round_add_79_4_n292 ) );
NOR2_X1 _sha1_round_add_79_4_U206  ( .A1(_sha1_round_add_79_4_n48 ), .A2(_sha1_round_add_79_4_n297 ), .ZN(_sha1_round_add_79_4_n300 ) );
NOR2_X2 _sha1_round_add_79_4_U205  ( .A1(_sha1_round_add_79_4_n275 ), .A2(_sha1_round_add_79_4_n300 ), .ZN(_sha1_round_add_79_4_n299 ) );
NOR2_X1 _sha1_round_add_79_4_U204  ( .A1(_sha1_round_add_79_4_n275 ), .A2(_sha1_round_add_79_4_n48 ), .ZN(_sha1_round_add_79_4_n301 ) );
NOR2_X2 _sha1_round_add_79_4_U203  ( .A1(_sha1_round_add_79_4_n59 ), .A2(_sha1_round_add_79_4_n60 ), .ZN(_sha1_round_add_79_4_n58 ) );
NOR2_X2 _sha1_round_add_79_4_U202  ( .A1(_sha1_round_add_79_4_n265 ), .A2(_sha1_round_add_79_4_n52 ), .ZN(_sha1_round_add_79_4_n262 ) );
NOR2_X1 _sha1_round_add_79_4_U201  ( .A1(_sha1_round_add_79_4_n218 ), .A2(_sha1_round_add_79_4_n51 ), .ZN(_sha1_round_add_79_4_n230 ) );
NOR2_X2 _sha1_round_add_79_4_U200  ( .A1(_sha1_round_add_79_4_n242 ), .A2(_sha1_round_add_79_4_n140 ), .ZN(_sha1_round_add_79_4_n241 ) );
NOR2_X2 _sha1_round_add_79_4_U199  ( .A1(_sha1_round_add_79_4_n335 ), .A2(_sha1_round_add_79_4_n140 ), .ZN(_sha1_round_add_79_4_n334 ) );
NAND3_X1 _sha1_round_add_79_4_U198  ( .A1(_sha1_round_add_79_4_n318 ), .A2(_sha1_round_add_79_4_n314 ), .A3(_sha1_round_add_79_4_n81 ), .ZN(_sha1_round_add_79_4_n330 ) );
NAND3_X2 _sha1_round_add_79_4_U197  ( .A1(_sha1_round_add_79_4_n312 ), .A2(_sha1_round_add_79_4_n329 ), .A3(_sha1_round_add_79_4_n330 ), .ZN(_sha1_round_add_79_4_n54 ) );
NOR2_X1 _sha1_round_add_79_4_U196  ( .A1(_sha1_round_add_79_4_n253 ), .A2(_sha1_round_add_79_4_n257 ), .ZN(_sha1_round_add_79_4_n256 ) );
NOR3_X2 _sha1_round_add_79_4_U195  ( .A1(_sha1_round_add_79_4_n7 ), .A2(_sha1_round_add_79_4_n284 ), .A3(_sha1_round_add_79_4_n285 ), .ZN(_sha1_round_add_79_4_n283 ) );
AND2_X2 _sha1_round_add_79_4_U194  ( .A1(_sha1_round_add_79_4_n43 ), .A2(_sha1_round_add_79_4_n79 ), .ZN(_sha1_round_add_79_4_n76 ) );
OR2_X2 _sha1_round_add_79_4_U193  ( .A1(_sha1_round_add_79_4_n140 ), .A2(_sha1_round_add_79_4_n243 ), .ZN(_sha1_round_add_79_4_n42 ) );
NOR2_X2 _sha1_round_add_79_4_U192  ( .A1(_sha1_round_add_79_4_n332 ), .A2(_sha1_round_add_79_4_n87 ), .ZN(_sha1_round_add_79_4_n285 ) );
NOR2_X1 _sha1_round_add_79_4_U191  ( .A1(_sha1_round_add_79_4_n278 ), .A2(_sha1_round_add_79_4_n296 ), .ZN(_sha1_round_add_79_4_n295 ) );
AND2_X2 _sha1_round_add_79_4_U190  ( .A1(_sha1_round_add_79_4_n204 ), .A2(_sha1_round_add_79_4_n225 ), .ZN(_sha1_round_add_79_4_n40 ) );
AND2_X2 _sha1_round_add_79_4_U189  ( .A1(_sha1_round_add_79_4_n260 ), .A2(_sha1_round_add_79_4_n252 ), .ZN(_sha1_round_add_79_4_n39 ) );
AND2_X2 _sha1_round_add_79_4_U188  ( .A1(_sha1_round_add_79_4_n150 ), .A2(_sha1_round_add_79_4_n210 ), .ZN(_sha1_round_add_79_4_n38 ) );
NOR2_X2 _sha1_round_add_79_4_U187  ( .A1(_sha1_round_add_79_4_n49 ), .A2(_sha1_round_add_79_4_n271 ), .ZN(_sha1_round_add_79_4_n270 ) );
NOR2_X2 _sha1_round_add_79_4_U186  ( .A1(_sha1_round_add_79_4_n7 ), .A2(_sha1_round_add_79_4_n285 ), .ZN(_sha1_round_add_79_4_n331 ) );
NOR2_X1 _sha1_round_add_79_4_U185  ( .A1(_sha1_round_add_79_4_n61 ), .A2(_sha1_round_add_79_4_n62 ), .ZN(_sha1_round_add_79_4_n57 ) );
NOR2_X2 _sha1_round_add_79_4_U184  ( .A1(_sha1_round_add_79_4_n27 ), .A2(_sha1_round_add_79_4_n151 ), .ZN(_sha1_round_add_79_4_n143 ) );
NOR2_X1 _sha1_round_add_79_4_U183  ( .A1(_sha1_round_add_79_4_n269 ), .A2(_sha1_round_add_79_4_n235 ), .ZN(_sha1_round_add_79_4_n268 ) );
OR2_X4 _sha1_round_add_79_4_U182  ( .A1(_sha1_round_N329 ), .A2(rnd_q[136]),.ZN(_sha1_round_add_79_4_n298 ) );
OR2_X4 _sha1_round_add_79_4_U181  ( .A1(_sha1_round_N345 ), .A2(rnd_q[152]),.ZN(_sha1_round_add_79_4_n127 ) );
OR2_X4 _sha1_round_add_79_4_U180  ( .A1(_sha1_round_N322 ), .A2(rnd_q[129]),.ZN(_sha1_round_add_79_4_n72 ) );
OR2_X1 _sha1_round_add_79_4_U179  ( .A1(_sha1_round_add_79_4_n63 ), .A2(_sha1_round_add_79_4_n80 ), .ZN(_sha1_round_add_79_4_n43 ) );
NOR2_X1 _sha1_round_add_79_4_U178  ( .A1(_sha1_round_add_79_4_n78 ), .A2(_sha1_round_add_79_4_n75 ), .ZN(_sha1_round_add_79_4_n77 ) );
OR2_X4 _sha1_round_add_79_4_U177  ( .A1(_sha1_round_add_79_4_n75 ), .A2(_sha1_round_add_79_4_n76 ), .ZN(_sha1_round_add_79_4_n41 ) );
AND2_X2 _sha1_round_add_79_4_U176  ( .A1(_sha1_round_add_79_4_n302 ), .A2(_sha1_round_add_79_4_n281 ), .ZN(_sha1_round_add_79_4_n37 ) );
NAND3_X4 _sha1_round_add_79_4_U175  ( .A1(_sha1_round_add_79_4_n279 ), .A2(_sha1_round_add_79_4_n280 ), .A3(_sha1_round_add_79_4_n281 ), .ZN(_sha1_round_add_79_4_n149 ) );
NOR2_X1 _sha1_round_add_79_4_U174  ( .A1(_sha1_round_add_79_4_n63 ), .A2(_sha1_round_add_79_4_n64 ), .ZN(_sha1_round_add_79_4_n61 ) );
OR2_X4 _sha1_round_add_79_4_U173  ( .A1(_sha1_round_N338 ), .A2(rnd_q[145]),.ZN(_sha1_round_add_79_4_n203 ) );
OR2_X4 _sha1_round_add_79_4_U172  ( .A1(_sha1_round_N339 ), .A2(rnd_q[146]),.ZN(_sha1_round_add_79_4_n154 ) );
NOR2_X2 _sha1_round_add_79_4_U171  ( .A1(_sha1_round_add_79_4_n245 ), .A2(_sha1_round_add_79_4_n209 ), .ZN(_sha1_round_add_79_4_n244 ) );
AND2_X4 _sha1_round_add_79_4_U170  ( .A1(_sha1_round_add_79_4_n21 ), .A2(_sha1_round_add_79_4_n150 ), .ZN(_sha1_round_add_79_4_n44 ) );
NOR2_X2 _sha1_round_add_79_4_U169  ( .A1(_sha1_round_add_79_4_n134 ), .A2(_sha1_round_add_79_4_n9 ), .ZN(_sha1_round_add_79_4_n121 ) );
NOR2_X2 _sha1_round_add_79_4_U168  ( .A1(rnd_q[131]), .A2(_sha1_round_N324 ),.ZN(_sha1_round_add_79_4_n60 ) );
NAND2_X2 _sha1_round_add_79_4_U167  ( .A1(_sha1_round_add_79_4_n21 ), .A2(_sha1_round_add_79_4_n150 ), .ZN(_sha1_round_add_79_4_n208 ) );
NOR2_X1 _sha1_round_add_79_4_U166  ( .A1(_sha1_round_add_79_4_n99 ), .A2(_sha1_round_add_79_4_n137 ), .ZN(_sha1_round_add_79_4_n134 ) );
NAND2_X2 _sha1_round_add_79_4_U165  ( .A1(_sha1_round_add_79_4_n208 ), .A2(_sha1_round_add_79_4_n136 ), .ZN(_sha1_round_add_79_4_n207 ) );
XNOR2_X1 _sha1_round_add_79_4_U164  ( .A(_sha1_round_add_79_4_n291 ), .B(_sha1_round_add_79_4_n292 ), .ZN(sha1_round_wire[142]) );
INV_X1 _sha1_round_add_79_4_U163  ( .A(_sha1_round_add_79_4_n271 ), .ZN(_sha1_round_add_79_4_n294 ) );
NOR2_X4 _sha1_round_add_79_4_U162  ( .A1(_sha1_round_add_79_4_n273 ), .A2(_sha1_round_add_79_4_n11 ), .ZN(_sha1_round_add_79_4_n148 ) );
NAND2_X4 _sha1_round_add_79_4_U161  ( .A1(_sha1_round_add_79_4_n156 ), .A2(_sha1_round_add_79_4_n110 ), .ZN(_sha1_round_add_79_4_n96 ) );
NOR2_X4 _sha1_round_add_79_4_U160  ( .A1(_sha1_round_add_79_4_n129 ), .A2(_sha1_round_add_79_4_n130 ), .ZN(_sha1_round_add_79_4_n106 ) );
NOR2_X2 _sha1_round_add_79_4_U159  ( .A1(_sha1_round_add_79_4_n106 ), .A2(_sha1_round_add_79_4_n107 ), .ZN(_sha1_round_add_79_4_n103 ) );
NAND2_X4 _sha1_round_add_79_4_U158  ( .A1(_sha1_round_add_79_4_n158 ), .A2(_sha1_round_add_79_4_n157 ), .ZN(_sha1_round_add_79_4_n36 ) );
INV_X4 _sha1_round_add_79_4_U157  ( .A(_sha1_round_add_79_4_n96 ), .ZN(_sha1_round_add_79_4_n145 ) );
NAND2_X2 _sha1_round_add_79_4_U156  ( .A1(_sha1_round_add_79_4_n2 ), .A2(_sha1_round_add_79_4_n146 ), .ZN(_sha1_round_add_79_4_n144 ) );
INV_X4 _sha1_round_add_79_4_U155  ( .A(_sha1_round_add_79_4_n92 ), .ZN(_sha1_round_add_79_4_n33 ) );
NAND2_X2 _sha1_round_add_79_4_U154  ( .A1(_sha1_round_add_79_4_n91 ), .A2(_sha1_round_add_79_4_n92 ), .ZN(_sha1_round_add_79_4_n34 ) );
NAND2_X2 _sha1_round_add_79_4_U153  ( .A1(_sha1_round_add_79_4_n17 ), .A2(_sha1_round_add_79_4_n165 ), .ZN(_sha1_round_add_79_4_n182 ) );
NAND2_X2 _sha1_round_add_79_4_U152  ( .A1(_sha1_round_add_79_4_n156 ), .A2(_sha1_round_add_79_4_n165 ), .ZN(_sha1_round_add_79_4_n170 ) );
NAND2_X2 _sha1_round_add_79_4_U151  ( .A1(_sha1_round_add_79_4_n178 ), .A2(_sha1_round_add_79_4_n165 ), .ZN(_sha1_round_add_79_4_n190 ) );
NAND3_X4 _sha1_round_add_79_4_U150  ( .A1(_sha1_round_add_79_4_n215 ), .A2(_sha1_round_add_79_4_n201 ), .A3(_sha1_round_add_79_4_n6 ), .ZN(_sha1_round_add_79_4_n213 ) );
NAND2_X2 _sha1_round_add_79_4_U149  ( .A1(_sha1_round_add_79_4_n1 ), .A2(_sha1_round_add_79_4_n165 ), .ZN(_sha1_round_add_79_4_n161 ) );
NAND3_X1 _sha1_round_add_79_4_U148  ( .A1(_sha1_round_add_79_4_n68 ), .A2(_sha1_round_add_79_4_n316 ), .A3(_sha1_round_add_79_4_n274 ), .ZN(_sha1_round_add_79_4_n315 ) );
NAND3_X1 _sha1_round_add_79_4_U147  ( .A1(_sha1_round_add_79_4_n314 ), .A2(_sha1_round_add_79_4_n274 ), .A3(_sha1_round_add_79_4_n81 ), .ZN(_sha1_round_add_79_4_n302 ) );
NAND3_X4 _sha1_round_add_79_4_U146  ( .A1(_sha1_round_add_79_4_n153 ), .A2(_sha1_round_add_79_4_n145 ), .A3(_sha1_round_add_79_4_n154 ), .ZN(_sha1_round_add_79_4_n105 ) );
NAND2_X2 _sha1_round_add_79_4_U145  ( .A1(_sha1_round_add_79_4_n183 ), .A2(_sha1_round_add_79_4_n179 ), .ZN(_sha1_round_add_79_4_n173 ) );
INV_X1 _sha1_round_add_79_4_U144  ( .A(_sha1_round_add_79_4_n176 ), .ZN(_sha1_round_add_79_4_n172 ) );
NOR2_X4 _sha1_round_add_79_4_U143  ( .A1(_sha1_round_add_79_4_n112 ), .A2(_sha1_round_add_79_4_n113 ), .ZN(_sha1_round_add_79_4_n101 ) );
NAND3_X2 _sha1_round_add_79_4_U142  ( .A1(_sha1_round_add_79_4_n152 ), .A2(_sha1_round_add_79_4_n105 ), .A3(_sha1_round_add_79_4_n131 ), .ZN(_sha1_round_add_79_4_n151 ) );
NAND2_X2 _sha1_round_add_79_4_U141  ( .A1(_sha1_round_add_79_4_n182 ), .A2(_sha1_round_add_79_4_n173 ), .ZN(_sha1_round_add_79_4_n180 ) );
INV_X2 _sha1_round_add_79_4_U140  ( .A(_sha1_round_add_79_4_n253 ), .ZN(_sha1_round_add_79_4_n249 ) );
NAND2_X4 _sha1_round_add_79_4_U139  ( .A1(_sha1_round_add_79_4_n128 ), .A2(_sha1_round_add_79_4_n127 ), .ZN(_sha1_round_add_79_4_n124 ) );
NOR2_X4 _sha1_round_add_79_4_U138  ( .A1(rnd_q[141]), .A2(_sha1_round_N334 ),.ZN(_sha1_round_add_79_4_n253 ) );
NAND2_X4 _sha1_round_add_79_4_U137  ( .A1(_sha1_round_add_79_4_n93 ), .A2(_sha1_round_add_79_4_n94 ), .ZN(_sha1_round_add_79_4_n91 ) );
NOR2_X2 _sha1_round_add_79_4_U136  ( .A1(_sha1_round_add_79_4_n107 ), .A2(_sha1_round_add_79_4_n100 ), .ZN(_sha1_round_add_79_4_n95 ) );
NAND2_X2 _sha1_round_add_79_4_U135  ( .A1(_sha1_round_add_79_4_n126 ), .A2(_sha1_round_add_79_4_n127 ), .ZN(_sha1_round_add_79_4_n125 ) );
AND2_X4 _sha1_round_add_79_4_U134  ( .A1(_sha1_round_add_79_4_n132 ), .A2(_sha1_round_add_79_4_n117 ), .ZN(_sha1_round_add_79_4_n123 ) );
NOR2_X1 _sha1_round_add_79_4_U133  ( .A1(_sha1_round_add_79_4_n218 ), .A2(_sha1_round_add_79_4_n216 ), .ZN(_sha1_round_add_79_4_n229 ) );
NAND2_X4 _sha1_round_add_79_4_U132  ( .A1(_sha1_round_add_79_4_n15 ), .A2(_sha1_round_add_79_4_n238 ), .ZN(_sha1_round_add_79_4_n147 ) );
NOR2_X1 _sha1_round_add_79_4_U131  ( .A1(_sha1_round_add_79_4_n216 ), .A2(_sha1_round_add_79_4_n14 ), .ZN(_sha1_round_add_79_4_n222 ) );
INV_X4 _sha1_round_add_79_4_U130  ( .A(_sha1_round_add_79_4_n214 ), .ZN(_sha1_round_add_79_4_n29 ) );
NAND2_X2 _sha1_round_add_79_4_U129  ( .A1(_sha1_round_add_79_4_n213 ), .A2(_sha1_round_add_79_4_n214 ), .ZN(_sha1_round_add_79_4_n30 ) );
OR2_X4 _sha1_round_add_79_4_U128  ( .A1(_sha1_round_N323 ), .A2(rnd_q[130]),.ZN(_sha1_round_add_79_4_n68 ) );
AND2_X4 _sha1_round_add_79_4_U127  ( .A1(_sha1_round_add_79_4_n315 ), .A2(_sha1_round_add_79_4_n37 ), .ZN(_sha1_round_add_79_4_n297 ) );
NAND2_X2 _sha1_round_add_79_4_U126  ( .A1(_sha1_round_add_79_4_n27 ), .A2(_sha1_round_add_79_4_n101 ), .ZN(_sha1_round_add_79_4_n109 ) );
NAND2_X2 _sha1_round_add_79_4_U125  ( .A1(_sha1_round_add_79_4_n111 ), .A2(_sha1_round_add_79_4_n20 ), .ZN(_sha1_round_add_79_4_n26 ) );
INV_X2 _sha1_round_add_79_4_U124  ( .A(_sha1_round_add_79_4_n142 ), .ZN(_sha1_round_add_79_4_n23 ) );
INV_X4 _sha1_round_add_79_4_U123  ( .A(_sha1_round_add_79_4_n141 ), .ZN(_sha1_round_add_79_4_n22 ) );
NAND2_X4 _sha1_round_add_79_4_U122  ( .A1(_sha1_round_add_79_4_n276 ), .A2(_sha1_round_add_79_4_n277 ), .ZN(_sha1_round_add_79_4_n240 ) );
NAND2_X2 _sha1_round_add_79_4_U121  ( .A1(_sha1_round_add_79_4_n133 ), .A2(_sha1_round_add_79_4_n111 ), .ZN(_sha1_round_add_79_4_n132 ) );
NOR2_X4 _sha1_round_add_79_4_U120  ( .A1(_sha1_round_add_79_4_n235 ), .A2(_sha1_round_add_79_4_n236 ), .ZN(_sha1_round_add_79_4_n234 ) );
NAND2_X4 _sha1_round_add_79_4_U119  ( .A1(_sha1_round_add_79_4_n4 ), .A2(_sha1_round_add_79_4_n234 ), .ZN(_sha1_round_add_79_4_n21 ) );
NOR3_X4 _sha1_round_add_79_4_U118  ( .A1(_sha1_round_add_79_4_n270 ), .A2(_sha1_round_add_79_4_n3 ), .A3(_sha1_round_add_79_4_n5 ), .ZN(_sha1_round_add_79_4_n235 ) );
NAND2_X2 _sha1_round_add_79_4_U117  ( .A1(_sha1_round_add_79_4_n306 ), .A2(_sha1_round_add_79_4_n307 ), .ZN(_sha1_round_add_79_4_n305 ) );
NOR2_X2 _sha1_round_add_79_4_U116  ( .A1(_sha1_round_add_79_4_n258 ), .A2(_sha1_round_add_79_4_n248 ), .ZN(_sha1_round_add_79_4_n255 ) );
INV_X2 _sha1_round_add_79_4_U115  ( .A(_sha1_round_add_79_4_n149 ), .ZN(_sha1_round_add_79_4_n237 ) );
NAND2_X1 _sha1_round_add_79_4_U114  ( .A1(_sha1_round_N327 ), .A2(rnd_q[134]), .ZN(_sha1_round_add_79_4_n303 ) );
NAND3_X2 _sha1_round_add_79_4_U113  ( .A1(_sha1_round_add_79_4_n44 ), .A2(_sha1_round_add_79_4_n97 ), .A3(_sha1_round_add_79_4_n98 ), .ZN(_sha1_round_add_79_4_n146 ) );
INV_X2 _sha1_round_add_79_4_U112  ( .A(_sha1_round_add_79_4_n19 ), .ZN(_sha1_round_add_79_4_n20 ) );
INV_X1 _sha1_round_add_79_4_U111  ( .A(_sha1_round_add_79_4_n110 ), .ZN(_sha1_round_add_79_4_n19 ) );
XNOR2_X1 _sha1_round_add_79_4_U110  ( .A(_sha1_round_add_79_4_n216 ), .B(_sha1_round_add_79_4_n230 ), .ZN(sha1_round_wire[148]) );
NOR2_X2 _sha1_round_add_79_4_U109  ( .A1(_sha1_round_add_79_4_n283 ), .A2(_sha1_round_add_79_4_n64 ), .ZN(_sha1_round_add_79_4_n282 ) );
NOR2_X4 _sha1_round_add_79_4_U108  ( .A1(_sha1_round_add_79_4_n282 ), .A2(_sha1_round_add_79_4_n275 ), .ZN(_sha1_round_add_79_4_n279 ) );
INV_X4 _sha1_round_add_79_4_U107  ( .A(_sha1_round_add_79_4_n236 ), .ZN(_sha1_round_add_79_4_n239 ) );
NAND2_X1 _sha1_round_add_79_4_U106  ( .A1(_sha1_round_add_79_4_n114 ), .A2(_sha1_round_add_79_4_n115 ), .ZN(_sha1_round_add_79_4_n108 ) );
INV_X2 _sha1_round_add_79_4_U105  ( .A(_sha1_round_add_79_4_n47 ), .ZN(_sha1_round_add_79_4_n210 ) );
INV_X2 _sha1_round_add_79_4_U104  ( .A(_sha1_round_add_79_4_n26 ), .ZN(_sha1_round_add_79_4_n27 ) );
OR2_X2 _sha1_round_add_79_4_U103  ( .A1(_sha1_round_N346 ), .A2(rnd_q[153]),.ZN(_sha1_round_add_79_4_n115 ) );
INV_X4 _sha1_round_add_79_4_U102  ( .A(_sha1_round_add_79_4_n115 ), .ZN(_sha1_round_add_79_4_n112 ) );
NOR2_X4 _sha1_round_add_79_4_U101  ( .A1(rnd_q[149]), .A2(_sha1_round_N342 ),.ZN(_sha1_round_add_79_4_n176 ) );
NAND2_X2 _sha1_round_add_79_4_U100  ( .A1(_sha1_round_N323 ), .A2(rnd_q[130]), .ZN(_sha1_round_add_79_4_n67 ) );
NOR2_X2 _sha1_round_add_79_4_U99  ( .A1(_sha1_round_add_79_4_n229 ), .A2(_sha1_round_add_79_4_n51 ), .ZN(_sha1_round_add_79_4_n226 ) );
NOR2_X2 _sha1_round_add_79_4_U98  ( .A1(_sha1_round_add_79_4_n197 ), .A2(_sha1_round_add_79_4_n198 ), .ZN(_sha1_round_add_79_4_n194 ) );
AND2_X4 _sha1_round_add_79_4_U97  ( .A1(_sha1_round_add_79_4_n318 ), .A2(_sha1_round_add_79_4_n313 ), .ZN(_sha1_round_add_79_4_n18 ) );
INV_X4 _sha1_round_add_79_4_U96  ( .A(_sha1_round_add_79_4_n205 ), .ZN(_sha1_round_add_79_4_n220 ) );
AND2_X4 _sha1_round_add_79_4_U95  ( .A1(_sha1_round_add_79_4_n178 ), .A2(_sha1_round_add_79_4_n179 ), .ZN(_sha1_round_add_79_4_n17 ) );
AND2_X4 _sha1_round_add_79_4_U94  ( .A1(_sha1_round_add_79_4_n243 ), .A2(_sha1_round_add_79_4_n50 ), .ZN(sha1_round_wire[128]) );
NOR2_X2 _sha1_round_add_79_4_U93  ( .A1(rnd_q[132]), .A2(_sha1_round_N325 ),.ZN(_sha1_round_add_79_4_n56 ) );
AND2_X2 _sha1_round_add_79_4_U92  ( .A1(_sha1_round_add_79_4_n239 ), .A2(_sha1_round_add_79_4_n210 ), .ZN(_sha1_round_add_79_4_n15 ) );
OR2_X4 _sha1_round_add_79_4_U91  ( .A1(_sha1_round_add_79_4_n219 ), .A2(_sha1_round_add_79_4_n218 ), .ZN(_sha1_round_add_79_4_n14 ) );
AND2_X4 _sha1_round_add_79_4_U90  ( .A1(_sha1_round_add_79_4_n150 ), .A2(_sha1_round_add_79_4_n21 ), .ZN(_sha1_round_add_79_4_n13 ) );
AND2_X4 _sha1_round_add_79_4_U89  ( .A1(_sha1_round_add_79_4_n303 ), .A2(_sha1_round_add_79_4_n305 ), .ZN(_sha1_round_add_79_4_n12 ) );
OR2_X4 _sha1_round_add_79_4_U88  ( .A1(_sha1_round_add_79_4_n274 ), .A2(_sha1_round_add_79_4_n275 ), .ZN(_sha1_round_add_79_4_n11 ) );
OR2_X4 _sha1_round_add_79_4_U87  ( .A1(_sha1_round_add_79_4_n295 ), .A2(_sha1_round_add_79_4_n294 ), .ZN(_sha1_round_add_79_4_n10 ) );
OR2_X1 _sha1_round_add_79_4_U86  ( .A1(_sha1_round_add_79_4_n135 ), .A2(_sha1_round_add_79_4_n96 ), .ZN(_sha1_round_add_79_4_n9 ) );
OR2_X4 _sha1_round_add_79_4_U85  ( .A1(_sha1_round_add_79_4_n278 ), .A2(_sha1_round_add_79_4_n48 ), .ZN(_sha1_round_add_79_4_n8 ) );
AND3_X4 _sha1_round_add_79_4_U84  ( .A1(_sha1_round_add_79_4_n85 ), .A2(_sha1_round_add_79_4_n333 ), .A3(_sha1_round_add_79_4_n334 ), .ZN(_sha1_round_add_79_4_n7 ) );
OR2_X4 _sha1_round_add_79_4_U83  ( .A1(_sha1_round_add_79_4_n216 ), .A2(_sha1_round_add_79_4_n212 ), .ZN(_sha1_round_add_79_4_n6 ) );
AND2_X4 _sha1_round_add_79_4_U82  ( .A1(_sha1_round_add_79_4_n233 ), .A2(_sha1_round_add_79_4_n210 ), .ZN(_sha1_round_add_79_4_n4 ) );
AND2_X4 _sha1_round_add_79_4_U81  ( .A1(_sha1_round_N330 ), .A2(rnd_q[137]),.ZN(_sha1_round_add_79_4_n3 ) );
NOR3_X4 _sha1_round_add_79_4_U80  ( .A1(_sha1_round_add_79_4_n102 ), .A2(_sha1_round_add_79_4_n103 ), .A3(_sha1_round_add_79_4_n104 ), .ZN(_sha1_round_add_79_4_n93 ) );
NAND2_X1 _sha1_round_add_79_4_U79  ( .A1(_sha1_round_N345 ), .A2(rnd_q[152]),.ZN(_sha1_round_add_79_4_n117 ) );
INV_X2 _sha1_round_add_79_4_U78  ( .A(_sha1_round_N340 ), .ZN(_sha1_round_add_79_4_n192 ) );
NAND2_X1 _sha1_round_add_79_4_U77  ( .A1(_sha1_round_add_79_4_n111 ), .A2(_sha1_round_add_79_4_n157 ), .ZN(_sha1_round_add_79_4_n162 ) );
INV_X4 _sha1_round_add_79_4_U76  ( .A(_sha1_round_add_79_4_n101 ), .ZN(_sha1_round_add_79_4_n107 ) );
NAND2_X1 _sha1_round_add_79_4_U75  ( .A1(_sha1_round_N335 ), .A2(rnd_q[142]),.ZN(_sha1_round_add_79_4_n150 ) );
AND2_X2 _sha1_round_add_79_4_U74  ( .A1(_sha1_round_N331 ), .A2(rnd_q[138]),.ZN(_sha1_round_add_79_4_n5 ) );
INV_X4 _sha1_round_add_79_4_U73  ( .A(_sha1_round_add_79_4_n91 ), .ZN(_sha1_round_add_79_4_n32 ) );
NAND2_X2 _sha1_round_add_79_4_U72  ( .A1(_sha1_round_add_79_4_n24 ), .A2(_sha1_round_add_79_4_n25 ), .ZN(sha1_round_wire[157]) );
NOR3_X2 _sha1_round_add_79_4_U71  ( .A1(_sha1_round_add_79_4_n237 ), .A2(_sha1_round_add_79_4_n147 ), .A3(_sha1_round_add_79_4_n148 ), .ZN(_sha1_round_add_79_4_n231 ) );
NOR2_X2 _sha1_round_add_79_4_U70  ( .A1(_sha1_round_add_79_4_n49 ), .A2(_sha1_round_add_79_4_n291 ), .ZN(_sha1_round_add_79_4_n290 ) );
NOR2_X2 _sha1_round_add_79_4_U69  ( .A1(_sha1_round_add_79_4_n3 ), .A2(_sha1_round_add_79_4_n290 ), .ZN(_sha1_round_add_79_4_n286 ) );
INV_X4 _sha1_round_add_79_4_U68  ( .A(_sha1_round_add_79_4_n213 ), .ZN(_sha1_round_add_79_4_n28 ) );
NAND2_X2 _sha1_round_add_79_4_U67  ( .A1(_sha1_round_add_79_4_n32 ), .A2(_sha1_round_add_79_4_n33 ), .ZN(_sha1_round_add_79_4_n35 ) );
NAND2_X2 _sha1_round_add_79_4_U66  ( .A1(_sha1_round_add_79_4_n206 ), .A2(_sha1_round_add_79_4_n207 ), .ZN(_sha1_round_add_79_4_n197 ) );
NAND2_X2 _sha1_round_add_79_4_U65  ( .A1(_sha1_round_add_79_4_n227 ), .A2(_sha1_round_add_79_4_n228 ), .ZN(_sha1_round_add_79_4_n225 ) );
NOR2_X2 _sha1_round_add_79_4_U64  ( .A1(_sha1_round_N330 ), .A2(rnd_q[137]),.ZN(_sha1_round_add_79_4_n49 ) );
NOR2_X2 _sha1_round_add_79_4_U63  ( .A1(_sha1_round_add_79_4_n56 ), .A2(_sha1_round_add_79_4_n317 ), .ZN(_sha1_round_add_79_4_n274 ) );
INV_X4 _sha1_round_add_79_4_U62  ( .A(_sha1_round_add_79_4_n68 ), .ZN(_sha1_round_add_79_4_n340 ) );
NAND2_X2 _sha1_round_add_79_4_U61  ( .A1(_sha1_round_N341 ), .A2(rnd_q[148]),.ZN(_sha1_round_add_79_4_n184 ) );
NOR2_X2 _sha1_round_add_79_4_U60  ( .A1(_sha1_round_add_79_4_n219 ), .A2(_sha1_round_add_79_4_n224 ), .ZN(_sha1_round_add_79_4_n205 ) );
NOR2_X2 _sha1_round_add_79_4_U59  ( .A1(_sha1_round_add_79_4_n218 ), .A2(_sha1_round_add_79_4_n219 ), .ZN(_sha1_round_add_79_4_n217 ) );
NOR2_X2 _sha1_round_add_79_4_U58  ( .A1(_sha1_round_add_79_4_n107 ), .A2(_sha1_round_add_79_4_n105 ), .ZN(_sha1_round_add_79_4_n104 ) );
INV_X4 _sha1_round_add_79_4_U57  ( .A(_sha1_round_add_79_4_n127 ), .ZN(_sha1_round_add_79_4_n113 ) );
NOR2_X2 _sha1_round_add_79_4_U56  ( .A1(_sha1_round_add_79_4_n222 ), .A2(_sha1_round_add_79_4_n223 ), .ZN(_sha1_round_add_79_4_n221 ) );
NAND2_X2 _sha1_round_add_79_4_U55  ( .A1(_sha1_round_add_79_4_n22 ), .A2(_sha1_round_add_79_4_n23 ), .ZN(_sha1_round_add_79_4_n25 ) );
INV_X4 _sha1_round_add_79_4_U54  ( .A(_sha1_round_add_79_4_n240 ), .ZN(_sha1_round_add_79_4_n238 ) );
NOR2_X2 _sha1_round_add_79_4_U53  ( .A1(_sha1_round_N328 ), .A2(rnd_q[135]),.ZN(_sha1_round_add_79_4_n48 ) );
NAND2_X2 _sha1_round_add_79_4_U52  ( .A1(_sha1_round_add_79_4_n288 ), .A2(_sha1_round_add_79_4_n289 ), .ZN(_sha1_round_add_79_4_n233 ) );
INV_X4 _sha1_round_add_79_4_U51  ( .A(_sha1_round_add_79_4_n225 ), .ZN(_sha1_round_add_79_4_n219 ) );
XNOR2_X1 _sha1_round_add_79_4_U50  ( .A(_sha1_round_add_79_4_n266 ), .B(_sha1_round_add_79_4_n250 ), .ZN(sha1_round_wire[144]) );
NAND2_X1 _sha1_round_add_79_4_U49  ( .A1(_sha1_round_N324 ), .A2(rnd_q[131]),.ZN(_sha1_round_add_79_4_n312 ) );
OR2_X4 _sha1_round_add_79_4_U48  ( .A1(_sha1_round_N344 ), .A2(rnd_q[151]),.ZN(_sha1_round_add_79_4_n158 ) );
NAND3_X4 _sha1_round_add_79_4_U47  ( .A1(_sha1_round_add_79_4_n309 ), .A2(_sha1_round_add_79_4_n310 ), .A3(_sha1_round_add_79_4_n311 ), .ZN(_sha1_round_add_79_4_n304 ) );
NAND2_X4 _sha1_round_add_79_4_U46  ( .A1(_sha1_round_add_79_4_n12 ), .A2(_sha1_round_add_79_4_n304 ), .ZN(_sha1_round_add_79_4_n273 ) );
NAND2_X4 _sha1_round_add_79_4_U45  ( .A1(_sha1_round_add_79_4_n259 ), .A2(_sha1_round_add_79_4_n260 ), .ZN(_sha1_round_add_79_4_n248 ) );
INV_X2 _sha1_round_add_79_4_U44  ( .A(_sha1_round_N331 ), .ZN(_sha1_round_add_79_4_n288 ) );
AND2_X4 _sha1_round_add_79_4_U43  ( .A1(_sha1_round_add_79_4_n136 ), .A2(_sha1_round_add_79_4_n145 ), .ZN(_sha1_round_add_79_4_n2 ) );
NOR2_X2 _sha1_round_add_79_4_U42  ( .A1(_sha1_round_add_79_4_n297 ), .A2(_sha1_round_add_79_4_n8 ), .ZN(_sha1_round_add_79_4_n293 ) );
NOR2_X2 _sha1_round_add_79_4_U41  ( .A1(_sha1_round_add_79_4_n293 ), .A2(_sha1_round_add_79_4_n10 ), .ZN(_sha1_round_add_79_4_n291 ) );
NAND2_X2 _sha1_round_add_79_4_U40  ( .A1(_sha1_round_add_79_4_n141 ), .A2(_sha1_round_add_79_4_n142 ), .ZN(_sha1_round_add_79_4_n24 ) );
NAND2_X2 _sha1_round_add_79_4_U39  ( .A1(_sha1_round_add_79_4_n192 ), .A2(_sha1_round_add_79_4_n193 ), .ZN(_sha1_round_add_79_4_n178 ) );
NOR2_X2 _sha1_round_add_79_4_U38  ( .A1(rnd_q[143]), .A2(_sha1_round_N336 ),.ZN(_sha1_round_add_79_4_n218 ) );
NAND2_X2 _sha1_round_add_79_4_U37  ( .A1(_sha1_round_add_79_4_n209 ), .A2(_sha1_round_add_79_4_n210 ), .ZN(_sha1_round_add_79_4_n97 ) );
NOR2_X2 _sha1_round_add_79_4_U36  ( .A1(_sha1_round_N335 ), .A2(rnd_q[142]),.ZN(_sha1_round_add_79_4_n47 ) );
INV_X4 _sha1_round_add_79_4_U35  ( .A(_sha1_round_N327 ), .ZN(_sha1_round_add_79_4_n321 ) );
NAND2_X2 _sha1_round_add_79_4_U34  ( .A1(_sha1_round_add_79_4_n321 ), .A2(_sha1_round_add_79_4_n322 ), .ZN(_sha1_round_add_79_4_n307 ) );
NAND2_X2 _sha1_round_add_79_4_U33  ( .A1(_sha1_round_add_79_4_n326 ), .A2(_sha1_round_add_79_4_n327 ), .ZN(_sha1_round_add_79_4_n313 ) );
NOR2_X2 _sha1_round_add_79_4_U32  ( .A1(_sha1_round_add_79_4_n339 ), .A2(_sha1_round_add_79_4_n340 ), .ZN(_sha1_round_add_79_4_n338 ) );
NAND2_X2 _sha1_round_add_79_4_U31  ( .A1(_sha1_round_add_79_4_n143 ), .A2(_sha1_round_add_79_4_n144 ), .ZN(_sha1_round_add_79_4_n141 ) );
NOR2_X2 _sha1_round_add_79_4_U30  ( .A1(_sha1_round_add_79_4_n278 ), .A2(_sha1_round_add_79_4_n48 ), .ZN(_sha1_round_add_79_4_n276 ) );
NOR2_X4 _sha1_round_add_79_4_U29  ( .A1(_sha1_round_add_79_4_n96 ), .A2(_sha1_round_add_79_4_n155 ), .ZN(_sha1_round_add_79_4_n130 ) );
NAND2_X4 _sha1_round_add_79_4_U28  ( .A1(_sha1_round_add_79_4_n248 ), .A2(_sha1_round_add_79_4_n249 ), .ZN(_sha1_round_add_79_4_n246 ) );
NAND2_X4 _sha1_round_add_79_4_U27  ( .A1(_sha1_round_add_79_4_n246 ), .A2(_sha1_round_add_79_4_n247 ), .ZN(_sha1_round_add_79_4_n209 ) );
NAND2_X4 _sha1_round_add_79_4_U26  ( .A1(_sha1_round_add_79_4_n200 ), .A2(_sha1_round_add_79_4_n201 ), .ZN(_sha1_round_add_79_4_n153 ) );
NAND2_X4 _sha1_round_add_79_4_U25  ( .A1(_sha1_round_add_79_4_n153 ), .A2(_sha1_round_add_79_4_n154 ), .ZN(_sha1_round_add_79_4_n199 ) );
NOR2_X4 _sha1_round_add_79_4_U24  ( .A1(_sha1_round_add_79_4_n267 ), .A2(_sha1_round_add_79_4_n268 ), .ZN(_sha1_round_add_79_4_n250 ) );
XNOR2_X1 _sha1_round_add_79_4_U23  ( .A(_sha1_round_add_79_4_n165 ), .B(_sha1_round_add_79_4_n191 ), .ZN(sha1_round_wire[152]) );
NOR2_X4 _sha1_round_add_79_4_U22  ( .A1(_sha1_round_add_79_4_n122 ), .A2(_sha1_round_add_79_4_n121 ), .ZN(_sha1_round_add_79_4_n118 ) );
NAND2_X4 _sha1_round_add_79_4_U21  ( .A1(_sha1_round_add_79_4_n161 ), .A2(_sha1_round_add_79_4_n162 ), .ZN(_sha1_round_add_79_4_n159 ) );
NAND2_X4 _sha1_round_add_79_4_U20  ( .A1(_sha1_round_add_79_4_n171 ), .A2(_sha1_round_add_79_4_n172 ), .ZN(_sha1_round_add_79_4_n163 ) );
NAND2_X4 _sha1_round_add_79_4_U19  ( .A1(_sha1_round_add_79_4_n170 ), .A2(_sha1_round_add_79_4_n163 ), .ZN(_sha1_round_add_79_4_n166 ) );
NAND2_X4 _sha1_round_add_79_4_U18  ( .A1(_sha1_round_add_79_4_n211 ), .A2(_sha1_round_add_79_4_n154 ), .ZN(_sha1_round_add_79_4_n100 ) );
INV_X8 _sha1_round_add_79_4_U17  ( .A(_sha1_round_add_79_4_n100 ), .ZN(_sha1_round_add_79_4_n136 ) );
NAND2_X4 _sha1_round_add_79_4_U16  ( .A1(_sha1_round_add_79_4_n13 ), .A2(_sha1_round_add_79_4_n97 ), .ZN(_sha1_round_add_79_4_n232 ) );
NAND2_X1 _sha1_round_add_79_4_U15  ( .A1(_sha1_round_add_79_4_n44 ), .A2(_sha1_round_add_79_4_n97 ), .ZN(_sha1_round_add_79_4_n137 ) );
NAND2_X1 _sha1_round_add_79_4_U14  ( .A1(_sha1_round_N342 ), .A2(rnd_q[149]),.ZN(_sha1_round_add_79_4_n174 ) );
NAND3_X4 _sha1_round_add_79_4_U13  ( .A1(_sha1_round_add_79_4_n336 ), .A2(_sha1_round_add_79_4_n337 ), .A3(_sha1_round_add_79_4_n338 ), .ZN(_sha1_round_add_79_4_n64 ) );
AND2_X2 _sha1_round_add_79_4_U12  ( .A1(_sha1_round_add_79_4_n157 ), .A2(_sha1_round_add_79_4_n156 ), .ZN(_sha1_round_add_79_4_n1 ) );
INV_X1 _sha1_round_add_79_4_U11  ( .A(_sha1_round_add_79_4_n130 ), .ZN(_sha1_round_add_79_4_n152 ) );
AND2_X4 _sha1_round_add_79_4_U10  ( .A1(_sha1_round_add_79_4_n307 ), .A2(_sha1_round_add_79_4_n313 ), .ZN(_sha1_round_add_79_4_n309 ) );
INV_X4 _sha1_round_add_79_4_U9  ( .A(_sha1_round_add_79_4_n36 ), .ZN(_sha1_round_add_79_4_n110 ) );
NOR2_X1 _sha1_round_add_79_4_U8  ( .A1(_sha1_round_add_79_4_n113 ), .A2(_sha1_round_add_79_4_n36 ), .ZN(_sha1_round_add_79_4_n133 ) );
NAND2_X4 _sha1_round_add_79_4_U7  ( .A1(_sha1_round_add_79_4_n34 ), .A2(_sha1_round_add_79_4_n35 ), .ZN(sha1_round_wire[159]) );
NOR2_X4 _sha1_round_add_79_4_U6  ( .A1(_sha1_round_add_79_4_n253 ), .A2(_sha1_round_add_79_4_n254 ), .ZN(_sha1_round_add_79_4_n251 ) );
NAND2_X1 _sha1_round_add_79_4_U5  ( .A1(_sha1_round_add_79_4_n18 ), .A2(_sha1_round_add_79_4_n307 ), .ZN(_sha1_round_add_79_4_n317 ) );
INV_X4 _sha1_round_add_79_4_U4  ( .A(_sha1_round_N343 ), .ZN(_sha1_round_add_79_4_n168 ) );
NAND2_X4 _sha1_round_add_79_4_U3  ( .A1(_sha1_round_add_79_4_n30 ), .A2(_sha1_round_add_79_4_n31 ), .ZN(sha1_round_wire[151]) );
NAND2_X4 _sha1_round_add_79_4_U2  ( .A1(_sha1_round_add_79_4_n28 ), .A2(_sha1_round_add_79_4_n29 ), .ZN(_sha1_round_add_79_4_n31 ) );
INV_X4 _sha1_round_add_79_3_U418  ( .A(_sha1_round_N256 ), .ZN(_sha1_round_add_79_3_n386 ) );
INV_X4 _sha1_round_add_79_3_U417  ( .A(_sha1_round_N288 ), .ZN(_sha1_round_add_79_3_n387 ) );
NAND3_X4 _sha1_round_add_79_3_U416  ( .A1(_sha1_round_add_79_3_n383 ), .A2(_sha1_round_add_79_3_n378 ), .A3(_sha1_round_add_79_3_n384 ), .ZN(_sha1_round_add_79_3_n239 ) );
NOR2_X4 _sha1_round_add_79_3_U415  ( .A1(_sha1_round_N259 ), .A2(_sha1_round_N291 ), .ZN(_sha1_round_add_79_3_n88 ) );
NAND3_X4 _sha1_round_add_79_3_U414  ( .A1(_sha1_round_add_79_3_n239 ), .A2(_sha1_round_add_79_3_n16 ), .A3(_sha1_round_add_79_3_n380 ), .ZN(_sha1_round_add_79_3_n81 ) );
NAND2_X2 _sha1_round_add_79_3_U413  ( .A1(_sha1_round_N284 ), .A2(_sha1_round_N252 ), .ZN(_sha1_round_add_79_3_n375 ) );
NAND2_X2 _sha1_round_add_79_3_U412  ( .A1(_sha1_round_N285 ), .A2(_sha1_round_N253 ), .ZN(_sha1_round_add_79_3_n376 ) );
NAND2_X2 _sha1_round_add_79_3_U411  ( .A1(_sha1_round_add_79_3_n375 ), .A2(_sha1_round_add_79_3_n376 ), .ZN(_sha1_round_add_79_3_n372 ) );
INV_X4 _sha1_round_add_79_3_U410  ( .A(_sha1_round_add_79_3_n146 ), .ZN(_sha1_round_add_79_3_n373 ) );
INV_X4 _sha1_round_add_79_3_U409  ( .A(_sha1_round_add_79_3_n111 ), .ZN(_sha1_round_add_79_3_n374 ) );
NAND4_X2 _sha1_round_add_79_3_U408  ( .A1(_sha1_round_add_79_3_n372 ), .A2(_sha1_round_add_79_3_n314 ), .A3(_sha1_round_add_79_3_n373 ), .A4(_sha1_round_add_79_3_n374 ), .ZN(_sha1_round_add_79_3_n371 ) );
NAND2_X2 _sha1_round_add_79_3_U407  ( .A1(_sha1_round_N287 ), .A2(_sha1_round_N255 ), .ZN(_sha1_round_add_79_3_n309 ) );
INV_X4 _sha1_round_add_79_3_U406  ( .A(_sha1_round_N293 ), .ZN(_sha1_round_add_79_3_n367 ) );
INV_X4 _sha1_round_add_79_3_U405  ( .A(_sha1_round_N261 ), .ZN(_sha1_round_add_79_3_n368 ) );
INV_X4 _sha1_round_add_79_3_U404  ( .A(_sha1_round_add_79_3_n74 ), .ZN(_sha1_round_add_79_3_n365 ) );
NOR2_X4 _sha1_round_add_79_3_U403  ( .A1(_sha1_round_add_79_3_n364 ), .A2(_sha1_round_add_79_3_n365 ), .ZN(_sha1_round_add_79_3_n360 ) );
INV_X4 _sha1_round_add_79_3_U402  ( .A(_sha1_round_add_79_3_n348 ), .ZN(_sha1_round_add_79_3_n359 ) );
INV_X4 _sha1_round_add_79_3_U401  ( .A(_sha1_round_N294 ), .ZN(_sha1_round_add_79_3_n362 ) );
XNOR2_X2 _sha1_round_add_79_3_U400  ( .A(_sha1_round_add_79_3_n360 ), .B(_sha1_round_add_79_3_n361 ), .ZN(_sha1_round_N326 ) );
INV_X4 _sha1_round_add_79_3_U399  ( .A(_sha1_round_N295 ), .ZN(_sha1_round_add_79_3_n356 ) );
NAND2_X2 _sha1_round_add_79_3_U398  ( .A1(_sha1_round_add_79_3_n76 ), .A2(_sha1_round_add_79_3_n74 ), .ZN(_sha1_round_add_79_3_n346 ) );
NOR2_X4 _sha1_round_add_79_3_U397  ( .A1(_sha1_round_add_79_3_n321 ), .A2(_sha1_round_add_79_3_n322 ), .ZN(_sha1_round_add_79_3_n347 ) );
NAND3_X4 _sha1_round_add_79_3_U396  ( .A1(_sha1_round_add_79_3_n347 ), .A2(_sha1_round_add_79_3_n346 ), .A3(_sha1_round_add_79_3_n73 ), .ZN(_sha1_round_add_79_3_n245 ) );
INV_X4 _sha1_round_add_79_3_U395  ( .A(_sha1_round_add_79_3_n84 ), .ZN(_sha1_round_add_79_3_n342 ) );
INV_X4 _sha1_round_add_79_3_U394  ( .A(_sha1_round_N297 ), .ZN(_sha1_round_add_79_3_n336 ) );
NAND2_X2 _sha1_round_add_79_3_U393  ( .A1(_sha1_round_add_79_3_n336 ), .A2(_sha1_round_add_79_3_n337 ), .ZN(_sha1_round_add_79_3_n298 ) );
NAND2_X2 _sha1_round_add_79_3_U392  ( .A1(_sha1_round_N297 ), .A2(_sha1_round_N265 ), .ZN(_sha1_round_add_79_3_n294 ) );
NAND2_X2 _sha1_round_add_79_3_U391  ( .A1(_sha1_round_add_79_3_n52 ), .A2(_sha1_round_add_79_3_n294 ), .ZN(_sha1_round_add_79_3_n335 ) );
INV_X4 _sha1_round_add_79_3_U390  ( .A(_sha1_round_N298 ), .ZN(_sha1_round_add_79_3_n331 ) );
XNOR2_X2 _sha1_round_add_79_3_U389  ( .A(_sha1_round_add_79_3_n329 ), .B(_sha1_round_add_79_3_n330 ), .ZN(_sha1_round_N330 ) );
INV_X4 _sha1_round_add_79_3_U388  ( .A(_sha1_round_N299 ), .ZN(_sha1_round_add_79_3_n326 ) );
INV_X4 _sha1_round_add_79_3_U387  ( .A(_sha1_round_N267 ), .ZN(_sha1_round_add_79_3_n327 ) );
XNOR2_X2 _sha1_round_add_79_3_U386  ( .A(_sha1_round_add_79_3_n324 ), .B(_sha1_round_add_79_3_n325 ), .ZN(_sha1_round_N331 ) );
INV_X4 _sha1_round_add_79_3_U385  ( .A(_sha1_round_add_79_3_n323 ), .ZN(_sha1_round_add_79_3_n246 ) );
INV_X4 _sha1_round_add_79_3_U384  ( .A(_sha1_round_add_79_3_n314 ), .ZN(_sha1_round_add_79_3_n107 ) );
NAND2_X2 _sha1_round_add_79_3_U383  ( .A1(_sha1_round_N284 ), .A2(_sha1_round_N252 ), .ZN(_sha1_round_add_79_3_n313 ) );
NAND2_X2 _sha1_round_add_79_3_U382  ( .A1(_sha1_round_N254 ), .A2(_sha1_round_N286 ), .ZN(_sha1_round_add_79_3_n312 ) );
INV_X4 _sha1_round_add_79_3_U381  ( .A(_sha1_round_add_79_3_n309 ), .ZN(_sha1_round_add_79_3_n106 ) );
NAND2_X2 _sha1_round_add_79_3_U380  ( .A1(_sha1_round_add_79_3_n306 ), .A2(_sha1_round_add_79_3_n307 ), .ZN(_sha1_round_add_79_3_n240 ) );
INV_X4 _sha1_round_add_79_3_U379  ( .A(_sha1_round_add_79_3_n235 ), .ZN(_sha1_round_add_79_3_n296 ) );
NOR2_X4 _sha1_round_add_79_3_U378  ( .A1(_sha1_round_add_79_3_n58 ), .A2(_sha1_round_add_79_3_n295 ), .ZN(_sha1_round_add_79_3_n277 ) );
NOR2_X4 _sha1_round_add_79_3_U377  ( .A1(_sha1_round_N268 ), .A2(_sha1_round_N300 ), .ZN(_sha1_round_add_79_3_n276 ) );
XNOR2_X2 _sha1_round_add_79_3_U376  ( .A(_sha1_round_add_79_3_n288 ), .B(_sha1_round_add_79_3_n289 ), .ZN(_sha1_round_N332 ) );
INV_X4 _sha1_round_add_79_3_U375  ( .A(_sha1_round_N301 ), .ZN(_sha1_round_add_79_3_n285 ) );
XNOR2_X2 _sha1_round_add_79_3_U374  ( .A(_sha1_round_add_79_3_n284 ), .B(_sha1_round_add_79_3_n8 ), .ZN(_sha1_round_N333 ) );
NAND2_X2 _sha1_round_add_79_3_U373  ( .A1(_sha1_round_add_79_3_n269 ), .A2(_sha1_round_add_79_3_n259 ), .ZN(_sha1_round_add_79_3_n268 ) );
INV_X4 _sha1_round_add_79_3_U372  ( .A(_sha1_round_N303 ), .ZN(_sha1_round_add_79_3_n265 ) );
INV_X4 _sha1_round_add_79_3_U371  ( .A(_sha1_round_N271 ), .ZN(_sha1_round_add_79_3_n266 ) );
XNOR2_X2 _sha1_round_add_79_3_U370  ( .A(_sha1_round_add_79_3_n262 ), .B(_sha1_round_add_79_3_n263 ), .ZN(_sha1_round_N335 ) );
INV_X4 _sha1_round_add_79_3_U369  ( .A(_sha1_round_add_79_3_n376 ), .ZN(_sha1_round_add_79_3_n261 ) );
XNOR2_X2 _sha1_round_add_79_3_U368  ( .A(_sha1_round_add_79_3_n313 ), .B(_sha1_round_add_79_3_n260 ), .ZN(_sha1_round_N317 ) );
NAND2_X2 _sha1_round_add_79_3_U367  ( .A1(_sha1_round_N304 ), .A2(_sha1_round_N272 ), .ZN(_sha1_round_add_79_3_n226 ) );
NAND2_X2 _sha1_round_add_79_3_U366  ( .A1(_sha1_round_add_79_3_n226 ), .A2(_sha1_round_add_79_3_n228 ), .ZN(_sha1_round_add_79_3_n229 ) );
INV_X4 _sha1_round_add_79_3_U365  ( .A(_sha1_round_add_79_3_n257 ), .ZN(_sha1_round_add_79_3_n256 ) );
NOR2_X4 _sha1_round_add_79_3_U364  ( .A1(_sha1_round_add_79_3_n253 ), .A2(_sha1_round_add_79_3_n252 ), .ZN(_sha1_round_add_79_3_n230 ) );
INV_X4 _sha1_round_add_79_3_U363  ( .A(_sha1_round_add_79_3_n250 ), .ZN(_sha1_round_add_79_3_n249 ) );
NAND3_X4 _sha1_round_add_79_3_U362  ( .A1(_sha1_round_add_79_3_n232 ), .A2(_sha1_round_add_79_3_n230 ), .A3(_sha1_round_add_79_3_n231 ), .ZN(_sha1_round_add_79_3_n148 ) );
INV_X4 _sha1_round_add_79_3_U361  ( .A(_sha1_round_add_79_3_n218 ), .ZN(_sha1_round_add_79_3_n228 ) );
INV_X4 _sha1_round_add_79_3_U360  ( .A(_sha1_round_N305 ), .ZN(_sha1_round_add_79_3_n224 ) );
INV_X4 _sha1_round_add_79_3_U359  ( .A(_sha1_round_N273 ), .ZN(_sha1_round_add_79_3_n225 ) );
XNOR2_X2 _sha1_round_add_79_3_U358  ( .A(_sha1_round_add_79_3_n222 ), .B(_sha1_round_add_79_3_n223 ), .ZN(_sha1_round_N337 ) );
INV_X4 _sha1_round_add_79_3_U357  ( .A(_sha1_round_add_79_3_n208 ), .ZN(_sha1_round_add_79_3_n220 ) );
NAND2_X2 _sha1_round_add_79_3_U356  ( .A1(_sha1_round_add_79_3_n215 ), .A2(_sha1_round_add_79_3_n216 ), .ZN(_sha1_round_add_79_3_n211 ) );
INV_X4 _sha1_round_add_79_3_U355  ( .A(_sha1_round_N306 ), .ZN(_sha1_round_add_79_3_n213 ) );
INV_X4 _sha1_round_add_79_3_U354  ( .A(_sha1_round_N274 ), .ZN(_sha1_round_add_79_3_n214 ) );
NAND2_X2 _sha1_round_add_79_3_U353  ( .A1(_sha1_round_N306 ), .A2(_sha1_round_N274 ), .ZN(_sha1_round_add_79_3_n209 ) );
NAND2_X2 _sha1_round_add_79_3_U352  ( .A1(_sha1_round_add_79_3_n200 ), .A2(_sha1_round_add_79_3_n209 ), .ZN(_sha1_round_add_79_3_n212 ) );
XNOR2_X2 _sha1_round_add_79_3_U351  ( .A(_sha1_round_add_79_3_n211 ), .B(_sha1_round_add_79_3_n212 ), .ZN(_sha1_round_N338 ) );
INV_X4 _sha1_round_add_79_3_U350  ( .A(_sha1_round_add_79_3_n198 ), .ZN(_sha1_round_add_79_3_n206 ) );
NAND2_X2 _sha1_round_add_79_3_U349  ( .A1(_sha1_round_add_79_3_n204 ), .A2(_sha1_round_add_79_3_n205 ), .ZN(_sha1_round_add_79_3_n202 ) );
NAND2_X2 _sha1_round_add_79_3_U348  ( .A1(_sha1_round_N307 ), .A2(_sha1_round_N275 ), .ZN(_sha1_round_add_79_3_n150 ) );
NAND2_X2 _sha1_round_add_79_3_U347  ( .A1(_sha1_round_add_79_3_n197 ), .A2(_sha1_round_add_79_3_n150 ), .ZN(_sha1_round_add_79_3_n203 ) );
NAND2_X2 _sha1_round_add_79_3_U346  ( .A1(_sha1_round_N308 ), .A2(_sha1_round_N276 ), .ZN(_sha1_round_add_79_3_n174 ) );
INV_X4 _sha1_round_add_79_3_U345  ( .A(_sha1_round_N308 ), .ZN(_sha1_round_add_79_3_n195 ) );
INV_X4 _sha1_round_add_79_3_U344  ( .A(_sha1_round_N276 ), .ZN(_sha1_round_add_79_3_n196 ) );
XNOR2_X2 _sha1_round_add_79_3_U343  ( .A(_sha1_round_add_79_3_n186 ), .B(_sha1_round_add_79_3_n194 ), .ZN(_sha1_round_N340 ) );
NAND2_X2 _sha1_round_add_79_3_U342  ( .A1(_sha1_round_add_79_3_n178 ), .A2(_sha1_round_add_79_3_n186 ), .ZN(_sha1_round_add_79_3_n193 ) );
INV_X4 _sha1_round_add_79_3_U341  ( .A(_sha1_round_N309 ), .ZN(_sha1_round_add_79_3_n191 ) );
INV_X4 _sha1_round_add_79_3_U340  ( .A(_sha1_round_N277 ), .ZN(_sha1_round_add_79_3_n192 ) );
NAND2_X2 _sha1_round_add_79_3_U339  ( .A1(_sha1_round_add_79_3_n172 ), .A2(_sha1_round_add_79_3_n179 ), .ZN(_sha1_round_add_79_3_n183 ) );
INV_X4 _sha1_round_add_79_3_U338  ( .A(_sha1_round_add_79_3_n179 ), .ZN(_sha1_round_add_79_3_n176 ) );
NAND2_X2 _sha1_round_add_79_3_U337  ( .A1(_sha1_round_add_79_3_n185 ), .A2(_sha1_round_add_79_3_n186 ), .ZN(_sha1_round_add_79_3_n184 ) );
NAND2_X2 _sha1_round_add_79_3_U336  ( .A1(_sha1_round_add_79_3_n183 ), .A2(_sha1_round_add_79_3_n184 ), .ZN(_sha1_round_add_79_3_n181 ) );
NAND2_X2 _sha1_round_add_79_3_U335  ( .A1(_sha1_round_N311 ), .A2(_sha1_round_N279 ), .ZN(_sha1_round_add_79_3_n157 ) );
INV_X4 _sha1_round_add_79_3_U334  ( .A(_sha1_round_N311 ), .ZN(_sha1_round_add_79_3_n166 ) );
INV_X4 _sha1_round_add_79_3_U333  ( .A(_sha1_round_N279 ), .ZN(_sha1_round_add_79_3_n167 ) );
NAND2_X2 _sha1_round_add_79_3_U332  ( .A1(_sha1_round_add_79_3_n166 ), .A2(_sha1_round_add_79_3_n167 ), .ZN(_sha1_round_add_79_3_n158 ) );
NOR2_X4 _sha1_round_add_79_3_U331  ( .A1(_sha1_round_add_79_3_n164 ), .A2(_sha1_round_add_79_3_n165 ), .ZN(_sha1_round_add_79_3_n161 ) );
NAND2_X2 _sha1_round_add_79_3_U330  ( .A1(_sha1_round_N312 ), .A2(_sha1_round_N280 ), .ZN(_sha1_round_add_79_3_n136 ) );
INV_X4 _sha1_round_add_79_3_U329  ( .A(_sha1_round_add_79_3_n153 ), .ZN(_sha1_round_add_79_3_n151 ) );
NAND2_X2 _sha1_round_add_79_3_U328  ( .A1(_sha1_round_add_79_3_n64 ), .A2(_sha1_round_add_79_3_n65 ), .ZN(_sha1_round_add_79_3_n127 ) );
INV_X4 _sha1_round_add_79_3_U327  ( .A(_sha1_round_add_79_3_n150 ), .ZN(_sha1_round_add_79_3_n149 ) );
NAND4_X2 _sha1_round_add_79_3_U326  ( .A1(_sha1_round_add_79_3_n129 ), .A2(_sha1_round_add_79_3_n136 ), .A3(_sha1_round_add_79_3_n127 ), .A4(_sha1_round_add_79_3_n126 ), .ZN(_sha1_round_add_79_3_n147 ) );
NAND2_X2 _sha1_round_add_79_3_U325  ( .A1(_sha1_round_N313 ), .A2(_sha1_round_N281 ), .ZN(_sha1_round_add_79_3_n134 ) );
NAND2_X2 _sha1_round_add_79_3_U324  ( .A1(_sha1_round_N286 ), .A2(_sha1_round_N254 ), .ZN(_sha1_round_add_79_3_n110 ) );
NAND2_X2 _sha1_round_add_79_3_U323  ( .A1(_sha1_round_add_79_3_n374 ), .A2(_sha1_round_add_79_3_n110 ), .ZN(_sha1_round_add_79_3_n145 ) );
NAND2_X2 _sha1_round_add_79_3_U322  ( .A1(_sha1_round_add_79_3_n62 ), .A2(_sha1_round_add_79_3_n376 ), .ZN(_sha1_round_add_79_3_n113 ) );
XNOR2_X2 _sha1_round_add_79_3_U321  ( .A(_sha1_round_add_79_3_n145 ), .B(_sha1_round_add_79_3_n113 ), .ZN(_sha1_round_N318 ) );
NAND2_X2 _sha1_round_add_79_3_U320  ( .A1(_sha1_round_N314 ), .A2(_sha1_round_N282 ), .ZN(_sha1_round_add_79_3_n135 ) );
NAND2_X2 _sha1_round_add_79_3_U319  ( .A1(_sha1_round_add_79_3_n135 ), .A2(_sha1_round_add_79_3_n139 ), .ZN(_sha1_round_add_79_3_n141 ) );
XNOR2_X2 _sha1_round_add_79_3_U318  ( .A(_sha1_round_add_79_3_n140 ), .B(_sha1_round_add_79_3_n141 ), .ZN(_sha1_round_N346 ) );
INV_X4 _sha1_round_add_79_3_U317  ( .A(_sha1_round_add_79_3_n139 ), .ZN(_sha1_round_add_79_3_n133 ) );
INV_X4 _sha1_round_add_79_3_U316  ( .A(_sha1_round_add_79_3_n138 ), .ZN(_sha1_round_add_79_3_n137 ) );
INV_X4 _sha1_round_add_79_3_U315  ( .A(_sha1_round_add_79_3_n135 ), .ZN(_sha1_round_add_79_3_n131 ) );
NAND2_X2 _sha1_round_add_79_3_U314  ( .A1(_sha1_round_add_79_3_n128 ), .A2(_sha1_round_add_79_3_n121 ), .ZN(_sha1_round_add_79_3_n117 ) );
INV_X4 _sha1_round_add_79_3_U313  ( .A(_sha1_round_add_79_3_n121 ), .ZN(_sha1_round_add_79_3_n125 ) );
NAND2_X2 _sha1_round_add_79_3_U312  ( .A1(_sha1_round_add_79_3_n120 ), .A2(_sha1_round_add_79_3_n121 ), .ZN(_sha1_round_add_79_3_n119 ) );
NAND4_X2 _sha1_round_add_79_3_U311  ( .A1(_sha1_round_add_79_3_n116 ), .A2(_sha1_round_add_79_3_n117 ), .A3(_sha1_round_add_79_3_n118 ), .A4(_sha1_round_add_79_3_n119 ), .ZN(_sha1_round_add_79_3_n114 ) );
XNOR2_X2 _sha1_round_add_79_3_U310  ( .A(_sha1_round_N315 ), .B(_sha1_round_N283 ), .ZN(_sha1_round_add_79_3_n115 ) );
XNOR2_X2 _sha1_round_add_79_3_U309  ( .A(_sha1_round_add_79_3_n114 ), .B(_sha1_round_add_79_3_n115 ), .ZN(_sha1_round_N347 ) );
INV_X4 _sha1_round_add_79_3_U308  ( .A(_sha1_round_add_79_3_n113 ), .ZN(_sha1_round_add_79_3_n112 ) );
INV_X4 _sha1_round_add_79_3_U307  ( .A(_sha1_round_add_79_3_n110 ), .ZN(_sha1_round_add_79_3_n109 ) );
XNOR2_X2 _sha1_round_add_79_3_U306  ( .A(_sha1_round_add_79_3_n104 ), .B(_sha1_round_add_79_3_n105 ), .ZN(_sha1_round_N319 ) );
NAND2_X2 _sha1_round_add_79_3_U305  ( .A1(_sha1_round_N288 ), .A2(_sha1_round_N256 ), .ZN(_sha1_round_add_79_3_n98 ) );
NAND2_X2 _sha1_round_add_79_3_U304  ( .A1(_sha1_round_add_79_3_n98 ), .A2(_sha1_round_add_79_3_n100 ), .ZN(_sha1_round_add_79_3_n103 ) );
NAND2_X2 _sha1_round_add_79_3_U303  ( .A1(_sha1_round_add_79_3_n93 ), .A2(_sha1_round_add_79_3_n95 ), .ZN(_sha1_round_add_79_3_n97 ) );
INV_X4 _sha1_round_add_79_3_U302  ( .A(_sha1_round_add_79_3_n102 ), .ZN(_sha1_round_add_79_3_n100 ) );
XNOR2_X2 _sha1_round_add_79_3_U301  ( .A(_sha1_round_add_79_3_n97 ), .B(_sha1_round_add_79_3_n94 ), .ZN(_sha1_round_N321 ) );
NAND2_X2 _sha1_round_add_79_3_U300  ( .A1(_sha1_round_add_79_3_n94 ), .A2(_sha1_round_add_79_3_n95 ), .ZN(_sha1_round_add_79_3_n92 ) );
XNOR2_X2 _sha1_round_add_79_3_U299  ( .A(_sha1_round_add_79_3_n63 ), .B(_sha1_round_add_79_3_n91 ), .ZN(_sha1_round_N322 ) );
NAND2_X2 _sha1_round_add_79_3_U298  ( .A1(_sha1_round_add_79_3_n76 ), .A2(_sha1_round_add_79_3_n77 ), .ZN(_sha1_round_add_79_3_n82 ) );
INV_X4 _sha1_round_add_79_3_U297  ( .A(_sha1_round_add_79_3_n81 ), .ZN(_sha1_round_add_79_3_n79 ) );
NAND2_X2 _sha1_round_add_79_3_U296  ( .A1(_sha1_round_add_79_3_n77 ), .A2(_sha1_round_add_79_3_n78 ), .ZN(_sha1_round_add_79_3_n75 ) );
NAND2_X2 _sha1_round_add_79_3_U295  ( .A1(_sha1_round_add_79_3_n75 ), .A2(_sha1_round_add_79_3_n76 ), .ZN(_sha1_round_add_79_3_n71 ) );
XNOR2_X2 _sha1_round_add_79_3_U294  ( .A(_sha1_round_add_79_3_n71 ), .B(_sha1_round_add_79_3_n72 ), .ZN(_sha1_round_N325 ) );
NAND2_X4 _sha1_round_add_79_3_U293  ( .A1(_sha1_round_add_79_3_n234 ), .A2(_sha1_round_add_79_3_n233 ), .ZN(_sha1_round_add_79_3_n232 ) );
NAND3_X2 _sha1_round_add_79_3_U292  ( .A1(_sha1_round_add_79_3_n19 ), .A2(_sha1_round_add_79_3_n350 ), .A3(_sha1_round_add_79_3_n351 ), .ZN(_sha1_round_add_79_3_n303 ) );
NAND2_X4 _sha1_round_add_79_3_U291  ( .A1(_sha1_round_add_79_3_n66 ), .A2(_sha1_round_add_79_3_n148 ), .ZN(_sha1_round_add_79_3_n180 ) );
NAND2_X1 _sha1_round_add_79_3_U290  ( .A1(_sha1_round_add_79_3_n148 ), .A2(_sha1_round_add_79_3_n207 ), .ZN(_sha1_round_add_79_3_n216 ) );
NAND2_X1 _sha1_round_add_79_3_U289  ( .A1(_sha1_round_add_79_3_n206 ), .A2(_sha1_round_add_79_3_n148 ), .ZN(_sha1_round_add_79_3_n205 ) );
NAND2_X1 _sha1_round_add_79_3_U288  ( .A1(_sha1_round_N299 ), .A2(_sha1_round_N267 ), .ZN(_sha1_round_add_79_3_n291 ) );
NAND2_X1 _sha1_round_add_79_3_U287  ( .A1(_sha1_round_add_79_3_n291 ), .A2(_sha1_round_add_79_3_n247 ), .ZN(_sha1_round_add_79_3_n325 ) );
NAND3_X2 _sha1_round_add_79_3_U286  ( .A1(_sha1_round_add_79_3_n249 ), .A2(_sha1_round_add_79_3_n248 ), .A3(_sha1_round_add_79_3_n247 ), .ZN(_sha1_round_add_79_3_n231 ) );
NAND2_X4 _sha1_round_add_79_3_U285  ( .A1(_sha1_round_add_79_3_n286 ), .A2(_sha1_round_add_79_3_n285 ), .ZN(_sha1_round_add_79_3_n274 ) );
NOR2_X1 _sha1_round_add_79_3_U284  ( .A1(_sha1_round_add_79_3_n87 ), .A2(_sha1_round_add_79_3_n385 ), .ZN(_sha1_round_add_79_3_n86 ) );
NAND3_X2 _sha1_round_add_79_3_U283  ( .A1(_sha1_round_add_79_3_n50 ), .A2(_sha1_round_add_79_3_n302 ), .A3(_sha1_round_add_79_3_n245 ), .ZN(_sha1_round_add_79_3_n341 ) );
NAND2_X1 _sha1_round_add_79_3_U282  ( .A1(_sha1_round_add_79_3_n302 ), .A2(_sha1_round_add_79_3_n20 ), .ZN(_sha1_round_add_79_3_n355 ) );
NAND2_X2 _sha1_round_add_79_3_U281  ( .A1(_sha1_round_add_79_3_n148 ), .A2(_sha1_round_add_79_3_n228 ), .ZN(_sha1_round_add_79_3_n227 ) );
NAND2_X4 _sha1_round_add_79_3_U280  ( .A1(_sha1_round_add_79_3_n327 ), .A2(_sha1_round_add_79_3_n326 ), .ZN(_sha1_round_add_79_3_n247 ) );
NOR2_X2 _sha1_round_add_79_3_U279  ( .A1(_sha1_round_add_79_3_n276 ), .A2(_sha1_round_add_79_3_n69 ), .ZN(_sha1_round_add_79_3_n289 ) );
NAND2_X1 _sha1_round_add_79_3_U278  ( .A1(_sha1_round_add_79_3_n208 ), .A2(_sha1_round_add_79_3_n219 ), .ZN(_sha1_round_add_79_3_n223 ) );
NAND3_X2 _sha1_round_add_79_3_U277  ( .A1(_sha1_round_N272 ), .A2(_sha1_round_N304 ), .A3(_sha1_round_add_79_3_n219 ), .ZN(_sha1_round_add_79_3_n210 ) );
NAND2_X1 _sha1_round_add_79_3_U276  ( .A1(_sha1_round_N309 ), .A2(_sha1_round_N277 ), .ZN(_sha1_round_add_79_3_n173 ) );
NAND2_X1 _sha1_round_add_79_3_U275  ( .A1(_sha1_round_N258 ), .A2(_sha1_round_N290 ), .ZN(_sha1_round_add_79_3_n381 ) );
NAND2_X1 _sha1_round_add_79_3_U274  ( .A1(_sha1_round_add_79_3_n73 ), .A2(_sha1_round_add_79_3_n74 ), .ZN(_sha1_round_add_79_3_n72 ) );
NAND2_X4 _sha1_round_add_79_3_U273  ( .A1(_sha1_round_add_79_3_n266 ), .A2(_sha1_round_add_79_3_n265 ), .ZN(_sha1_round_add_79_3_n251 ) );
NAND2_X1 _sha1_round_add_79_3_U272  ( .A1(_sha1_round_N310 ), .A2(_sha1_round_N278 ), .ZN(_sha1_round_add_79_3_n160 ) );
NOR3_X2 _sha1_round_add_79_3_U271  ( .A1(_sha1_round_add_79_3_n13 ), .A2(_sha1_round_add_79_3_n146 ), .A3(_sha1_round_add_79_3_n111 ), .ZN(_sha1_round_add_79_3_n310 ) );
OR2_X4 _sha1_round_add_79_3_U270  ( .A1(_sha1_round_N252 ), .A2(_sha1_round_N284 ), .ZN(_sha1_round_add_79_3_n70 ) );
AND2_X2 _sha1_round_add_79_3_U269  ( .A1(_sha1_round_add_79_3_n313 ), .A2(_sha1_round_add_79_3_n70 ), .ZN(_sha1_round_N316 ) );
AND2_X2 _sha1_round_add_79_3_U268  ( .A1(_sha1_round_N300 ), .A2(_sha1_round_N268 ), .ZN(_sha1_round_add_79_3_n69 ) );
AND2_X2 _sha1_round_add_79_3_U267  ( .A1(_sha1_round_N290 ), .A2(_sha1_round_N258 ), .ZN(_sha1_round_add_79_3_n68 ) );
NOR2_X2 _sha1_round_add_79_3_U266  ( .A1(_sha1_round_add_79_3_n275 ), .A2(_sha1_round_add_79_3_n276 ), .ZN(_sha1_round_add_79_3_n273 ) );
NOR2_X2 _sha1_round_add_79_3_U265  ( .A1(_sha1_round_add_79_3_n310 ), .A2(_sha1_round_add_79_3_n311 ), .ZN(_sha1_round_add_79_3_n306 ) );
NOR2_X2 _sha1_round_add_79_3_U264  ( .A1(_sha1_round_add_79_3_n106 ), .A2(_sha1_round_add_79_3_n308 ), .ZN(_sha1_round_add_79_3_n307 ) );
NAND2_X1 _sha1_round_add_79_3_U263  ( .A1(_sha1_round_N302 ), .A2(_sha1_round_N270 ), .ZN(_sha1_round_add_79_3_n259 ) );
NOR2_X2 _sha1_round_add_79_3_U262  ( .A1(_sha1_round_add_79_3_n88 ), .A2(_sha1_round_add_79_3_n381 ), .ZN(_sha1_round_add_79_3_n323 ) );
OR2_X2 _sha1_round_add_79_3_U261  ( .A1(_sha1_round_N314 ), .A2(_sha1_round_N282 ), .ZN(_sha1_round_add_79_3_n139 ) );
OR2_X2 _sha1_round_add_79_3_U260  ( .A1(_sha1_round_N312 ), .A2(_sha1_round_N280 ), .ZN(_sha1_round_add_79_3_n152 ) );
OR2_X2 _sha1_round_add_79_3_U259  ( .A1(_sha1_round_N313 ), .A2(_sha1_round_N281 ), .ZN(_sha1_round_add_79_3_n138 ) );
NOR2_X2 _sha1_round_add_79_3_U258  ( .A1(_sha1_round_N253 ), .A2(_sha1_round_N285 ), .ZN(_sha1_round_add_79_3_n146 ) );
NOR2_X1 _sha1_round_add_79_3_U257  ( .A1(_sha1_round_add_79_3_n111 ), .A2(_sha1_round_add_79_3_n112 ), .ZN(_sha1_round_add_79_3_n108 ) );
INV_X4 _sha1_round_add_79_3_U256  ( .A(_sha1_round_add_79_3_n244 ), .ZN(_sha1_round_add_79_3_n87 ) );
NOR2_X1 _sha1_round_add_79_3_U255  ( .A1(_sha1_round_add_79_3_n102 ), .A2(_sha1_round_add_79_3_n96 ), .ZN(_sha1_round_add_79_3_n318 ) );
AND2_X2 _sha1_round_add_79_3_U254  ( .A1(_sha1_round_add_79_3_n92 ), .A2(_sha1_round_add_79_3_n93 ), .ZN(_sha1_round_add_79_3_n63 ) );
NOR2_X1 _sha1_round_add_79_3_U253  ( .A1(_sha1_round_add_79_3_n176 ), .A2(_sha1_round_add_79_3_n188 ), .ZN(_sha1_round_add_79_3_n185 ) );
NOR2_X2 _sha1_round_add_79_3_U252  ( .A1(_sha1_round_add_79_3_n258 ), .A2(_sha1_round_add_79_3_n259 ), .ZN(_sha1_round_add_79_3_n252 ) );
NOR3_X2 _sha1_round_add_79_3_U251  ( .A1(_sha1_round_add_79_3_n241 ), .A2(_sha1_round_add_79_3_n4 ), .A3(_sha1_round_add_79_3_n243 ), .ZN(_sha1_round_add_79_3_n304 ) );
AND2_X2 _sha1_round_add_79_3_U250  ( .A1(_sha1_round_add_79_3_n136 ), .A2(_sha1_round_add_79_3_n129 ), .ZN(_sha1_round_add_79_3_n144 ) );
NOR2_X2 _sha1_round_add_79_3_U249  ( .A1(_sha1_round_add_79_3_n133 ), .A2(_sha1_round_add_79_3_n137 ), .ZN(_sha1_round_add_79_3_n121 ) );
NAND2_X2 _sha1_round_add_79_3_U248  ( .A1(_sha1_round_add_79_3_n341 ), .A2(_sha1_round_add_79_3_n299 ), .ZN(_sha1_round_add_79_3_n340 ) );
NOR2_X2 _sha1_round_add_79_3_U247  ( .A1(_sha1_round_add_79_3_n322 ), .A2(_sha1_round_add_79_3_n348 ), .ZN(_sha1_round_add_79_3_n242 ) );
NOR2_X1 _sha1_round_add_79_3_U246  ( .A1(_sha1_round_add_79_3_n68 ), .A2(_sha1_round_add_79_3_n90 ), .ZN(_sha1_round_add_79_3_n91 ) );
NOR2_X2 _sha1_round_add_79_3_U245  ( .A1(_sha1_round_add_79_3_n89 ), .A2(_sha1_round_add_79_3_n68 ), .ZN(_sha1_round_add_79_3_n85 ) );
NOR2_X2 _sha1_round_add_79_3_U244  ( .A1(_sha1_round_add_79_3_n220 ), .A2(_sha1_round_add_79_3_n221 ), .ZN(_sha1_round_add_79_3_n215 ) );
NOR2_X2 _sha1_round_add_79_3_U243  ( .A1(_sha1_round_add_79_3_n108 ), .A2(_sha1_round_add_79_3_n109 ), .ZN(_sha1_round_add_79_3_n104 ) );
NOR2_X2 _sha1_round_add_79_3_U242  ( .A1(_sha1_round_add_79_3_n319 ), .A2(_sha1_round_add_79_3_n320 ), .ZN(_sha1_round_add_79_3_n351 ) );
XNOR2_X2 _sha1_round_add_79_3_U241  ( .A(_sha1_round_add_79_3_n202 ), .B(_sha1_round_add_79_3_n203 ), .ZN(_sha1_round_N339 ) );
NOR2_X1 _sha1_round_add_79_3_U240  ( .A1(_sha1_round_add_79_3_n125 ), .A2(_sha1_round_add_79_3_n126 ), .ZN(_sha1_round_add_79_3_n124 ) );
NOR2_X1 _sha1_round_add_79_3_U239  ( .A1(_sha1_round_add_79_3_n125 ), .A2(_sha1_round_add_79_3_n127 ), .ZN(_sha1_round_add_79_3_n123 ) );
NOR2_X2 _sha1_round_add_79_3_U238  ( .A1(_sha1_round_add_79_3_n123 ), .A2(_sha1_round_add_79_3_n124 ), .ZN(_sha1_round_add_79_3_n118 ) );
NOR2_X1 _sha1_round_add_79_3_U237  ( .A1(_sha1_round_add_79_3_n352 ), .A2(_sha1_round_add_79_3_n81 ), .ZN(_sha1_round_add_79_3_n349 ) );
AND4_X2 _sha1_round_add_79_3_U236  ( .A1(_sha1_round_add_79_3_n304 ), .A2(_sha1_round_add_79_3_n5 ), .A3(_sha1_round_add_79_3_n239 ), .A4(_sha1_round_add_79_3_n305 ), .ZN(_sha1_round_add_79_3_n58 ) );
NOR2_X1 _sha1_round_add_79_3_U235  ( .A1(_sha1_round_add_79_3_n359 ), .A2(_sha1_round_add_79_3_n321 ), .ZN(_sha1_round_add_79_3_n361 ) );
NOR2_X1 _sha1_round_add_79_3_U234  ( .A1(_sha1_round_add_79_3_n107 ), .A2(_sha1_round_add_79_3_n312 ), .ZN(_sha1_round_add_79_3_n311 ) );
NOR3_X1 _sha1_round_add_79_3_U233  ( .A1(_sha1_round_add_79_3_n376 ), .A2(_sha1_round_add_79_3_n107 ), .A3(_sha1_round_add_79_3_n111 ), .ZN(_sha1_round_add_79_3_n308 ) );
NAND3_X2 _sha1_round_add_79_3_U232  ( .A1(_sha1_round_N254 ), .A2(_sha1_round_N286 ), .A3(_sha1_round_add_79_3_n314 ), .ZN(_sha1_round_add_79_3_n370 ) );
OR2_X4 _sha1_round_add_79_3_U231  ( .A1(_sha1_round_N296 ), .A2(_sha1_round_N264 ), .ZN(_sha1_round_add_79_3_n299 ) );
NAND3_X2 _sha1_round_add_79_3_U230  ( .A1(_sha1_round_N257 ), .A2(_sha1_round_N289 ), .A3(_sha1_round_add_79_3_n378 ), .ZN(_sha1_round_add_79_3_n382 ) );
OR2_X4 _sha1_round_add_79_3_U229  ( .A1(_sha1_round_N307 ), .A2(_sha1_round_N275 ), .ZN(_sha1_round_add_79_3_n197 ) );
INV_X1 _sha1_round_add_79_3_U228  ( .A(_sha1_round_add_79_3_n96 ), .ZN(_sha1_round_add_79_3_n95 ) );
AND2_X2 _sha1_round_add_79_3_U227  ( .A1(_sha1_round_add_79_3_n157 ), .A2(_sha1_round_add_79_3_n158 ), .ZN(_sha1_round_add_79_3_n60 ) );
INV_X1 _sha1_round_add_79_3_U226  ( .A(_sha1_round_add_79_3_n251 ), .ZN(_sha1_round_add_79_3_n258 ) );
INV_X4 _sha1_round_add_79_3_U225  ( .A(_sha1_round_add_79_3_n197 ), .ZN(_sha1_round_add_79_3_n67 ) );
INV_X1 _sha1_round_add_79_3_U224  ( .A(_sha1_round_add_79_3_n177 ), .ZN(_sha1_round_add_79_3_n175 ) );
AND2_X2 _sha1_round_add_79_3_U223  ( .A1(_sha1_round_add_79_3_n301 ), .A2(_sha1_round_add_79_3_n299 ), .ZN(_sha1_round_add_79_3_n57 ) );
XNOR2_X2 _sha1_round_add_79_3_U222  ( .A(_sha1_round_add_79_3_n344 ), .B(_sha1_round_add_79_3_n57 ), .ZN(_sha1_round_N328 ) );
NOR2_X1 _sha1_round_add_79_3_U221  ( .A1(_sha1_round_add_79_3_n133 ), .A2(_sha1_round_add_79_3_n134 ), .ZN(_sha1_round_add_79_3_n132 ) );
NOR3_X1 _sha1_round_add_79_3_U220  ( .A1(_sha1_round_add_79_3_n130 ), .A2(_sha1_round_add_79_3_n131 ), .A3(_sha1_round_add_79_3_n132 ), .ZN(_sha1_round_add_79_3_n116 ) );
NOR2_X1 _sha1_round_add_79_3_U219  ( .A1(_sha1_round_add_79_3_n125 ), .A2(_sha1_round_add_79_3_n136 ), .ZN(_sha1_round_add_79_3_n130 ) );
OR2_X4 _sha1_round_add_79_3_U218  ( .A1(_sha1_round_add_79_3_n146 ), .A2(_sha1_round_add_79_3_n313 ), .ZN(_sha1_round_add_79_3_n62 ) );
NOR2_X1 _sha1_round_add_79_3_U217  ( .A1(_sha1_round_add_79_3_n106 ), .A2(_sha1_round_add_79_3_n107 ), .ZN(_sha1_round_add_79_3_n105 ) );
INV_X1 _sha1_round_add_79_3_U216  ( .A(_sha1_round_add_79_3_n259 ), .ZN(_sha1_round_add_79_3_n280 ) );
INV_X1 _sha1_round_add_79_3_U215  ( .A(_sha1_round_add_79_3_n254 ), .ZN(_sha1_round_add_79_3_n264 ) );
NOR2_X1 _sha1_round_add_79_3_U214  ( .A1(_sha1_round_add_79_3_n261 ), .A2(_sha1_round_add_79_3_n146 ), .ZN(_sha1_round_add_79_3_n260 ) );
XOR2_X2 _sha1_round_add_79_3_U213  ( .A(_sha1_round_add_79_3_n349 ), .B(_sha1_round_add_79_3_n82 ), .Z(_sha1_round_N324 ) );
NOR2_X1 _sha1_round_add_79_3_U212  ( .A1(_sha1_round_add_79_3_n83 ), .A2(_sha1_round_add_79_3_n84 ), .ZN(_sha1_round_add_79_3_n352 ) );
NOR2_X1 _sha1_round_add_79_3_U211  ( .A1(_sha1_round_add_79_3_n264 ), .A2(_sha1_round_add_79_3_n258 ), .ZN(_sha1_round_add_79_3_n263 ) );
AND3_X4 _sha1_round_add_79_3_U210  ( .A1(_sha1_round_add_79_3_n200 ), .A2(_sha1_round_add_79_3_n197 ), .A3(_sha1_round_add_79_3_n201 ), .ZN(_sha1_round_add_79_3_n64 ) );
NAND2_X1 _sha1_round_add_79_3_U209  ( .A1(_sha1_round_N298 ), .A2(_sha1_round_N266 ), .ZN(_sha1_round_add_79_3_n292 ) );
XNOR2_X2 _sha1_round_add_79_3_U208  ( .A(_sha1_round_add_79_3_n51 ), .B(_sha1_round_add_79_3_n1 ), .ZN(_sha1_round_N344 ) );
INV_X1 _sha1_round_add_79_3_U207  ( .A(_sha1_round_add_79_3_n101 ), .ZN(_sha1_round_add_79_3_n83 ) );
INV_X1 _sha1_round_add_79_3_U206  ( .A(_sha1_round_add_79_3_n122 ), .ZN(_sha1_round_add_79_3_n120 ) );
NOR2_X2 _sha1_round_add_79_3_U205  ( .A1(_sha1_round_add_79_3_n272 ), .A2(_sha1_round_add_79_3_n18 ), .ZN(_sha1_round_add_79_3_n267 ) );
NOR2_X2 _sha1_round_add_79_3_U204  ( .A1(_sha1_round_add_79_3_n276 ), .A2(_sha1_round_add_79_3_n272 ), .ZN(_sha1_round_add_79_3_n287 ) );
NAND2_X2 _sha1_round_add_79_3_U203  ( .A1(_sha1_round_N291 ), .A2(_sha1_round_N259 ), .ZN(_sha1_round_add_79_3_n244 ) );
NOR2_X2 _sha1_round_add_79_3_U202  ( .A1(_sha1_round_add_79_3_n250 ), .A2(_sha1_round_add_79_3_n290 ), .ZN(_sha1_round_add_79_3_n55 ) );
INV_X4 _sha1_round_add_79_3_U201  ( .A(_sha1_round_add_79_3_n4 ), .ZN(_sha1_round_add_79_3_n50 ) );
INV_X1 _sha1_round_add_79_3_U200  ( .A(_sha1_round_add_79_3_n274 ), .ZN(_sha1_round_add_79_3_n283 ) );
NOR2_X2 _sha1_round_add_79_3_U199  ( .A1(_sha1_round_add_79_3_n161 ), .A2(_sha1_round_add_79_3_n163 ), .ZN(_sha1_round_add_79_3_n169 ) );
NAND2_X4 _sha1_round_add_79_3_U198  ( .A1(_sha1_round_add_79_3_n331 ), .A2(_sha1_round_add_79_3_n332 ), .ZN(_sha1_round_add_79_3_n297 ) );
NAND2_X1 _sha1_round_add_79_3_U197  ( .A1(_sha1_round_add_79_3_n297 ), .A2(_sha1_round_add_79_3_n292 ), .ZN(_sha1_round_add_79_3_n330 ) );
NAND2_X1 _sha1_round_add_79_3_U196  ( .A1(_sha1_round_N305 ), .A2(_sha1_round_N273 ), .ZN(_sha1_round_add_79_3_n208 ) );
NOR2_X4 _sha1_round_add_79_3_U195  ( .A1(_sha1_round_add_79_3_n277 ), .A2(_sha1_round_add_79_3_n55 ), .ZN(_sha1_round_add_79_3_n288 ) );
NOR2_X4 _sha1_round_add_79_3_U194  ( .A1(_sha1_round_add_79_3_n277 ), .A2(_sha1_round_add_79_3_n55 ), .ZN(_sha1_round_add_79_3_n272 ) );
NAND2_X1 _sha1_round_add_79_3_U193  ( .A1(_sha1_round_add_79_3_n201 ), .A2(_sha1_round_add_79_3_n200 ), .ZN(_sha1_round_add_79_3_n204 ) );
INV_X4 _sha1_round_add_79_3_U192  ( .A(_sha1_round_add_79_3_n165 ), .ZN(_sha1_round_add_79_3_n187 ) );
NOR2_X2 _sha1_round_add_79_3_U191  ( .A1(_sha1_round_add_79_3_n287 ), .A2(_sha1_round_add_79_3_n69 ), .ZN(_sha1_round_add_79_3_n284 ) );
INV_X4 _sha1_round_add_79_3_U190  ( .A(_sha1_round_add_79_3_n180 ), .ZN(_sha1_round_add_79_3_n164 ) );
INV_X4 _sha1_round_add_79_3_U189  ( .A(_sha1_round_add_79_3_n178 ), .ZN(_sha1_round_add_79_3_n188 ) );
NAND2_X1 _sha1_round_add_79_3_U188  ( .A1(_sha1_round_add_79_3_n174 ), .A2(_sha1_round_add_79_3_n178 ), .ZN(_sha1_round_add_79_3_n194 ) );
NAND2_X2 _sha1_round_add_79_3_U187  ( .A1(_sha1_round_add_79_3_n69 ), .A2(_sha1_round_add_79_3_n274 ), .ZN(_sha1_round_add_79_3_n270 ) );
INV_X4 _sha1_round_add_79_3_U186  ( .A(_sha1_round_add_79_3_n279 ), .ZN(_sha1_round_add_79_3_n47 ) );
NAND2_X4 _sha1_round_add_79_3_U185  ( .A1(_sha1_round_add_79_3_n48 ), .A2(_sha1_round_add_79_3_n49 ), .ZN(_sha1_round_N334 ) );
NAND2_X4 _sha1_round_add_79_3_U184  ( .A1(_sha1_round_add_79_3_n46 ), .A2(_sha1_round_add_79_3_n47 ), .ZN(_sha1_round_add_79_3_n49 ) );
NAND2_X2 _sha1_round_add_79_3_U183  ( .A1(_sha1_round_add_79_3_n278 ), .A2(_sha1_round_add_79_3_n279 ), .ZN(_sha1_round_add_79_3_n48 ) );
NAND2_X4 _sha1_round_add_79_3_U182  ( .A1(_sha1_round_add_79_3_n10 ), .A2(_sha1_round_add_79_3_n178 ), .ZN(_sha1_round_add_79_3_n163 ) );
NAND4_X2 _sha1_round_add_79_3_U181  ( .A1(_sha1_round_add_79_3_n126 ), .A2(_sha1_round_add_79_3_n144 ), .A3(_sha1_round_add_79_3_n127 ), .A4(_sha1_round_add_79_3_n122 ), .ZN(_sha1_round_add_79_3_n143 ) );
NOR2_X2 _sha1_round_add_79_3_U180  ( .A1(_sha1_round_add_79_3_n198 ), .A2(_sha1_round_add_79_3_n67 ), .ZN(_sha1_round_add_79_3_n66 ) );
AND2_X4 _sha1_round_add_79_3_U179  ( .A1(_sha1_round_add_79_3_n151 ), .A2(_sha1_round_add_79_3_n152 ), .ZN(_sha1_round_add_79_3_n65 ) );
INV_X4 _sha1_round_add_79_3_U178  ( .A(_sha1_round_add_79_3_n60 ), .ZN(_sha1_round_add_79_3_n43 ) );
INV_X4 _sha1_round_add_79_3_U177  ( .A(_sha1_round_add_79_3_n168 ), .ZN(_sha1_round_add_79_3_n42 ) );
NAND2_X4 _sha1_round_add_79_3_U176  ( .A1(_sha1_round_add_79_3_n45 ), .A2(_sha1_round_add_79_3_n44 ), .ZN(_sha1_round_N343 ) );
NAND2_X4 _sha1_round_add_79_3_U175  ( .A1(_sha1_round_add_79_3_n42 ), .A2(_sha1_round_add_79_3_n43 ), .ZN(_sha1_round_add_79_3_n45 ) );
NAND2_X2 _sha1_round_add_79_3_U174  ( .A1(_sha1_round_add_79_3_n168 ), .A2(_sha1_round_add_79_3_n60 ), .ZN(_sha1_round_add_79_3_n44 ) );
NAND2_X1 _sha1_round_add_79_3_U173  ( .A1(_sha1_round_add_79_3_n173 ), .A2(_sha1_round_add_79_3_n179 ), .ZN(_sha1_round_add_79_3_n190 ) );
INV_X2 _sha1_round_add_79_3_U172  ( .A(_sha1_round_add_79_3_n190 ), .ZN(_sha1_round_add_79_3_n39 ) );
INV_X4 _sha1_round_add_79_3_U171  ( .A(_sha1_round_add_79_3_n189 ), .ZN(_sha1_round_add_79_3_n38 ) );
NAND2_X4 _sha1_round_add_79_3_U170  ( .A1(_sha1_round_add_79_3_n40 ), .A2(_sha1_round_add_79_3_n41 ), .ZN(_sha1_round_N341 ) );
NAND2_X4 _sha1_round_add_79_3_U169  ( .A1(_sha1_round_add_79_3_n38 ), .A2(_sha1_round_add_79_3_n39 ), .ZN(_sha1_round_add_79_3_n41 ) );
NAND2_X2 _sha1_round_add_79_3_U168  ( .A1(_sha1_round_add_79_3_n189 ), .A2(_sha1_round_add_79_3_n190 ), .ZN(_sha1_round_add_79_3_n40 ) );
NAND3_X2 _sha1_round_add_79_3_U167  ( .A1(_sha1_round_add_79_3_n238 ), .A2(_sha1_round_add_79_3_n305 ), .A3(_sha1_round_add_79_3_n15 ), .ZN(_sha1_round_add_79_3_n233 ) );
NAND2_X1 _sha1_round_add_79_3_U166  ( .A1(_sha1_round_add_79_3_n160 ), .A2(_sha1_round_add_79_3_n177 ), .ZN(_sha1_round_add_79_3_n182 ) );
INV_X1 _sha1_round_add_79_3_U165  ( .A(_sha1_round_add_79_3_n182 ), .ZN(_sha1_round_add_79_3_n35 ) );
INV_X4 _sha1_round_add_79_3_U164  ( .A(_sha1_round_add_79_3_n181 ), .ZN(_sha1_round_add_79_3_n34 ) );
INV_X1 _sha1_round_add_79_3_U163  ( .A(_sha1_round_add_79_3_n86 ), .ZN(_sha1_round_add_79_3_n31 ) );
INV_X4 _sha1_round_add_79_3_U162  ( .A(_sha1_round_add_79_3_n85 ), .ZN(_sha1_round_add_79_3_n30 ) );
NAND2_X4 _sha1_round_add_79_3_U161  ( .A1(_sha1_round_add_79_3_n32 ), .A2(_sha1_round_add_79_3_n33 ), .ZN(_sha1_round_N323 ) );
NAND2_X4 _sha1_round_add_79_3_U160  ( .A1(_sha1_round_add_79_3_n30 ), .A2(_sha1_round_add_79_3_n31 ), .ZN(_sha1_round_add_79_3_n33 ) );
NAND2_X2 _sha1_round_add_79_3_U159  ( .A1(_sha1_round_add_79_3_n85 ), .A2(_sha1_round_add_79_3_n86 ), .ZN(_sha1_round_add_79_3_n32 ) );
NAND3_X4 _sha1_round_add_79_3_U158  ( .A1(_sha1_round_add_79_3_n208 ), .A2(_sha1_round_add_79_3_n209 ), .A3(_sha1_round_add_79_3_n210 ), .ZN(_sha1_round_add_79_3_n201 ) );
NAND2_X4 _sha1_round_add_79_3_U157  ( .A1(_sha1_round_add_79_3_n29 ), .A2(_sha1_round_add_79_3_n201 ), .ZN(_sha1_round_add_79_3_n199 ) );
AND2_X2 _sha1_round_add_79_3_U156  ( .A1(_sha1_round_add_79_3_n200 ), .A2(_sha1_round_add_79_3_n197 ), .ZN(_sha1_round_add_79_3_n29 ) );
NAND3_X2 _sha1_round_add_79_3_U155  ( .A1(_sha1_round_add_79_3_n245 ), .A2(_sha1_round_add_79_3_n303 ), .A3(_sha1_round_add_79_3_n12 ), .ZN(_sha1_round_add_79_3_n300 ) );
NAND2_X4 _sha1_round_add_79_3_U154  ( .A1(_sha1_round_add_79_3_n328 ), .A2(_sha1_round_add_79_3_n292 ), .ZN(_sha1_round_add_79_3_n324 ) );
INV_X4 _sha1_round_add_79_3_U153  ( .A(_sha1_round_N262 ), .ZN(_sha1_round_add_79_3_n363 ) );
NAND2_X1 _sha1_round_add_79_3_U152  ( .A1(_sha1_round_N303 ), .A2(_sha1_round_N271 ), .ZN(_sha1_round_add_79_3_n254 ) );
NAND2_X1 _sha1_round_add_79_3_U151  ( .A1(_sha1_round_add_79_3_n282 ), .A2(_sha1_round_add_79_3_n256 ), .ZN(_sha1_round_add_79_3_n269 ) );
NOR2_X2 _sha1_round_add_79_3_U150  ( .A1(_sha1_round_add_79_3_n90 ), .A2(_sha1_round_add_79_3_n63 ), .ZN(_sha1_round_add_79_3_n89 ) );
NOR2_X2 _sha1_round_add_79_3_U149  ( .A1(_sha1_round_add_79_3_n267 ), .A2(_sha1_round_add_79_3_n268 ), .ZN(_sha1_round_add_79_3_n262 ) );
INV_X1 _sha1_round_add_79_3_U148  ( .A(_sha1_round_add_79_3_n88 ), .ZN(_sha1_round_add_79_3_n377 ) );
NAND2_X2 _sha1_round_add_79_3_U147  ( .A1(_sha1_round_add_79_3_n76 ), .A2(_sha1_round_add_79_3_n80 ), .ZN(_sha1_round_add_79_3_n28 ) );
NOR2_X2 _sha1_round_add_79_3_U146  ( .A1(_sha1_round_add_79_3_n319 ), .A2(_sha1_round_add_79_3_n320 ), .ZN(_sha1_round_add_79_3_n316 ) );
NOR2_X2 _sha1_round_add_79_3_U145  ( .A1(_sha1_round_N291 ), .A2(_sha1_round_N259 ), .ZN(_sha1_round_add_79_3_n385 ) );
NOR2_X2 _sha1_round_add_79_3_U144  ( .A1(_sha1_round_add_79_3_n321 ), .A2(_sha1_round_add_79_3_n322 ), .ZN(_sha1_round_add_79_3_n315 ) );
AND2_X4 _sha1_round_add_79_3_U143  ( .A1(_sha1_round_add_79_3_n134 ), .A2(_sha1_round_add_79_3_n138 ), .ZN(_sha1_round_add_79_3_n27 ) );
XNOR2_X2 _sha1_round_add_79_3_U142  ( .A(_sha1_round_add_79_3_n56 ), .B(_sha1_round_add_79_3_n27 ), .ZN(_sha1_round_N345 ) );
NOR2_X2 _sha1_round_add_79_3_U141  ( .A1(_sha1_round_add_79_3_n28 ), .A2(_sha1_round_add_79_3_n81 ), .ZN(_sha1_round_add_79_3_n26 ) );
OR2_X4 _sha1_round_add_79_3_U140  ( .A1(_sha1_round_N292 ), .A2(_sha1_round_N260 ), .ZN(_sha1_round_add_79_3_n77 ) );
INV_X1 _sha1_round_add_79_3_U139  ( .A(_sha1_round_add_79_3_n129 ), .ZN(_sha1_round_add_79_3_n128 ) );
NOR2_X2 _sha1_round_add_79_3_U138  ( .A1(_sha1_round_add_79_3_n26 ), .A2(_sha1_round_add_79_3_n366 ), .ZN(_sha1_round_add_79_3_n364 ) );
NOR2_X1 _sha1_round_add_79_3_U137  ( .A1(_sha1_round_add_79_3_n345 ), .A2(_sha1_round_add_79_3_n341 ), .ZN(_sha1_round_add_79_3_n344 ) );
NAND2_X2 _sha1_round_add_79_3_U136  ( .A1(_sha1_round_N294 ), .A2(_sha1_round_N262 ), .ZN(_sha1_round_add_79_3_n348 ) );
NAND2_X1 _sha1_round_add_79_3_U135  ( .A1(_sha1_round_add_79_3_n336 ), .A2(_sha1_round_add_79_3_n337 ), .ZN(_sha1_round_add_79_3_n52 ) );
OR2_X2 _sha1_round_add_79_3_U134  ( .A1(_sha1_round_add_79_3_n293 ), .A2(_sha1_round_add_79_3_n294 ), .ZN(_sha1_round_add_79_3_n61 ) );
AND3_X4 _sha1_round_add_79_3_U133  ( .A1(_sha1_round_add_79_3_n61 ), .A2(_sha1_round_add_79_3_n292 ), .A3(_sha1_round_add_79_3_n291 ), .ZN(_sha1_round_add_79_3_n250 ) );
OR2_X4 _sha1_round_add_79_3_U132  ( .A1(_sha1_round_N310 ), .A2(_sha1_round_N278 ), .ZN(_sha1_round_add_79_3_n177 ) );
INV_X4 _sha1_round_add_79_3_U131  ( .A(_sha1_round_add_79_3_n353 ), .ZN(_sha1_round_add_79_3_n23 ) );
NAND2_X4 _sha1_round_add_79_3_U130  ( .A1(_sha1_round_add_79_3_n24 ), .A2(_sha1_round_add_79_3_n25 ), .ZN(_sha1_round_N327 ) );
NAND2_X4 _sha1_round_add_79_3_U129  ( .A1(_sha1_round_add_79_3_n23 ), .A2(_sha1_round_add_79_3_n355 ), .ZN(_sha1_round_add_79_3_n25 ) );
NAND2_X2 _sha1_round_add_79_3_U128  ( .A1(_sha1_round_add_79_3_n353 ), .A2(_sha1_round_add_79_3_n354 ), .ZN(_sha1_round_add_79_3_n24 ) );
NAND2_X2 _sha1_round_add_79_3_U127  ( .A1(_sha1_round_add_79_3_n14 ), .A2(_sha1_round_add_79_3_n377 ), .ZN(_sha1_round_add_79_3_n84 ) );
INV_X4 _sha1_round_add_79_3_U126  ( .A(_sha1_round_N269 ), .ZN(_sha1_round_add_79_3_n286 ) );
NAND2_X1 _sha1_round_add_79_3_U125  ( .A1(_sha1_round_N301 ), .A2(_sha1_round_N269 ), .ZN(_sha1_round_add_79_3_n271 ) );
NAND2_X2 _sha1_round_add_79_3_U124  ( .A1(_sha1_round_add_79_3_n181 ), .A2(_sha1_round_add_79_3_n182 ), .ZN(_sha1_round_add_79_3_n36 ) );
OR2_X4 _sha1_round_add_79_3_U123  ( .A1(_sha1_round_N287 ), .A2(_sha1_round_N255 ), .ZN(_sha1_round_add_79_3_n314 ) );
INV_X4 _sha1_round_add_79_3_U122  ( .A(_sha1_round_add_79_3_n297 ), .ZN(_sha1_round_add_79_3_n293 ) );
INV_X4 _sha1_round_add_79_3_U121  ( .A(_sha1_round_add_79_3_n21 ), .ZN(_sha1_round_add_79_3_n237 ) );
NAND3_X2 _sha1_round_add_79_3_U120  ( .A1(_sha1_round_add_79_3_n22 ), .A2(_sha1_round_add_79_3_n247 ), .A3(_sha1_round_add_79_3_n297 ), .ZN(_sha1_round_add_79_3_n21 ) );
NAND2_X2 _sha1_round_add_79_3_U119  ( .A1(_sha1_round_add_79_3_n164 ), .A2(_sha1_round_add_79_3_n65 ), .ZN(_sha1_round_add_79_3_n122 ) );
NAND2_X1 _sha1_round_add_79_3_U118  ( .A1(_sha1_round_add_79_3_n79 ), .A2(_sha1_round_add_79_3_n80 ), .ZN(_sha1_round_add_79_3_n78 ) );
NAND2_X1 _sha1_round_add_79_3_U117  ( .A1(_sha1_round_add_79_3_n17 ), .A2(_sha1_round_add_79_3_n356 ), .ZN(_sha1_round_add_79_3_n20 ) );
INV_X1 _sha1_round_add_79_3_U116  ( .A(_sha1_round_add_79_3_n7 ), .ZN(_sha1_round_add_79_3_n18 ) );
INV_X4 _sha1_round_add_79_3_U115  ( .A(_sha1_round_add_79_3_n219 ), .ZN(_sha1_round_add_79_3_n217 ) );
INV_X1 _sha1_round_add_79_3_U114  ( .A(_sha1_round_N263 ), .ZN(_sha1_round_add_79_3_n17 ) );
INV_X4 _sha1_round_add_79_3_U113  ( .A(_sha1_round_N266 ), .ZN(_sha1_round_add_79_3_n332 ) );
AND2_X2 _sha1_round_add_79_3_U112  ( .A1(_sha1_round_add_79_3_n298 ), .A2(_sha1_round_add_79_3_n299 ), .ZN(_sha1_round_add_79_3_n22 ) );
NAND2_X1 _sha1_round_add_79_3_U111  ( .A1(_sha1_round_N293 ), .A2(_sha1_round_N261 ), .ZN(_sha1_round_add_79_3_n74 ) );
NAND2_X1 _sha1_round_add_79_3_U110  ( .A1(_sha1_round_add_79_3_n73 ), .A2(_sha1_round_add_79_3_n77 ), .ZN(_sha1_round_add_79_3_n366 ) );
INV_X4 _sha1_round_add_79_3_U109  ( .A(_sha1_round_add_79_3_n163 ), .ZN(_sha1_round_add_79_3_n162 ) );
NAND4_X1 _sha1_round_add_79_3_U108  ( .A1(_sha1_round_add_79_3_n342 ), .A2(_sha1_round_add_79_3_n343 ), .A3(_sha1_round_add_79_3_n299 ), .A4(_sha1_round_add_79_3_n101 ), .ZN(_sha1_round_add_79_3_n338 ) );
NAND3_X1 _sha1_round_add_79_3_U107  ( .A1(_sha1_round_add_79_3_n81 ), .A2(_sha1_round_add_79_3_n343 ), .A3(_sha1_round_add_79_3_n299 ), .ZN(_sha1_round_add_79_3_n339 ) );
INV_X1 _sha1_round_add_79_3_U106  ( .A(_sha1_round_add_79_3_n303 ), .ZN(_sha1_round_add_79_3_n343 ) );
NOR2_X1 _sha1_round_add_79_3_U105  ( .A1(_sha1_round_add_79_3_n349 ), .A2(_sha1_round_add_79_3_n303 ), .ZN(_sha1_round_add_79_3_n345 ) );
NAND2_X2 _sha1_round_add_79_3_U104  ( .A1(_sha1_round_add_79_3_n173 ), .A2(_sha1_round_add_79_3_n174 ), .ZN(_sha1_round_add_79_3_n172 ) );
XNOR2_X1 _sha1_round_add_79_3_U103  ( .A(_sha1_round_add_79_3_n334 ), .B(_sha1_round_add_79_3_n335 ), .ZN(_sha1_round_N329 ) );
NAND2_X2 _sha1_round_add_79_3_U102  ( .A1(_sha1_round_add_79_3_n142 ), .A2(_sha1_round_add_79_3_n134 ), .ZN(_sha1_round_add_79_3_n140 ) );
INV_X4 _sha1_round_add_79_3_U101  ( .A(_sha1_round_N265 ), .ZN(_sha1_round_add_79_3_n337 ) );
NAND2_X2 _sha1_round_add_79_3_U100  ( .A1(_sha1_round_N296 ), .A2(_sha1_round_N264 ), .ZN(_sha1_round_add_79_3_n301 ) );
NOR2_X2 _sha1_round_add_79_3_U99  ( .A1(_sha1_round_add_79_3_n257 ), .A2(_sha1_round_add_79_3_n280 ), .ZN(_sha1_round_add_79_3_n279 ) );
NOR2_X2 _sha1_round_add_79_3_U98  ( .A1(_sha1_round_N270 ), .A2(_sha1_round_N302 ), .ZN(_sha1_round_add_79_3_n257 ) );
NOR2_X2 _sha1_round_add_79_3_U97  ( .A1(_sha1_round_N270 ), .A2(_sha1_round_N302 ), .ZN(_sha1_round_add_79_3_n275 ) );
OR2_X4 _sha1_round_add_79_3_U96  ( .A1(_sha1_round_add_79_3_n382 ), .A2(_sha1_round_add_79_3_n88 ), .ZN(_sha1_round_add_79_3_n16 ) );
NAND2_X2 _sha1_round_add_79_3_U95  ( .A1(_sha1_round_add_79_3_n296 ), .A2(_sha1_round_add_79_3_n237 ), .ZN(_sha1_round_add_79_3_n295 ) );
AND2_X4 _sha1_round_add_79_3_U94  ( .A1(_sha1_round_add_79_3_n239 ), .A2(_sha1_round_add_79_3_n5 ), .ZN(_sha1_round_add_79_3_n15 ) );
INV_X4 _sha1_round_add_79_3_U93  ( .A(_sha1_round_add_79_3_n355 ), .ZN(_sha1_round_add_79_3_n354 ) );
AND2_X4 _sha1_round_add_79_3_U92  ( .A1(_sha1_round_add_79_3_n378 ), .A2(_sha1_round_add_79_3_n379 ), .ZN(_sha1_round_add_79_3_n14 ) );
OR2_X4 _sha1_round_add_79_3_U91  ( .A1(_sha1_round_add_79_3_n107 ), .A2(_sha1_round_add_79_3_n313 ), .ZN(_sha1_round_add_79_3_n13 ) );
AND2_X4 _sha1_round_add_79_3_U90  ( .A1(_sha1_round_add_79_3_n301 ), .A2(_sha1_round_add_79_3_n302 ), .ZN(_sha1_round_add_79_3_n12 ) );
AND2_X4 _sha1_round_add_79_3_U89  ( .A1(_sha1_round_add_79_3_n256 ), .A2(_sha1_round_add_79_3_n251 ), .ZN(_sha1_round_add_79_3_n11 ) );
AND2_X4 _sha1_round_add_79_3_U88  ( .A1(_sha1_round_add_79_3_n179 ), .A2(_sha1_round_add_79_3_n177 ), .ZN(_sha1_round_add_79_3_n10 ) );
NOR2_X2 _sha1_round_add_79_3_U87  ( .A1(_sha1_round_N272 ), .A2(_sha1_round_N304 ), .ZN(_sha1_round_add_79_3_n218 ) );
NAND2_X2 _sha1_round_add_79_3_U86  ( .A1(_sha1_round_add_79_3_n199 ), .A2(_sha1_round_add_79_3_n150 ), .ZN(_sha1_round_add_79_3_n165 ) );
AND4_X4 _sha1_round_add_79_3_U85  ( .A1(_sha1_round_add_79_3_n315 ), .A2(_sha1_round_add_79_3_n316 ), .A3(_sha1_round_add_79_3_n317 ), .A4(_sha1_round_add_79_3_n318 ), .ZN(_sha1_round_add_79_3_n9 ) );
NOR2_X2 _sha1_round_add_79_3_U84  ( .A1(_sha1_round_N256 ), .A2(_sha1_round_N288 ), .ZN(_sha1_round_add_79_3_n102 ) );
NOR2_X2 _sha1_round_add_79_3_U83  ( .A1(_sha1_round_N254 ), .A2(_sha1_round_N286 ), .ZN(_sha1_round_add_79_3_n111 ) );
INV_X4 _sha1_round_add_79_3_U82  ( .A(_sha1_round_N263 ), .ZN(_sha1_round_add_79_3_n357 ) );
AND2_X4 _sha1_round_add_79_3_U81  ( .A1(_sha1_round_add_79_3_n271 ), .A2(_sha1_round_add_79_3_n274 ), .ZN(_sha1_round_add_79_3_n8 ) );
AND2_X4 _sha1_round_add_79_3_U80  ( .A1(_sha1_round_add_79_3_n273 ), .A2(_sha1_round_add_79_3_n274 ), .ZN(_sha1_round_add_79_3_n7 ) );
OR2_X4 _sha1_round_add_79_3_U79  ( .A1(_sha1_round_add_79_3_n283 ), .A2(_sha1_round_add_79_3_n276 ), .ZN(_sha1_round_add_79_3_n6 ) );
AND2_X4 _sha1_round_add_79_3_U78  ( .A1(_sha1_round_add_79_3_n302 ), .A2(_sha1_round_add_79_3_n301 ), .ZN(_sha1_round_add_79_3_n5 ) );
INV_X2 _sha1_round_add_79_3_U77  ( .A(_sha1_round_add_79_3_n247 ), .ZN(_sha1_round_add_79_3_n290 ) );
NOR2_X2 _sha1_round_add_79_3_U76  ( .A1(_sha1_round_add_79_3_n102 ), .A2(_sha1_round_add_79_3_n96 ), .ZN(_sha1_round_add_79_3_n379 ) );
NOR2_X2 _sha1_round_add_79_3_U75  ( .A1(_sha1_round_add_79_3_n96 ), .A2(_sha1_round_add_79_3_n385 ), .ZN(_sha1_round_add_79_3_n384 ) );
NAND2_X2 _sha1_round_add_79_3_U74  ( .A1(_sha1_round_add_79_3_n143 ), .A2(_sha1_round_add_79_3_n138 ), .ZN(_sha1_round_add_79_3_n142 ) );
NAND2_X2 _sha1_round_add_79_3_U73  ( .A1(_sha1_round_N263 ), .A2(_sha1_round_N295 ), .ZN(_sha1_round_add_79_3_n302 ) );
NAND3_X4 _sha1_round_add_79_3_U72  ( .A1(_sha1_round_add_79_3_n244 ), .A2(_sha1_round_add_79_3_n245 ), .A3(_sha1_round_add_79_3_n246 ), .ZN(_sha1_round_add_79_3_n241 ) );
NAND2_X4 _sha1_round_add_79_3_U71  ( .A1(_sha1_round_add_79_3_n329 ), .A2(_sha1_round_add_79_3_n297 ), .ZN(_sha1_round_add_79_3_n328 ) );
NAND2_X2 _sha1_round_add_79_3_U70  ( .A1(_sha1_round_add_79_3_n149 ), .A2(_sha1_round_add_79_3_n65 ), .ZN(_sha1_round_add_79_3_n126 ) );
NAND2_X2 _sha1_round_add_79_3_U69  ( .A1(_sha1_round_add_79_3_n195 ), .A2(_sha1_round_add_79_3_n196 ), .ZN(_sha1_round_add_79_3_n178 ) );
NAND2_X2 _sha1_round_add_79_3_U68  ( .A1(_sha1_round_add_79_3_n213 ), .A2(_sha1_round_add_79_3_n214 ), .ZN(_sha1_round_add_79_3_n200 ) );
INV_X4 _sha1_round_add_79_3_U67  ( .A(_sha1_round_add_79_3_n278 ), .ZN(_sha1_round_add_79_3_n46 ) );
NAND2_X2 _sha1_round_add_79_3_U66  ( .A1(_sha1_round_add_79_3_n98 ), .A2(_sha1_round_add_79_3_n99 ), .ZN(_sha1_round_add_79_3_n94 ) );
NAND2_X2 _sha1_round_add_79_3_U65  ( .A1(_sha1_round_N292 ), .A2(_sha1_round_N260 ), .ZN(_sha1_round_add_79_3_n76 ) );
NOR2_X2 _sha1_round_add_79_3_U64  ( .A1(_sha1_round_add_79_3_n147 ), .A2(_sha1_round_add_79_3_n120 ), .ZN(_sha1_round_add_79_3_n56 ) );
NOR3_X2 _sha1_round_add_79_3_U63  ( .A1(_sha1_round_add_79_3_n241 ), .A2(_sha1_round_add_79_3_n4 ), .A3(_sha1_round_add_79_3_n243 ), .ZN(_sha1_round_add_79_3_n238 ) );
INV_X4 _sha1_round_add_79_3_U62  ( .A(_sha1_round_add_79_3_n53 ), .ZN(_sha1_round_add_79_3_n54 ) );
NOR2_X2 _sha1_round_add_79_3_U61  ( .A1(_sha1_round_add_79_3_n235 ), .A2(_sha1_round_add_79_3_n54 ), .ZN(_sha1_round_add_79_3_n234 ) );
NAND2_X2 _sha1_round_add_79_3_U60  ( .A1(_sha1_round_add_79_3_n11 ), .A2(_sha1_round_add_79_3_n282 ), .ZN(_sha1_round_add_79_3_n255 ) );
NAND2_X2 _sha1_round_add_79_3_U59  ( .A1(_sha1_round_add_79_3_n255 ), .A2(_sha1_round_add_79_3_n254 ), .ZN(_sha1_round_add_79_3_n253 ) );
INV_X4 _sha1_round_add_79_3_U58  ( .A(_sha1_round_add_79_3_n77 ), .ZN(_sha1_round_add_79_3_n319 ) );
NOR2_X2 _sha1_round_add_79_3_U57  ( .A1(_sha1_round_add_79_3_n217 ), .A2(_sha1_round_add_79_3_n218 ), .ZN(_sha1_round_add_79_3_n207 ) );
NOR2_X2 _sha1_round_add_79_3_U56  ( .A1(_sha1_round_add_79_3_n175 ), .A2(_sha1_round_add_79_3_n176 ), .ZN(_sha1_round_add_79_3_n171 ) );
NAND2_X2 _sha1_round_add_79_3_U55  ( .A1(_sha1_round_add_79_3_n171 ), .A2(_sha1_round_add_79_3_n172 ), .ZN(_sha1_round_add_79_3_n159 ) );
NAND2_X2 _sha1_round_add_79_3_U54  ( .A1(_sha1_round_add_79_3_n162 ), .A2(_sha1_round_add_79_3_n158 ), .ZN(_sha1_round_add_79_3_n153 ) );
NOR2_X2 _sha1_round_add_79_3_U53  ( .A1(_sha1_round_add_79_3_n4 ), .A2(_sha1_round_add_79_3_n300 ), .ZN(_sha1_round_add_79_3_n235 ) );
INV_X4 _sha1_round_add_79_3_U52  ( .A(_sha1_round_add_79_3_n19 ), .ZN(_sha1_round_add_79_3_n322 ) );
NAND2_X2 _sha1_round_add_79_3_U51  ( .A1(_sha1_round_add_79_3_n207 ), .A2(_sha1_round_add_79_3_n200 ), .ZN(_sha1_round_add_79_3_n198 ) );
NOR2_X2 _sha1_round_add_79_3_U50  ( .A1(_sha1_round_add_79_3_n386 ), .A2(_sha1_round_add_79_3_n387 ), .ZN(_sha1_round_add_79_3_n383 ) );
INV_X4 _sha1_round_add_79_3_U49  ( .A(_sha1_round_add_79_3_n16 ), .ZN(_sha1_round_add_79_3_n243 ) );
AND2_X4 _sha1_round_add_79_3_U48  ( .A1(_sha1_round_add_79_3_n371 ), .A2(_sha1_round_add_79_3_n370 ), .ZN(_sha1_round_add_79_3_n369 ) );
NAND2_X4 _sha1_round_add_79_3_U47  ( .A1(_sha1_round_add_79_3_n226 ), .A2(_sha1_round_add_79_3_n227 ), .ZN(_sha1_round_add_79_3_n222 ) );
NOR2_X4 _sha1_round_add_79_3_U46  ( .A1(_sha1_round_add_79_3_n87 ), .A2(_sha1_round_add_79_3_n323 ), .ZN(_sha1_round_add_79_3_n380 ) );
NOR2_X4 _sha1_round_add_79_3_U45  ( .A1(_sha1_round_add_79_3_n288 ), .A2(_sha1_round_add_79_3_n6 ), .ZN(_sha1_round_add_79_3_n281 ) );
NOR2_X4 _sha1_round_add_79_3_U44  ( .A1(_sha1_round_add_79_3_n281 ), .A2(_sha1_round_add_79_3_n282 ), .ZN(_sha1_round_add_79_3_n278 ) );
NAND2_X4 _sha1_round_add_79_3_U43  ( .A1(_sha1_round_add_79_3_n7 ), .A2(_sha1_round_add_79_3_n251 ), .ZN(_sha1_round_add_79_3_n236 ) );
INV_X4 _sha1_round_add_79_3_U42  ( .A(_sha1_round_add_79_3_n236 ), .ZN(_sha1_round_add_79_3_n248 ) );
INV_X1 _sha1_round_add_79_3_U41  ( .A(_sha1_round_add_79_3_n210 ), .ZN(_sha1_round_add_79_3_n221 ) );
NAND2_X4 _sha1_round_add_79_3_U40  ( .A1(_sha1_round_add_79_3_n357 ), .A2(_sha1_round_add_79_3_n356 ), .ZN(_sha1_round_add_79_3_n19 ) );
NAND2_X2 _sha1_round_add_79_3_U39  ( .A1(_sha1_round_add_79_3_n34 ), .A2(_sha1_round_add_79_3_n35 ), .ZN(_sha1_round_add_79_3_n37 ) );
NAND2_X2 _sha1_round_add_79_3_U38  ( .A1(_sha1_round_add_79_3_n294 ), .A2(_sha1_round_add_79_3_n333 ), .ZN(_sha1_round_add_79_3_n329 ) );
NOR2_X2 _sha1_round_add_79_3_U37  ( .A1(_sha1_round_add_79_3_n360 ), .A2(_sha1_round_add_79_3_n321 ), .ZN(_sha1_round_add_79_3_n358 ) );
INV_X4 _sha1_round_add_79_3_U36  ( .A(_sha1_round_add_79_3_n350 ), .ZN(_sha1_round_add_79_3_n321 ) );
NAND2_X2 _sha1_round_add_79_3_U35  ( .A1(_sha1_round_add_79_3_n170 ), .A2(_sha1_round_add_79_3_n158 ), .ZN(_sha1_round_add_79_3_n156 ) );
NAND2_X2 _sha1_round_add_79_3_U34  ( .A1(_sha1_round_add_79_3_n156 ), .A2(_sha1_round_add_79_3_n157 ), .ZN(_sha1_round_add_79_3_n154 ) );
NOR2_X2 _sha1_round_add_79_3_U33  ( .A1(_sha1_round_add_79_3_n161 ), .A2(_sha1_round_add_79_3_n153 ), .ZN(_sha1_round_add_79_3_n155 ) );
NAND2_X2 _sha1_round_add_79_3_U32  ( .A1(_sha1_round_add_79_3_n191 ), .A2(_sha1_round_add_79_3_n192 ), .ZN(_sha1_round_add_79_3_n179 ) );
NAND2_X2 _sha1_round_add_79_3_U31  ( .A1(_sha1_round_add_79_3_n9 ), .A2(_sha1_round_add_79_3_n240 ), .ZN(_sha1_round_add_79_3_n305 ) );
NOR2_X4 _sha1_round_add_79_3_U30  ( .A1(_sha1_round_N258 ), .A2(_sha1_round_N290 ), .ZN(_sha1_round_add_79_3_n90 ) );
NOR2_X1 _sha1_round_add_79_3_U29  ( .A1(_sha1_round_add_79_3_n90 ), .A2(_sha1_round_add_79_3_n88 ), .ZN(_sha1_round_add_79_3_n317 ) );
INV_X8 _sha1_round_add_79_3_U28  ( .A(_sha1_round_add_79_3_n90 ), .ZN(_sha1_round_add_79_3_n378 ) );
NAND2_X4 _sha1_round_add_79_3_U27  ( .A1(_sha1_round_add_79_3_n369 ), .A2(_sha1_round_add_79_3_n309 ), .ZN(_sha1_round_add_79_3_n101 ) );
NAND2_X4 _sha1_round_add_79_3_U26  ( .A1(_sha1_round_add_79_3_n100 ), .A2(_sha1_round_add_79_3_n101 ), .ZN(_sha1_round_add_79_3_n99 ) );
XNOR2_X1 _sha1_round_add_79_3_U25  ( .A(_sha1_round_add_79_3_n103 ), .B(_sha1_round_add_79_3_n101 ), .ZN(_sha1_round_N320 ) );
NAND2_X4 _sha1_round_add_79_3_U24  ( .A1(_sha1_round_add_79_3_n342 ), .A2(_sha1_round_add_79_3_n101 ), .ZN(_sha1_round_add_79_3_n80 ) );
NAND2_X4 _sha1_round_add_79_3_U23  ( .A1(_sha1_round_add_79_3_n367 ), .A2(_sha1_round_add_79_3_n368 ), .ZN(_sha1_round_add_79_3_n73 ) );
INV_X8 _sha1_round_add_79_3_U22  ( .A(_sha1_round_add_79_3_n73 ), .ZN(_sha1_round_add_79_3_n320 ) );
NOR2_X4 _sha1_round_add_79_3_U21  ( .A1(_sha1_round_N257 ), .A2(_sha1_round_N289 ), .ZN(_sha1_round_add_79_3_n96 ) );
NAND2_X1 _sha1_round_add_79_3_U20  ( .A1(_sha1_round_N289 ), .A2(_sha1_round_N257 ), .ZN(_sha1_round_add_79_3_n93 ) );
NAND2_X4 _sha1_round_add_79_3_U19  ( .A1(_sha1_round_add_79_3_n187 ), .A2(_sha1_round_add_79_3_n180 ), .ZN(_sha1_round_add_79_3_n186 ) );
NOR2_X2 _sha1_round_add_79_3_U18  ( .A1(_sha1_round_add_79_3_n155 ), .A2(_sha1_round_add_79_3_n154 ), .ZN(_sha1_round_add_79_3_n51 ) );
NOR2_X4 _sha1_round_add_79_3_U17  ( .A1(_sha1_round_add_79_3_n358 ), .A2(_sha1_round_add_79_3_n359 ), .ZN(_sha1_round_add_79_3_n353 ) );
INV_X8 _sha1_round_add_79_3_U16  ( .A(_sha1_round_add_79_3_n3 ), .ZN(_sha1_round_add_79_3_n4 ) );
INV_X4 _sha1_round_add_79_3_U15  ( .A(_sha1_round_add_79_3_n242 ), .ZN(_sha1_round_add_79_3_n3 ) );
NAND4_X4 _sha1_round_add_79_3_U14  ( .A1(_sha1_round_add_79_3_n338 ), .A2(_sha1_round_add_79_3_n339 ), .A3(_sha1_round_add_79_3_n301 ), .A4(_sha1_round_add_79_3_n340 ), .ZN(_sha1_round_add_79_3_n334 ) );
NAND2_X4 _sha1_round_add_79_3_U13  ( .A1(_sha1_round_add_79_3_n334 ), .A2(_sha1_round_add_79_3_n52 ), .ZN(_sha1_round_add_79_3_n333 ) );
NAND2_X4 _sha1_round_add_79_3_U12  ( .A1(_sha1_round_add_79_3_n193 ), .A2(_sha1_round_add_79_3_n174 ), .ZN(_sha1_round_add_79_3_n189 ) );
NAND2_X4 _sha1_round_add_79_3_U11  ( .A1(_sha1_round_add_79_3_n36 ), .A2(_sha1_round_add_79_3_n37 ), .ZN(_sha1_round_N342 ) );
NOR2_X4 _sha1_round_add_79_3_U10  ( .A1(_sha1_round_add_79_3_n236 ), .A2(_sha1_round_add_79_3_n21 ), .ZN(_sha1_round_add_79_3_n53 ) );
NAND2_X4 _sha1_round_add_79_3_U9  ( .A1(_sha1_round_add_79_3_n363 ), .A2(_sha1_round_add_79_3_n362 ), .ZN(_sha1_round_add_79_3_n350 ) );
NAND2_X4 _sha1_round_add_79_3_U8  ( .A1(_sha1_round_add_79_3_n224 ), .A2(_sha1_round_add_79_3_n225 ), .ZN(_sha1_round_add_79_3_n219 ) );
NAND2_X4 _sha1_round_add_79_3_U7  ( .A1(_sha1_round_add_79_3_n154 ), .A2(_sha1_round_add_79_3_n152 ), .ZN(_sha1_round_add_79_3_n129 ) );
NAND2_X4 _sha1_round_add_79_3_U6  ( .A1(_sha1_round_add_79_3_n159 ), .A2(_sha1_round_add_79_3_n160 ), .ZN(_sha1_round_add_79_3_n170 ) );
XNOR2_X1 _sha1_round_add_79_3_U5  ( .A(_sha1_round_add_79_3_n229 ), .B(_sha1_round_add_79_3_n148 ), .ZN(_sha1_round_N336 ) );
AND2_X4 _sha1_round_add_79_3_U4  ( .A1(_sha1_round_add_79_3_n136 ), .A2(_sha1_round_add_79_3_n152 ), .ZN(_sha1_round_add_79_3_n1 ) );
NAND2_X2 _sha1_round_add_79_3_U3  ( .A1(_sha1_round_add_79_3_n270 ), .A2(_sha1_round_add_79_3_n271 ), .ZN(_sha1_round_add_79_3_n282 ) );
NOR2_X4 _sha1_round_add_79_3_U2  ( .A1(_sha1_round_add_79_3_n169 ), .A2(_sha1_round_add_79_3_n170 ), .ZN(_sha1_round_add_79_3_n168 ) );
NAND2_X2 _sha1_round_add_79_U405  ( .A1(_sha1_round_k_23 ), .A2(_sha1_round_f [0]), .ZN(_sha1_round_add_79_n270 ) );
NOR2_X4 _sha1_round_add_79_U404  ( .A1(_sha1_round_add_79_n377 ), .A2(_sha1_round_add_79_n83 ), .ZN(_sha1_round_add_79_n376 ) );
NAND3_X4 _sha1_round_add_79_U403  ( .A1(_sha1_round_add_79_n374 ), .A2(_sha1_round_add_79_n375 ), .A3(_sha1_round_add_79_n376 ), .ZN(_sha1_round_add_79_n109 ) );
INV_X4 _sha1_round_add_79_U402  ( .A(_sha1_round_add_79_n380 ), .ZN(_sha1_round_add_79_n121 ) );
INV_X4 _sha1_round_add_79_U401  ( .A(_sha1_round_add_79_n306 ), .ZN(_sha1_round_add_79_n129 ) );
INV_X4 _sha1_round_add_79_U400  ( .A(_sha1_round_k[13] ), .ZN(_sha1_round_add_79_n354 ) );
INV_X4 _sha1_round_add_79_U399  ( .A(_sha1_round_f [11]), .ZN(_sha1_round_add_79_n355 ) );
INV_X4 _sha1_round_add_79_U398  ( .A(_sha1_round_add_79_n343 ), .ZN(_sha1_round_add_79_n345 ) );
XNOR2_X2 _sha1_round_add_79_U397  ( .A(_sha1_round_add_79_n352 ), .B(_sha1_round_add_79_n353 ), .ZN(_sha1_round_add_79_n351 ) );
INV_X4 _sha1_round_add_79_U396  ( .A(_sha1_round_f [12]), .ZN(_sha1_round_add_79_n350 ) );
NAND2_X2 _sha1_round_add_79_U395  ( .A1(_sha1_round_add_79_n92 ), .A2(_sha1_round_add_79_n350 ), .ZN(_sha1_round_add_79_n313 ) );
NAND2_X2 _sha1_round_add_79_U394  ( .A1(_sha1_round_add_79_n313 ), .A2(_sha1_round_add_79_n302 ), .ZN(_sha1_round_add_79_n337 ) );
NAND2_X2 _sha1_round_add_79_U393  ( .A1(_sha1_round_k_30 ), .A2(_sha1_round_f [8]), .ZN(_sha1_round_add_79_n341 ) );
NAND4_X2 _sha1_round_add_79_U392  ( .A1(_sha1_round_add_79_n341 ), .A2(_sha1_round_add_79_n342 ), .A3(_sha1_round_add_79_n343 ), .A4(_sha1_round_add_79_n344 ), .ZN(_sha1_round_add_79_n339 ) );
XNOR2_X2 _sha1_round_add_79_U391  ( .A(_sha1_round_add_79_n336 ), .B(_sha1_round_add_79_n337 ), .ZN(_sha1_round_N264 ) );
INV_X4 _sha1_round_add_79_U390  ( .A(_sha1_round_add_79_n323 ), .ZN(_sha1_round_add_79_n334 ) );
XNOR2_X2 _sha1_round_add_79_U389  ( .A(_sha1_round_add_79_n333 ), .B(_sha1_round_add_79_n20 ), .ZN(_sha1_round_N265 ) );
INV_X4 _sha1_round_add_79_U388  ( .A(_sha1_round_add_79_n313 ), .ZN(_sha1_round_add_79_n330 ) );
NAND2_X2 _sha1_round_add_79_U387  ( .A1(_sha1_round_add_79_n294 ), .A2(_sha1_round_add_79_n327 ), .ZN(_sha1_round_add_79_n326 ) );
NAND2_X2 _sha1_round_add_79_U386  ( .A1(_sha1_round_k[15] ), .A2(_sha1_round_f [15]), .ZN(_sha1_round_add_79_n295 ) );
INV_X4 _sha1_round_add_79_U385  ( .A(_sha1_round_add_79_n318 ), .ZN(_sha1_round_add_79_n314 ) );
INV_X4 _sha1_round_add_79_U384  ( .A(_sha1_round_add_79_n289 ), .ZN(_sha1_round_add_79_n316 ) );
INV_X4 _sha1_round_add_79_U383  ( .A(_sha1_round_add_79_n238 ), .ZN(_sha1_round_add_79_n297 ) );
NAND3_X2 _sha1_round_add_79_U382  ( .A1(_sha1_round_add_79_n70 ), .A2(_sha1_round_add_79_n306 ), .A3(_sha1_round_add_79_n307 ), .ZN(_sha1_round_add_79_n305 ) );
NAND2_X2 _sha1_round_add_79_U381  ( .A1(_sha1_round_add_79_n304 ), .A2(_sha1_round_add_79_n305 ), .ZN(_sha1_round_add_79_n298 ) );
INV_X4 _sha1_round_add_79_U380  ( .A(_sha1_round_add_79_n303 ), .ZN(_sha1_round_add_79_n300 ) );
INV_X4 _sha1_round_add_79_U379  ( .A(_sha1_round_add_79_n302 ), .ZN(_sha1_round_add_79_n301 ) );
NAND2_X2 _sha1_round_add_79_U378  ( .A1(_sha1_round_k[13] ), .A2(_sha1_round_f [13]), .ZN(_sha1_round_add_79_n296 ) );
INV_X4 _sha1_round_add_79_U377  ( .A(_sha1_round_k_26 ), .ZN(_sha1_round_add_79_n201 ) );
INV_X4 _sha1_round_add_79_U376  ( .A(_sha1_round_f [16]), .ZN(_sha1_round_add_79_n292 ) );
NAND2_X2 _sha1_round_add_79_U375  ( .A1(_sha1_round_add_79_n201 ), .A2(_sha1_round_add_79_n292 ), .ZN(_sha1_round_add_79_n280 ) );
NAND2_X2 _sha1_round_add_79_U374  ( .A1(_sha1_round_add_79_n293 ), .A2(_sha1_round_add_79_n233 ), .ZN(_sha1_round_add_79_n279 ) );
NAND2_X2 _sha1_round_add_79_U373  ( .A1(_sha1_round_add_79_n279 ), .A2(_sha1_round_add_79_n280 ), .ZN(_sha1_round_add_79_n284 ) );
INV_X4 _sha1_round_add_79_U372  ( .A(_sha1_round_add_79_n275 ), .ZN(_sha1_round_add_79_n239 ) );
INV_X4 _sha1_round_add_79_U371  ( .A(_sha1_round_add_79_n280 ), .ZN(_sha1_round_add_79_n278 ) );
NAND2_X2 _sha1_round_add_79_U370  ( .A1(_sha1_round_add_79_n231 ), .A2(_sha1_round_add_79_n279 ), .ZN(_sha1_round_add_79_n274 ) );
XNOR2_X2 _sha1_round_add_79_U369  ( .A(_sha1_round_add_79_n250 ), .B(_sha1_round_add_79_n262 ), .ZN(_sha1_round_N270 ) );
INV_X4 _sha1_round_add_79_U368  ( .A(_sha1_round_add_79_n266 ), .ZN(_sha1_round_add_79_n272 ) );
XNOR2_X2 _sha1_round_add_79_U367  ( .A(_sha1_round_add_79_n270 ), .B(_sha1_round_add_79_n268 ), .ZN(_sha1_round_N253 ) );
INV_X4 _sha1_round_add_79_U366  ( .A(_sha1_round_f [20]), .ZN(_sha1_round_add_79_n265 ) );
NAND2_X2 _sha1_round_add_79_U365  ( .A1(_sha1_round_add_79_n201 ), .A2(_sha1_round_add_79_n265 ), .ZN(_sha1_round_add_79_n259 ) );
NAND2_X2 _sha1_round_add_79_U364  ( .A1(_sha1_round_add_79_n258 ), .A2(_sha1_round_add_79_n259 ), .ZN(_sha1_round_add_79_n264 ) );
NAND2_X2 _sha1_round_add_79_U363  ( .A1(_sha1_round_f [19]), .A2(_sha1_round_k_26 ), .ZN(_sha1_round_add_79_n257 ) );
XNOR2_X2 _sha1_round_add_79_U362  ( .A(_sha1_round_add_79_n254 ), .B(_sha1_round_add_79_n15 ), .ZN(_sha1_round_N273 ) );
INV_X4 _sha1_round_add_79_U361  ( .A(_sha1_round_add_79_n240 ), .ZN(_sha1_round_add_79_n253 ) );
INV_X4 _sha1_round_add_79_U360  ( .A(_sha1_round_add_79_n251 ), .ZN(_sha1_round_add_79_n242 ) );
NAND2_X2 _sha1_round_add_79_U359  ( .A1(_sha1_round_add_79_n248 ), .A2(_sha1_round_add_79_n249 ), .ZN(_sha1_round_add_79_n245 ) );
INV_X4 _sha1_round_add_79_U358  ( .A(_sha1_round_f [22]), .ZN(_sha1_round_add_79_n247 ) );
NAND2_X2 _sha1_round_add_79_U357  ( .A1(_sha1_round_add_79_n91 ), .A2(_sha1_round_add_79_n247 ), .ZN(_sha1_round_add_79_n241 ) );
NAND2_X2 _sha1_round_add_79_U356  ( .A1(_sha1_round_n3370 ), .A2(_sha1_round_f [22]), .ZN(_sha1_round_add_79_n243 ) );
NAND2_X2 _sha1_round_add_79_U355  ( .A1(_sha1_round_add_79_n241 ), .A2(_sha1_round_add_79_n243 ), .ZN(_sha1_round_add_79_n246 ) );
NAND2_X2 _sha1_round_add_79_U354  ( .A1(_sha1_round_add_79_n219 ), .A2(_sha1_round_add_79_n222 ), .ZN(_sha1_round_add_79_n228 ) );
INV_X4 _sha1_round_add_79_U353  ( .A(_sha1_round_add_79_n243 ), .ZN(_sha1_round_add_79_n227 ) );
INV_X4 _sha1_round_add_79_U352  ( .A(_sha1_round_add_79_n237 ), .ZN(_sha1_round_add_79_n230 ) );
INV_X4 _sha1_round_add_79_U351  ( .A(_sha1_round_add_79_n213 ), .ZN(_sha1_round_add_79_n222 ) );
NAND2_X2 _sha1_round_add_79_U350  ( .A1(_sha1_round_add_79_n221 ), .A2(_sha1_round_add_79_n222 ), .ZN(_sha1_round_add_79_n220 ) );
NAND2_X2 _sha1_round_add_79_U349  ( .A1(_sha1_round_add_79_n219 ), .A2(_sha1_round_add_79_n220 ), .ZN(_sha1_round_add_79_n217 ) );
NAND2_X2 _sha1_round_add_79_U348  ( .A1(_sha1_round_f [24]), .A2(_sha1_round_add_79_n89 ), .ZN(_sha1_round_add_79_n196 ) );
XNOR2_X2 _sha1_round_add_79_U347  ( .A(_sha1_round_add_79_n217 ), .B(_sha1_round_add_79_n218 ), .ZN(_sha1_round_add_79_n216 ) );
INV_X4 _sha1_round_add_79_U346  ( .A(_sha1_round_add_79_n216 ), .ZN(_sha1_round_N276 ) );
INV_X4 _sha1_round_add_79_U345  ( .A(_sha1_round_add_79_n196 ), .ZN(_sha1_round_add_79_n214 ) );
INV_X4 _sha1_round_add_79_U344  ( .A(_sha1_round_add_79_n197 ), .ZN(_sha1_round_add_79_n215 ) );
INV_X4 _sha1_round_add_79_U343  ( .A(_sha1_round_f [25]), .ZN(_sha1_round_add_79_n209 ) );
NAND2_X2 _sha1_round_add_79_U342  ( .A1(_sha1_round_add_79_n55 ), .A2(_sha1_round_add_79_n209 ), .ZN(_sha1_round_add_79_n193 ) );
NAND2_X2 _sha1_round_add_79_U341  ( .A1(_sha1_round_add_79_n193 ), .A2(_sha1_round_add_79_n198 ), .ZN(_sha1_round_add_79_n208 ) );
XNOR2_X2 _sha1_round_add_79_U340  ( .A(_sha1_round_add_79_n207 ), .B(_sha1_round_add_79_n208 ), .ZN(_sha1_round_N277 ) );
NAND2_X2 _sha1_round_add_79_U339  ( .A1(_sha1_round_add_79_n206 ), .A2(_sha1_round_add_79_n193 ), .ZN(_sha1_round_add_79_n203 ) );
NAND2_X2 _sha1_round_add_79_U338  ( .A1(_sha1_round_f [26]), .A2(_sha1_round_k_26 ), .ZN(_sha1_round_add_79_n192 ) );
INV_X4 _sha1_round_add_79_U337  ( .A(_sha1_round_f [26]), .ZN(_sha1_round_add_79_n202 ) );
NAND2_X2 _sha1_round_add_79_U336  ( .A1(_sha1_round_add_79_n201 ), .A2(_sha1_round_add_79_n202 ), .ZN(_sha1_round_add_79_n194 ) );
NAND2_X2 _sha1_round_add_79_U335  ( .A1(_sha1_round_add_79_n192 ), .A2(_sha1_round_add_79_n194 ), .ZN(_sha1_round_add_79_n200 ) );
XNOR2_X2 _sha1_round_add_79_U334  ( .A(_sha1_round_add_79_n199 ), .B(_sha1_round_add_79_n200 ), .ZN(_sha1_round_N278 ) );
NAND2_X2 _sha1_round_add_79_U333  ( .A1(_sha1_round_add_79_n1 ), .A2(_sha1_round_add_79_n194 ), .ZN(_sha1_round_add_79_n187 ) );
NAND2_X2 _sha1_round_add_79_U332  ( .A1(_sha1_round_add_79_n191 ), .A2(_sha1_round_add_79_n192 ), .ZN(_sha1_round_add_79_n183 ) );
INV_X4 _sha1_round_add_79_U331  ( .A(_sha1_round_f [27]), .ZN(_sha1_round_add_79_n189 ) );
NAND2_X2 _sha1_round_add_79_U330  ( .A1(_sha1_round_add_79_n55 ), .A2(_sha1_round_add_79_n189 ), .ZN(_sha1_round_add_79_n184 ) );
XNOR2_X2 _sha1_round_add_79_U329  ( .A(_sha1_round_add_79_n188 ), .B(_sha1_round_add_79_n22 ), .ZN(_sha1_round_N279 ) );
INV_X4 _sha1_round_add_79_U328  ( .A(_sha1_round_add_79_n187 ), .ZN(_sha1_round_add_79_n186 ) );
NAND2_X2 _sha1_round_add_79_U327  ( .A1(_sha1_round_add_79_n186 ), .A2(_sha1_round_add_79_n184 ), .ZN(_sha1_round_add_79_n146 ) );
NAND2_X2 _sha1_round_add_79_U326  ( .A1(_sha1_round_add_79_n183 ), .A2(_sha1_round_add_79_n184 ), .ZN(_sha1_round_add_79_n176 ) );
NAND2_X2 _sha1_round_add_79_U325  ( .A1(_sha1_round_add_79_n176 ), .A2(_sha1_round_add_79_n152 ), .ZN(_sha1_round_add_79_n182 ) );
NAND2_X2 _sha1_round_add_79_U324  ( .A1(_sha1_round_n511 ), .A2(_sha1_round_f [28]), .ZN(_sha1_round_add_79_n161 ) );
INV_X4 _sha1_round_add_79_U323  ( .A(_sha1_round_f [28]), .ZN(_sha1_round_add_79_n180 ) );
NAND2_X2 _sha1_round_add_79_U322  ( .A1(_sha1_round_add_79_n88 ), .A2(_sha1_round_add_79_n180 ), .ZN(_sha1_round_add_79_n175 ) );
NAND2_X2 _sha1_round_add_79_U321  ( .A1(_sha1_round_add_79_n161 ), .A2(_sha1_round_add_79_n175 ), .ZN(_sha1_round_add_79_n179 ) );
INV_X4 _sha1_round_add_79_U320  ( .A(_sha1_round_add_79_n161 ), .ZN(_sha1_round_add_79_n177 ) );
INV_X4 _sha1_round_add_79_U319  ( .A(_sha1_round_add_79_n175 ), .ZN(_sha1_round_add_79_n164 ) );
INV_X4 _sha1_round_add_79_U318  ( .A(_sha1_round_add_79_n176 ), .ZN(_sha1_round_add_79_n141 ) );
NAND2_X2 _sha1_round_add_79_U317  ( .A1(_sha1_round_add_79_n141 ), .A2(_sha1_round_add_79_n175 ), .ZN(_sha1_round_add_79_n174 ) );
NAND2_X2 _sha1_round_add_79_U316  ( .A1(_sha1_round_f [29]), .A2(_sha1_round_n825 ), .ZN(_sha1_round_add_79_n162 ) );
NAND2_X2 _sha1_round_add_79_U315  ( .A1(_sha1_round_add_79_n162 ), .A2(_sha1_round_add_79_n165 ), .ZN(_sha1_round_add_79_n171 ) );
XNOR2_X2 _sha1_round_add_79_U314  ( .A(_sha1_round_add_79_n170 ), .B(_sha1_round_add_79_n171 ), .ZN(_sha1_round_N281 ) );
NAND2_X2 _sha1_round_add_79_U313  ( .A1(_sha1_round_add_79_n169 ), .A2(_sha1_round_add_79_n311 ), .ZN(_sha1_round_add_79_n166 ) );
XNOR2_X2 _sha1_round_add_79_U312  ( .A(_sha1_round_add_79_n166 ), .B(_sha1_round_add_79_n134 ), .ZN(_sha1_round_N254 ) );
INV_X4 _sha1_round_add_79_U311  ( .A(_sha1_round_add_79_n165 ), .ZN(_sha1_round_add_79_n160 ) );
INV_X4 _sha1_round_add_79_U310  ( .A(_sha1_round_add_79_n151 ), .ZN(_sha1_round_add_79_n163 ) );
INV_X4 _sha1_round_add_79_U309  ( .A(_sha1_round_add_79_n148 ), .ZN(_sha1_round_add_79_n159 ) );
NAND2_X2 _sha1_round_add_79_U308  ( .A1(_sha1_round_add_79_n141 ), .A2(_sha1_round_add_79_n151 ), .ZN(_sha1_round_add_79_n157 ) );
NAND2_X2 _sha1_round_add_79_U307  ( .A1(_sha1_round_f [30]), .A2(_sha1_round_k_30 ), .ZN(_sha1_round_add_79_n150 ) );
NAND2_X2 _sha1_round_add_79_U306  ( .A1(_sha1_round_add_79_n150 ), .A2(_sha1_round_add_79_n149 ), .ZN(_sha1_round_add_79_n154 ) );
XNOR2_X2 _sha1_round_add_79_U305  ( .A(_sha1_round_add_79_n153 ), .B(_sha1_round_add_79_n154 ), .ZN(_sha1_round_N282 ) );
NAND2_X2 _sha1_round_add_79_U304  ( .A1(_sha1_round_add_79_n151 ), .A2(_sha1_round_add_79_n149 ), .ZN(_sha1_round_add_79_n143 ) );
INV_X4 _sha1_round_add_79_U303  ( .A(_sha1_round_add_79_n149 ), .ZN(_sha1_round_add_79_n147 ) );
INV_X4 _sha1_round_add_79_U302  ( .A(_sha1_round_add_79_n146 ), .ZN(_sha1_round_add_79_n144 ) );
INV_X4 _sha1_round_add_79_U301  ( .A(_sha1_round_add_79_n143 ), .ZN(_sha1_round_add_79_n142 ) );
NAND2_X2 _sha1_round_add_79_U300  ( .A1(_sha1_round_add_79_n141 ), .A2(_sha1_round_add_79_n142 ), .ZN(_sha1_round_add_79_n140 ) );
NAND4_X2 _sha1_round_add_79_U299  ( .A1(_sha1_round_add_79_n137 ), .A2(_sha1_round_add_79_n138 ), .A3(_sha1_round_add_79_n139 ), .A4(_sha1_round_add_79_n140 ), .ZN(_sha1_round_add_79_n135 ) );
XNOR2_X2 _sha1_round_add_79_U298  ( .A(_sha1_round_f [31]), .B(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n136 ) );
XNOR2_X2 _sha1_round_add_79_U297  ( .A(_sha1_round_add_79_n135 ), .B(_sha1_round_add_79_n136 ), .ZN(_sha1_round_N283 ) );
INV_X4 _sha1_round_add_79_U296  ( .A(_sha1_round_add_79_n134 ), .ZN(_sha1_round_add_79_n133 ) );
INV_X4 _sha1_round_add_79_U295  ( .A(_sha1_round_add_79_n311 ), .ZN(_sha1_round_add_79_n131 ) );
XNOR2_X2 _sha1_round_add_79_U294  ( .A(_sha1_round_add_79_n127 ), .B(_sha1_round_add_79_n128 ), .ZN(_sha1_round_N255 ) );
XNOR2_X2 _sha1_round_add_79_U293  ( .A(_sha1_round_add_79_n126 ), .B(_sha1_round_add_79_n63 ), .ZN(_sha1_round_N256 ) );
NAND2_X2 _sha1_round_add_79_U292  ( .A1(_sha1_round_add_79_n125 ), .A2(_sha1_round_add_79_n119 ), .ZN(_sha1_round_add_79_n122 ) );
INV_X4 _sha1_round_add_79_U291  ( .A(_sha1_round_add_79_n124 ), .ZN(_sha1_round_add_79_n123 ) );
XNOR2_X2 _sha1_round_add_79_U290  ( .A(_sha1_round_add_79_n122 ), .B(_sha1_round_add_79_n123 ), .ZN(_sha1_round_N257 ) );
INV_X4 _sha1_round_add_79_U289  ( .A(_sha1_round_add_79_n120 ), .ZN(_sha1_round_add_79_n117 ) );
XNOR2_X2 _sha1_round_add_79_U288  ( .A(_sha1_round_add_79_n115 ), .B(_sha1_round_add_79_n116 ), .ZN(_sha1_round_N258 ) );
NAND2_X2 _sha1_round_add_79_U287  ( .A1(_sha1_round_add_79_n104 ), .A2(_sha1_round_add_79_n105 ), .ZN(_sha1_round_add_79_n102 ) );
INV_X4 _sha1_round_add_79_U286  ( .A(_sha1_round_add_79_n100 ), .ZN(_sha1_round_add_79_n103 ) );
INV_X4 _sha1_round_add_79_U285  ( .A(_sha1_round_add_79_n96 ), .ZN(_sha1_round_add_79_n95 ) );
XNOR2_X2 _sha1_round_add_79_U284  ( .A(_sha1_round_add_79_n93 ), .B(_sha1_round_add_79_n94 ), .ZN(_sha1_round_N261 ) );
NAND2_X1 _sha1_round_add_79_U283  ( .A1(_sha1_round_n2 ), .A2(_sha1_round_f [4]), .ZN(_sha1_round_add_79_n119 ) );
NAND2_X1 _sha1_round_add_79_U282  ( .A1(_sha1_round_f [17]), .A2(_sha1_round_n2 ), .ZN(_sha1_round_add_79_n275 ) );
NAND3_X2 _sha1_round_add_79_U281  ( .A1(_sha1_round_add_79_n109 ), .A2(_sha1_round_add_79_n31 ), .A3(_sha1_round_add_79_n110 ), .ZN(_sha1_round_add_79_n332 ) );
NAND3_X1 _sha1_round_add_79_U280  ( .A1(_sha1_round_add_79_n31 ), .A2(_sha1_round_add_79_n107 ), .A3(_sha1_round_add_79_n106 ), .ZN(_sha1_round_add_79_n338 ) );
NOR2_X1 _sha1_round_add_79_U279  ( .A1(_sha1_round_add_79_n26 ), .A2(_sha1_round_add_79_n129 ), .ZN(_sha1_round_add_79_n128 ) );
NAND3_X2 _sha1_round_add_79_U278  ( .A1(_sha1_round_add_79_n107 ), .A2(_sha1_round_add_79_n121 ), .A3(_sha1_round_add_79_n8 ), .ZN(_sha1_round_add_79_n120 ) );
NAND3_X1 _sha1_round_add_79_U277  ( .A1(_sha1_round_add_79_n151 ), .A2(_sha1_round_add_79_n144 ), .A3(_sha1_round_add_79_n145 ), .ZN(_sha1_round_add_79_n156 ) );
NAND3_X1 _sha1_round_add_79_U276  ( .A1(_sha1_round_add_79_n142 ), .A2(_sha1_round_add_79_n144 ), .A3(_sha1_round_add_79_n145 ), .ZN(_sha1_round_add_79_n139 ) );
NAND2_X4 _sha1_round_add_79_U275  ( .A1(_sha1_round_add_79_n354 ), .A2(_sha1_round_add_79_n355 ), .ZN(_sha1_round_add_79_n340 ) );
INV_X2 _sha1_round_add_79_U274  ( .A(_sha1_round_add_79_n167 ), .ZN(_sha1_round_add_79_n269 ) );
NAND2_X2 _sha1_round_add_79_U273  ( .A1(_sha1_round_add_79_n1 ), .A2(_sha1_round_add_79_n145 ), .ZN(_sha1_round_add_79_n204 ) );
NAND2_X2 _sha1_round_add_79_U272  ( .A1(_sha1_round_add_79_n205 ), .A2(_sha1_round_add_79_n145 ), .ZN(_sha1_round_add_79_n211 ) );
INV_X2 _sha1_round_add_79_U271  ( .A(_sha1_round_add_79_n101 ), .ZN(_sha1_round_add_79_n97 ) );
NOR2_X2 _sha1_round_add_79_U270  ( .A1(_sha1_round_f [7]), .A2(_sha1_round_k_27 ), .ZN(_sha1_round_add_79_n111 ) );
NAND2_X1 _sha1_round_add_79_U269  ( .A1(_sha1_round_add_79_n2 ), .A2(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n375 ) );
NAND3_X2 _sha1_round_add_79_U268  ( .A1(_sha1_round_add_79_n234 ), .A2(_sha1_round_add_79_n235 ), .A3(_sha1_round_add_79_n236 ), .ZN(_sha1_round_add_79_n226 ) );
NOR2_X1 _sha1_round_add_79_U267  ( .A1(_sha1_round_f [0]), .A2(_sha1_round_k_23 ), .ZN(_sha1_round_add_79_n271 ) );
NAND2_X1 _sha1_round_add_79_U266  ( .A1(_sha1_round_add_79_n359 ), .A2(_sha1_round_add_79_n344 ), .ZN(_sha1_round_add_79_n361 ) );
NAND3_X1 _sha1_round_add_79_U265  ( .A1(_sha1_round_add_79_n144 ), .A2(_sha1_round_add_79_n175 ), .A3(_sha1_round_add_79_n145 ), .ZN(_sha1_round_add_79_n173 ) );
INV_X4 _sha1_round_add_79_U264  ( .A(_sha1_round_f [18]), .ZN(_sha1_round_add_79_n262 ) );
NAND2_X2 _sha1_round_add_79_U263  ( .A1(_sha1_round_add_79_n266 ), .A2(_sha1_round_add_79_n267 ), .ZN(_sha1_round_add_79_n263 ) );
AND2_X2 _sha1_round_add_79_U262  ( .A1(_sha1_round_k_27 ), .A2(_sha1_round_f [7]), .ZN(_sha1_round_add_79_n83 ) );
NOR3_X2 _sha1_round_add_79_U261  ( .A1(_sha1_round_add_79_n310 ), .A2(_sha1_round_add_79_n269 ), .A3(_sha1_round_add_79_n129 ), .ZN(_sha1_round_add_79_n309 ) );
NAND3_X1 _sha1_round_add_79_U260  ( .A1(_sha1_round_f [18]), .A2(_sha1_round_add_79_n27 ), .A3(_sha1_round_add_79_n250 ), .ZN(_sha1_round_add_79_n267 ) );
NAND3_X2 _sha1_round_add_79_U259  ( .A1(_sha1_round_add_79_n294 ), .A2(_sha1_round_add_79_n295 ), .A3(_sha1_round_add_79_n24 ), .ZN(_sha1_round_add_79_n288 ) );
AND2_X2 _sha1_round_add_79_U258  ( .A1(_sha1_round_add_79_n257 ), .A2(_sha1_round_add_79_n258 ), .ZN(_sha1_round_add_79_n82 ) );
AND2_X2 _sha1_round_add_79_U257  ( .A1(_sha1_round_add_79_n2 ), .A2(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n81 ) );
NOR2_X2 _sha1_round_add_79_U256  ( .A1(_sha1_round_f [8]), .A2(_sha1_round_k_30 ), .ZN(_sha1_round_add_79_n348 ) );
AND2_X2 _sha1_round_add_79_U255  ( .A1(_sha1_round_n825 ), .A2(_sha1_round_add_79_n33 ), .ZN(_sha1_round_add_79_n80 ) );
NOR2_X1 _sha1_round_add_79_U254  ( .A1(_sha1_round_n2 ), .A2(_sha1_round_f [17]), .ZN(_sha1_round_add_79_n79 ) );
NAND3_X1 _sha1_round_add_79_U253  ( .A1(_sha1_round_f [23]), .A2(_sha1_round_add_79_n25 ), .A3(_sha1_round_k_23 ), .ZN(_sha1_round_add_79_n197 ) );
NOR2_X1 _sha1_round_add_79_U252  ( .A1(_sha1_round_f [23]), .A2(_sha1_round_k_23 ), .ZN(_sha1_round_add_79_n213 ) );
NOR2_X2 _sha1_round_add_79_U251  ( .A1(_sha1_round_add_79_n381 ), .A2(_sha1_round_add_79_n271 ), .ZN(_sha1_round_N252 ) );
INV_X1 _sha1_round_add_79_U250  ( .A(_sha1_round_n511 ), .ZN(_sha1_round_add_79_n88 ) );
INV_X1 _sha1_round_add_79_U249  ( .A(_sha1_round_n3370 ), .ZN(_sha1_round_add_79_n91 ) );
OR2_X2 _sha1_round_add_79_U248  ( .A1(_sha1_round_add_79_n152 ), .A2(_sha1_round_add_79_n143 ), .ZN(_sha1_round_add_79_n137 ) );
INV_X4 _sha1_round_add_79_U247  ( .A(_sha1_round_add_79_n86 ), .ZN(_sha1_round_add_79_n87 ) );
OR2_X4 _sha1_round_add_79_U246  ( .A1(_sha1_round_add_79_n348 ), .A2(_sha1_round_add_79_n103 ), .ZN(_sha1_round_add_79_n77 ) );
XNOR2_X2 _sha1_round_add_79_U245  ( .A(_sha1_round_add_79_n102 ), .B(_sha1_round_add_79_n77 ), .ZN(_sha1_round_N260 ) );
NOR2_X2 _sha1_round_add_79_U244  ( .A1(_sha1_round_add_79_n212 ), .A2(_sha1_round_add_79_n214 ), .ZN(_sha1_round_add_79_n218 ) );
OR2_X4 _sha1_round_add_79_U243  ( .A1(_sha1_round_add_79_n147 ), .A2(_sha1_round_add_79_n148 ), .ZN(_sha1_round_add_79_n75 ) );
AND2_X2 _sha1_round_add_79_U242  ( .A1(_sha1_round_add_79_n150 ), .A2(_sha1_round_add_79_n75 ), .ZN(_sha1_round_add_79_n138 ) );
NAND3_X2 _sha1_round_add_79_U241  ( .A1(_sha1_round_add_79_n230 ), .A2(_sha1_round_add_79_n231 ), .A3(_sha1_round_add_79_n232 ), .ZN(_sha1_round_add_79_n225 ) );
NOR2_X1 _sha1_round_add_79_U240  ( .A1(_sha1_round_add_79_n74 ), .A2(_sha1_round_add_79_n227 ), .ZN(_sha1_round_add_79_n223 ) );
NAND3_X1 _sha1_round_add_79_U239  ( .A1(_sha1_round_add_79_n242 ), .A2(_sha1_round_add_79_n240 ), .A3(_sha1_round_add_79_n250 ), .ZN(_sha1_round_add_79_n249 ) );
OR2_X4 _sha1_round_add_79_U238  ( .A1(_sha1_round_add_79_n160 ), .A2(_sha1_round_add_79_n161 ), .ZN(_sha1_round_add_79_n73 ) );
AND2_X2 _sha1_round_add_79_U237  ( .A1(_sha1_round_add_79_n162 ), .A2(_sha1_round_add_79_n73 ), .ZN(_sha1_round_add_79_n148 ) );
XNOR2_X2 _sha1_round_add_79_U236  ( .A(_sha1_round_add_79_n263 ), .B(_sha1_round_add_79_n264 ), .ZN(_sha1_round_N272 ) );
NOR2_X2 _sha1_round_add_79_U235  ( .A1(_sha1_round_add_79_n163 ), .A2(_sha1_round_add_79_n152 ), .ZN(_sha1_round_add_79_n158 ) );
NOR2_X2 _sha1_round_add_79_U234  ( .A1(_sha1_round_add_79_n164 ), .A2(_sha1_round_add_79_n152 ), .ZN(_sha1_round_add_79_n178 ) );
NOR2_X1 _sha1_round_add_79_U233  ( .A1(_sha1_round_add_79_n349 ), .A2(_sha1_round_add_79_n346 ), .ZN(_sha1_round_add_79_n357 ) );
NOR2_X2 _sha1_round_add_79_U232  ( .A1(_sha1_round_add_79_n212 ), .A2(_sha1_round_add_79_n213 ), .ZN(_sha1_round_add_79_n205 ) );
OR2_X2 _sha1_round_add_79_U231  ( .A1(_sha1_round_add_79_n253 ), .A2(_sha1_round_add_79_n82 ), .ZN(_sha1_round_add_79_n69 ) );
NAND3_X2 _sha1_round_add_79_U230  ( .A1(_sha1_round_add_79_n196 ), .A2(_sha1_round_add_79_n197 ), .A3(_sha1_round_add_79_n198 ), .ZN(_sha1_round_add_79_n195 ) );
NAND3_X2 _sha1_round_add_79_U229  ( .A1(_sha1_round_add_79_n193 ), .A2(_sha1_round_add_79_n194 ), .A3(_sha1_round_add_79_n195 ), .ZN(_sha1_round_add_79_n191 ) );
NOR2_X2 _sha1_round_add_79_U228  ( .A1(_sha1_round_add_79_n214 ), .A2(_sha1_round_add_79_n215 ), .ZN(_sha1_round_add_79_n210 ) );
NOR2_X2 _sha1_round_add_79_U227  ( .A1(_sha1_round_add_79_n158 ), .A2(_sha1_round_add_79_n159 ), .ZN(_sha1_round_add_79_n155 ) );
NAND3_X2 _sha1_round_add_79_U226  ( .A1(_sha1_round_add_79_n155 ), .A2(_sha1_round_add_79_n156 ), .A3(_sha1_round_add_79_n157 ), .ZN(_sha1_round_add_79_n153 ) );
NOR2_X2 _sha1_round_add_79_U225  ( .A1(_sha1_round_add_79_n177 ), .A2(_sha1_round_add_79_n178 ), .ZN(_sha1_round_add_79_n172 ) );
NAND3_X2 _sha1_round_add_79_U224  ( .A1(_sha1_round_add_79_n172 ), .A2(_sha1_round_add_79_n173 ), .A3(_sha1_round_add_79_n174 ), .ZN(_sha1_round_add_79_n170 ) );
NOR2_X2 _sha1_round_add_79_U223  ( .A1(_sha1_round_add_79_n308 ), .A2(_sha1_round_add_79_n129 ), .ZN(_sha1_round_add_79_n367 ) );
INV_X1 _sha1_round_add_79_U222  ( .A(_sha1_round_n512 ), .ZN(_sha1_round_add_79_n90 ) );
XNOR2_X2 _sha1_round_add_79_U221  ( .A(_sha1_round_add_79_n245 ), .B(_sha1_round_add_79_n246 ), .ZN(_sha1_round_N274 ) );
NAND3_X2 _sha1_round_add_79_U220  ( .A1(_sha1_round_add_79_n235 ), .A2(_sha1_round_add_79_n297 ), .A3(_sha1_round_add_79_n236 ), .ZN(_sha1_round_add_79_n287 ) );
NOR2_X1 _sha1_round_add_79_U219  ( .A1(_sha1_round_add_79_n185 ), .A2(_sha1_round_add_79_n146 ), .ZN(_sha1_round_add_79_n181 ) );
NOR2_X2 _sha1_round_add_79_U218  ( .A1(_sha1_round_add_79_n160 ), .A2(_sha1_round_add_79_n164 ), .ZN(_sha1_round_add_79_n151 ) );
INV_X4 _sha1_round_add_79_U217  ( .A(_sha1_round_add_79_n90 ), .ZN(_sha1_round_add_79_n89 ) );
NAND2_X4 _sha1_round_add_79_U216  ( .A1(_sha1_round_add_79_n362 ), .A2(_sha1_round_add_79_n90 ), .ZN(_sha1_round_add_79_n359 ) );
INV_X1 _sha1_round_add_79_U215  ( .A(_sha1_round_add_79_n270 ), .ZN(_sha1_round_add_79_n381 ) );
OR2_X4 _sha1_round_add_79_U214  ( .A1(_sha1_round_n825 ), .A2(_sha1_round_f [29]), .ZN(_sha1_round_add_79_n165 ) );
OR2_X4 _sha1_round_add_79_U213  ( .A1(_sha1_round_k_30 ), .A2(_sha1_round_f [30]), .ZN(_sha1_round_add_79_n149 ) );
NOR2_X2 _sha1_round_add_79_U212  ( .A1(_sha1_round_add_79_n309 ), .A2(_sha1_round_add_79_n108 ), .ZN(_sha1_round_add_79_n304 ) );
OR2_X4 _sha1_round_add_79_U211  ( .A1(_sha1_round_n824 ), .A2(_sha1_round_f [21]), .ZN(_sha1_round_add_79_n240 ) );
NOR2_X2 _sha1_round_add_79_U210  ( .A1(_sha1_round_add_79_n181 ), .A2(_sha1_round_add_79_n182 ), .ZN(_sha1_round_add_79_n64 ) );
XOR2_X2 _sha1_round_add_79_U209  ( .A(_sha1_round_add_79_n64 ), .B(_sha1_round_add_79_n179 ), .Z(_sha1_round_N280 ) );
AND2_X4 _sha1_round_add_79_U208  ( .A1(_sha1_round_add_79_n244 ), .A2(_sha1_round_add_79_n241 ), .ZN(_sha1_round_add_79_n74 ) );
INV_X1 _sha1_round_add_79_U207  ( .A(_sha1_round_add_79_n308 ), .ZN(_sha1_round_add_79_n307 ) );
NAND3_X1 _sha1_round_add_79_U206  ( .A1(_sha1_round_add_79_n198 ), .A2(_sha1_round_add_79_n196 ), .A3(_sha1_round_add_79_n197 ), .ZN(_sha1_round_add_79_n206 ) );
NOR2_X2 _sha1_round_add_79_U205  ( .A1(_sha1_round_add_79_n12 ), .A2(_sha1_round_add_79_n238 ), .ZN(_sha1_round_add_79_n277 ) );
NAND4_X1 _sha1_round_add_79_U204  ( .A1(_sha1_round_add_79_n223 ), .A2(_sha1_round_add_79_n224 ), .A3(_sha1_round_add_79_n225 ), .A4(_sha1_round_add_79_n226 ), .ZN(_sha1_round_add_79_n221 ) );
NOR2_X1 _sha1_round_add_79_U203  ( .A1(_sha1_round_add_79_n79 ), .A2(_sha1_round_add_79_n278 ), .ZN(_sha1_round_add_79_n231 ) );
OR2_X4 _sha1_round_add_79_U202  ( .A1(_sha1_round_add_79_n168 ), .A2(_sha1_round_add_79_n270 ), .ZN(_sha1_round_add_79_n68 ) );
NOR2_X1 _sha1_round_add_79_U201  ( .A1(_sha1_round_add_79_n380 ), .A2(_sha1_round_add_79_n119 ), .ZN(_sha1_round_add_79_n118 ) );
NOR2_X1 _sha1_round_add_79_U200  ( .A1(_sha1_round_add_79_n347 ), .A2(_sha1_round_add_79_n345 ), .ZN(_sha1_round_add_79_n353 ) );
NAND3_X2 _sha1_round_add_79_U199  ( .A1(_sha1_round_add_79_n277 ), .A2(_sha1_round_add_79_n235 ), .A3(_sha1_round_add_79_n236 ), .ZN(_sha1_round_add_79_n276 ) );
INV_X1 _sha1_round_add_79_U198  ( .A(_sha1_round_n517 ), .ZN(_sha1_round_add_79_n92 ) );
NOR2_X1 _sha1_round_add_79_U197  ( .A1(_sha1_round_f [24]), .A2(_sha1_round_add_79_n89 ), .ZN(_sha1_round_add_79_n212 ) );
NAND3_X2 _sha1_round_add_79_U196  ( .A1(_sha1_round_add_79_n313 ), .A2(_sha1_round_add_79_n314 ), .A3(_sha1_round_add_79_n315 ), .ZN(_sha1_round_add_79_n238 ) );
INV_X4 _sha1_round_add_79_U195  ( .A(_sha1_round_add_79_n60 ), .ZN(_sha1_round_add_79_n61 ) );
NAND2_X2 _sha1_round_add_79_U194  ( .A1(_sha1_round_add_79_n13 ), .A2(_sha1_round_add_79_n319 ), .ZN(_sha1_round_add_79_n235 ) );
INV_X1 _sha1_round_add_79_U193  ( .A(_sha1_round_add_79_n317 ), .ZN(_sha1_round_add_79_n327 ) );
NOR2_X1 _sha1_round_add_79_U192  ( .A1(_sha1_round_add_79_n185 ), .A2(_sha1_round_add_79_n187 ), .ZN(_sha1_round_add_79_n190 ) );
NAND2_X1 _sha1_round_add_79_U191  ( .A1(_sha1_round_add_79_n233 ), .A2(_sha1_round_add_79_n280 ), .ZN(_sha1_round_add_79_n291 ) );
INV_X2 _sha1_round_add_79_U190  ( .A(_sha1_round_add_79_n291 ), .ZN(_sha1_round_add_79_n57 ) );
INV_X4 _sha1_round_add_79_U189  ( .A(_sha1_round_add_79_n290 ), .ZN(_sha1_round_add_79_n56 ) );
NAND2_X4 _sha1_round_add_79_U188  ( .A1(_sha1_round_add_79_n58 ), .A2(_sha1_round_add_79_n59 ), .ZN(_sha1_round_N268 ) );
NAND2_X4 _sha1_round_add_79_U187  ( .A1(_sha1_round_add_79_n56 ), .A2(_sha1_round_add_79_n57 ), .ZN(_sha1_round_add_79_n59 ) );
NAND2_X2 _sha1_round_add_79_U186  ( .A1(_sha1_round_add_79_n291 ), .A2(_sha1_round_add_79_n290 ), .ZN(_sha1_round_add_79_n58 ) );
NAND2_X4 _sha1_round_add_79_U185  ( .A1(_sha1_round_add_79_n322 ), .A2(_sha1_round_add_79_n294 ), .ZN(_sha1_round_add_79_n320 ) );
NAND3_X2 _sha1_round_add_79_U184  ( .A1(_sha1_round_add_79_n104 ), .A2(_sha1_round_add_79_n298 ), .A3(_sha1_round_add_79_n299 ), .ZN(_sha1_round_add_79_n236 ) );
NAND2_X1 _sha1_round_add_79_U183  ( .A1(_sha1_round_n517 ), .A2(_sha1_round_f [3]), .ZN(_sha1_round_add_79_n306 ) );
NAND2_X1 _sha1_round_add_79_U182  ( .A1(_sha1_round_add_79_n87 ), .A2(_sha1_round_f [2]), .ZN(_sha1_round_add_79_n311 ) );
NOR2_X4 _sha1_round_add_79_U181  ( .A1(_sha1_round_f [5]), .A2(_sha1_round_n825 ), .ZN(_sha1_round_add_79_n380 ) );
NAND2_X2 _sha1_round_add_79_U180  ( .A1(_sha1_round_add_79_n4 ), .A2(_sha1_round_add_79_n101 ), .ZN(_sha1_round_add_79_n364 ) );
XNOR2_X2 _sha1_round_add_79_U179  ( .A(_sha1_round_add_79_n325 ), .B(_sha1_round_add_79_n326 ), .ZN(_sha1_round_N266 ) );
NOR2_X4 _sha1_round_add_79_U178  ( .A1(_sha1_round_f [9]), .A2(_sha1_round_n825 ), .ZN(_sha1_round_add_79_n349 ) );
NAND2_X1 _sha1_round_add_79_U177  ( .A1(_sha1_round_f [9]), .A2(_sha1_round_n825 ), .ZN(_sha1_round_add_79_n96 ) );
NAND3_X2 _sha1_round_add_79_U176  ( .A1(_sha1_round_add_79_n33 ), .A2(_sha1_round_add_79_n85 ), .A3(_sha1_round_n825 ), .ZN(_sha1_round_add_79_n374 ) );
NOR2_X2 _sha1_round_add_79_U175  ( .A1(_sha1_round_add_79_n115 ), .A2(_sha1_round_add_79_n379 ), .ZN(_sha1_round_add_79_n114 ) );
OR2_X4 _sha1_round_add_79_U174  ( .A1(_sha1_round_add_79_n84 ), .A2(_sha1_round_add_79_n312 ), .ZN(_sha1_round_add_79_n78 ) );
NAND2_X4 _sha1_round_add_79_U173  ( .A1(_sha1_round_add_79_n53 ), .A2(_sha1_round_add_79_n54 ), .ZN(_sha1_round_N267 ) );
NAND2_X4 _sha1_round_add_79_U172  ( .A1(_sha1_round_add_79_n51 ), .A2(_sha1_round_add_79_n52 ), .ZN(_sha1_round_add_79_n54 ) );
INV_X4 _sha1_round_add_79_U171  ( .A(_sha1_round_add_79_n49 ), .ZN(_sha1_round_add_79_n50 ) );
NAND2_X4 _sha1_round_add_79_U170  ( .A1(_sha1_round_add_79_n50 ), .A2(_sha1_round_add_79_n226 ), .ZN(_sha1_round_add_79_n145 ) );
NAND2_X4 _sha1_round_add_79_U169  ( .A1(_sha1_round_add_79_n23 ), .A2(_sha1_round_add_79_n35 ), .ZN(_sha1_round_add_79_n303 ) );
NAND2_X4 _sha1_round_add_79_U168  ( .A1(_sha1_round_add_79_n61 ), .A2(_sha1_round_add_79_n63 ), .ZN(_sha1_round_add_79_n101 ) );
NAND2_X4 _sha1_round_add_79_U167  ( .A1(_sha1_round_add_79_n48 ), .A2(_sha1_round_add_79_n47 ), .ZN(_sha1_round_N259 ) );
NAND2_X4 _sha1_round_add_79_U166  ( .A1(_sha1_round_add_79_n45 ), .A2(_sha1_round_add_79_n46 ), .ZN(_sha1_round_add_79_n48 ) );
INV_X2 _sha1_round_add_79_U165  ( .A(_sha1_round_add_79_n361 ), .ZN(_sha1_round_add_79_n42 ) );
NAND2_X4 _sha1_round_add_79_U164  ( .A1(_sha1_round_add_79_n43 ), .A2(_sha1_round_add_79_n44 ), .ZN(_sha1_round_N262 ) );
NAND2_X4 _sha1_round_add_79_U163  ( .A1(_sha1_round_add_79_n41 ), .A2(_sha1_round_add_79_n42 ), .ZN(_sha1_round_add_79_n44 ) );
NOR2_X2 _sha1_round_add_79_U162  ( .A1(_sha1_round_add_79_n239 ), .A2(_sha1_round_add_79_n79 ), .ZN(_sha1_round_add_79_n283 ) );
INV_X4 _sha1_round_add_79_U161  ( .A(_sha1_round_add_79_n283 ), .ZN(_sha1_round_add_79_n38 ) );
NAND2_X4 _sha1_round_add_79_U160  ( .A1(_sha1_round_add_79_n39 ), .A2(_sha1_round_add_79_n40 ), .ZN(_sha1_round_add_79_n281 ) );
NAND2_X4 _sha1_round_add_79_U159  ( .A1(_sha1_round_add_79_n37 ), .A2(_sha1_round_add_79_n38 ), .ZN(_sha1_round_add_79_n40 ) );
NAND2_X2 _sha1_round_add_79_U158  ( .A1(_sha1_round_add_79_n282 ), .A2(_sha1_round_add_79_n283 ), .ZN(_sha1_round_add_79_n39 ) );
INV_X2 _sha1_round_add_79_U157  ( .A(_sha1_round_add_79_n348 ), .ZN(_sha1_round_add_79_n366 ) );
NAND2_X2 _sha1_round_add_79_U156  ( .A1(_sha1_round_f [1]), .A2(_sha1_round_n824 ), .ZN(_sha1_round_add_79_n370 ) );
NAND2_X2 _sha1_round_add_79_U155  ( .A1(_sha1_round_n824 ), .A2(_sha1_round_f [1]), .ZN(_sha1_round_add_79_n167 ) );
NAND2_X1 _sha1_round_add_79_U154  ( .A1(_sha1_round_f [13]), .A2(_sha1_round_k[13] ), .ZN(_sha1_round_add_79_n323 ) );
NAND2_X4 _sha1_round_add_79_U153  ( .A1(_sha1_round_add_79_n109 ), .A2(_sha1_round_add_79_n21 ), .ZN(_sha1_round_add_79_n99 ) );
NAND3_X2 _sha1_round_add_79_U152  ( .A1(_sha1_round_add_79_n36 ), .A2(_sha1_round_add_79_n344 ), .A3(_sha1_round_add_79_n343 ), .ZN(_sha1_round_add_79_n35 ) );
NOR3_X2 _sha1_round_add_79_U151  ( .A1(_sha1_round_add_79_n78 ), .A2(_sha1_round_add_79_n132 ), .A3(_sha1_round_add_79_n168 ), .ZN(_sha1_round_add_79_n369 ) );
NAND3_X2 _sha1_round_add_79_U150  ( .A1(_sha1_round_add_79_n101 ), .A2(_sha1_round_add_79_n99 ), .A3(_sha1_round_add_79_n14 ), .ZN(_sha1_round_add_79_n358 ) );
INV_X1 _sha1_round_add_79_U149  ( .A(_sha1_round_add_79_n82 ), .ZN(_sha1_round_add_79_n256 ) );
INV_X2 _sha1_round_add_79_U148  ( .A(_sha1_round_add_79_n132 ), .ZN(_sha1_round_add_79_n169 ) );
NAND2_X2 _sha1_round_add_79_U147  ( .A1(_sha1_round_add_79_n112 ), .A2(_sha1_round_add_79_n113 ), .ZN(_sha1_round_add_79_n47 ) );
INV_X4 _sha1_round_add_79_U146  ( .A(_sha1_round_add_79_n113 ), .ZN(_sha1_round_add_79_n46 ) );
NOR2_X2 _sha1_round_add_79_U145  ( .A1(_sha1_round_add_79_n111 ), .A2(_sha1_round_add_79_n83 ), .ZN(_sha1_round_add_79_n113 ) );
INV_X2 _sha1_round_add_79_U144  ( .A(_sha1_round_add_79_n111 ), .ZN(_sha1_round_add_79_n110 ) );
OR2_X4 _sha1_round_add_79_U143  ( .A1(_sha1_round_k[15] ), .A2(_sha1_round_f [15]), .ZN(_sha1_round_add_79_n289 ) );
NAND2_X1 _sha1_round_add_79_U142  ( .A1(_sha1_round_add_79_n295 ), .A2(_sha1_round_add_79_n289 ), .ZN(_sha1_round_add_79_n321 ) );
NOR2_X1 _sha1_round_add_79_U141  ( .A1(_sha1_round_add_79_n269 ), .A2(_sha1_round_add_79_n168 ), .ZN(_sha1_round_add_79_n268 ) );
INV_X2 _sha1_round_add_79_U140  ( .A(_sha1_round_n3170 ), .ZN(_sha1_round_add_79_n86 ) );
NAND2_X1 _sha1_round_add_79_U139  ( .A1(_sha1_round_f [21]), .A2(_sha1_round_n824 ), .ZN(_sha1_round_add_79_n252 ) );
NOR2_X4 _sha1_round_add_79_U138  ( .A1(_sha1_round_add_79_n300 ), .A2(_sha1_round_add_79_n301 ), .ZN(_sha1_round_add_79_n299 ) );
INV_X4 _sha1_round_add_79_U137  ( .A(_sha1_round_add_79_n324 ), .ZN(_sha1_round_add_79_n328 ) );
INV_X4 _sha1_round_add_79_U136  ( .A(_sha1_round_add_79_n282 ), .ZN(_sha1_round_add_79_n37 ) );
NAND2_X4 _sha1_round_add_79_U135  ( .A1(_sha1_round_f [11]), .A2(_sha1_round_k[13] ), .ZN(_sha1_round_add_79_n343 ) );
NOR2_X2 _sha1_round_add_79_U134  ( .A1(_sha1_round_add_79_n260 ), .A2(_sha1_round_add_79_n251 ), .ZN(_sha1_round_add_79_n255 ) );
INV_X4 _sha1_round_add_79_U133  ( .A(_sha1_round_add_79_n250 ), .ZN(_sha1_round_add_79_n260 ) );
NAND2_X4 _sha1_round_add_79_U132  ( .A1(_sha1_round_f [10]), .A2(_sha1_round_add_79_n89 ), .ZN(_sha1_round_add_79_n344 ) );
NOR2_X4 _sha1_round_add_79_U131  ( .A1(_sha1_round_add_79_n117 ), .A2(_sha1_round_add_79_n18 ), .ZN(_sha1_round_add_79_n115 ) );
NAND2_X1 _sha1_round_add_79_U130  ( .A1(_sha1_round_add_79_n311 ), .A2(_sha1_round_add_79_n312 ), .ZN(_sha1_round_add_79_n310 ) );
OR2_X4 _sha1_round_add_79_U129  ( .A1(_sha1_round_add_79_n261 ), .A2(_sha1_round_add_79_n272 ), .ZN(_sha1_round_add_79_n34 ) );
XNOR2_X2 _sha1_round_add_79_U128  ( .A(_sha1_round_add_79_n273 ), .B(_sha1_round_add_79_n34 ), .ZN(_sha1_round_N271 ) );
NOR2_X1 _sha1_round_add_79_U127  ( .A1(_sha1_round_add_79_n80 ), .A2(_sha1_round_add_79_n380 ), .ZN(_sha1_round_add_79_n124 ) );
INV_X2 _sha1_round_add_79_U126  ( .A(_sha1_round_add_79_n359 ), .ZN(_sha1_round_add_79_n346 ) );
NAND2_X2 _sha1_round_add_79_U125  ( .A1(_sha1_round_add_79_n365 ), .A2(_sha1_round_add_79_n359 ), .ZN(_sha1_round_add_79_n36 ) );
INV_X1 _sha1_round_add_79_U124  ( .A(_sha1_round_add_79_n244 ), .ZN(_sha1_round_add_79_n248 ) );
NAND2_X4 _sha1_round_add_79_U123  ( .A1(_sha1_round_add_79_n68 ), .A2(_sha1_round_add_79_n167 ), .ZN(_sha1_round_add_79_n134 ) );
NAND2_X2 _sha1_round_add_79_U122  ( .A1(_sha1_round_n825 ), .A2(_sha1_round_f [9]), .ZN(_sha1_round_add_79_n342 ) );
NAND2_X2 _sha1_round_add_79_U121  ( .A1(_sha1_round_add_79_n336 ), .A2(_sha1_round_add_79_n313 ), .ZN(_sha1_round_add_79_n335 ) );
INV_X4 _sha1_round_add_79_U120  ( .A(_sha1_round_add_79_n32 ), .ZN(_sha1_round_add_79_n33 ) );
INV_X1 _sha1_round_add_79_U119  ( .A(_sha1_round_f [5]), .ZN(_sha1_round_add_79_n32 ) );
NAND2_X1 _sha1_round_add_79_U118  ( .A1(_sha1_round_f [23]), .A2(_sha1_round_k_23 ), .ZN(_sha1_round_add_79_n219 ) );
NAND2_X1 _sha1_round_add_79_U117  ( .A1(_sha1_round_f [16]), .A2(_sha1_round_k_26 ), .ZN(_sha1_round_add_79_n233 ) );
NAND2_X1 _sha1_round_add_79_U116  ( .A1(_sha1_round_f [19]), .A2(_sha1_round_k_26 ), .ZN(_sha1_round_add_79_n266 ) );
NAND2_X1 _sha1_round_add_79_U115  ( .A1(_sha1_round_k_30 ), .A2(_sha1_round_f [8]), .ZN(_sha1_round_add_79_n100 ) );
OR2_X2 _sha1_round_add_79_U114  ( .A1(_sha1_round_f [6]), .A2(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n85 ) );
OR3_X1 _sha1_round_add_79_U113  ( .A1(_sha1_round_add_79_n132 ), .A2(_sha1_round_add_79_n26 ), .A3(_sha1_round_add_79_n168 ), .ZN(_sha1_round_add_79_n70 ) );
NAND2_X2 _sha1_round_add_79_U112  ( .A1(_sha1_round_add_79_n203 ), .A2(_sha1_round_add_79_n204 ), .ZN(_sha1_round_add_79_n199 ) );
XNOR2_X1 _sha1_round_add_79_U111  ( .A(_sha1_round_add_79_n228 ), .B(_sha1_round_add_79_n145 ), .ZN(_sha1_round_N275 ) );
NOR3_X2 _sha1_round_add_79_U110  ( .A1(_sha1_round_add_79_n349 ), .A2(_sha1_round_add_79_n348 ), .A3(_sha1_round_add_79_n71 ), .ZN(_sha1_round_add_79_n31 ) );
NAND2_X4 _sha1_round_add_79_U109  ( .A1(_sha1_round_add_79_n210 ), .A2(_sha1_round_add_79_n211 ), .ZN(_sha1_round_add_79_n207 ) );
NAND2_X2 _sha1_round_add_79_U108  ( .A1(_sha1_round_f [12]), .A2(_sha1_round_n3300 ), .ZN(_sha1_round_add_79_n302 ) );
INV_X4 _sha1_round_add_79_U107  ( .A(_sha1_round_add_79_n112 ), .ZN(_sha1_round_add_79_n45 ) );
NOR2_X2 _sha1_round_add_79_U106  ( .A1(_sha1_round_add_79_n255 ), .A2(_sha1_round_add_79_n256 ), .ZN(_sha1_round_add_79_n254 ) );
NAND2_X2 _sha1_round_add_79_U105  ( .A1(_sha1_round_add_79_n69 ), .A2(_sha1_round_add_79_n252 ), .ZN(_sha1_round_add_79_n244 ) );
AND2_X2 _sha1_round_add_79_U104  ( .A1(_sha1_round_add_79_n252 ), .A2(_sha1_round_add_79_n243 ), .ZN(_sha1_round_add_79_n30 ) );
OR2_X2 _sha1_round_add_79_U103  ( .A1(_sha1_round_add_79_n227 ), .A2(_sha1_round_add_79_n241 ), .ZN(_sha1_round_add_79_n29 ) );
NAND2_X2 _sha1_round_add_79_U102  ( .A1(_sha1_round_add_79_n28 ), .A2(_sha1_round_add_79_n29 ), .ZN(_sha1_round_add_79_n229 ) );
NAND2_X2 _sha1_round_add_79_U101  ( .A1(_sha1_round_add_79_n69 ), .A2(_sha1_round_add_79_n30 ), .ZN(_sha1_round_add_79_n28 ) );
INV_X1 _sha1_round_add_79_U100  ( .A(_sha1_round_add_79_n27 ), .ZN(_sha1_round_add_79_n261 ) );
NOR2_X2 _sha1_round_add_79_U99  ( .A1(_sha1_round_add_79_n262 ), .A2(_sha1_round_add_79_n260 ), .ZN(_sha1_round_add_79_n273 ) );
NAND2_X2 _sha1_round_add_79_U98  ( .A1(_sha1_round_n2 ), .A2(_sha1_round_f [4]), .ZN(_sha1_round_add_79_n378 ) );
INV_X4 _sha1_round_add_79_U97  ( .A(_sha1_round_add_79_n320 ), .ZN(_sha1_round_add_79_n51 ) );
INV_X2 _sha1_round_add_79_U96  ( .A(_sha1_round_f [10]), .ZN(_sha1_round_add_79_n362 ) );
NAND2_X2 _sha1_round_add_79_U95  ( .A1(_sha1_round_add_79_n360 ), .A2(_sha1_round_add_79_n361 ), .ZN(_sha1_round_add_79_n43 ) );
NAND2_X2 _sha1_round_add_79_U94  ( .A1(_sha1_round_add_79_n99 ), .A2(_sha1_round_add_79_n100 ), .ZN(_sha1_round_add_79_n98 ) );
NOR2_X4 _sha1_round_add_79_U93  ( .A1(_sha1_round_add_79_n97 ), .A2(_sha1_round_add_79_n98 ), .ZN(_sha1_round_add_79_n93 ) );
NAND2_X2 _sha1_round_add_79_U92  ( .A1(_sha1_round_add_79_n325 ), .A2(_sha1_round_add_79_n327 ), .ZN(_sha1_round_add_79_n322 ) );
NAND2_X2 _sha1_round_add_79_U91  ( .A1(_sha1_round_add_79_n320 ), .A2(_sha1_round_add_79_n321 ), .ZN(_sha1_round_add_79_n53 ) );
NOR2_X2 _sha1_round_add_79_U90  ( .A1(_sha1_round_add_79_n316 ), .A2(_sha1_round_add_79_n317 ), .ZN(_sha1_round_add_79_n315 ) );
NOR2_X2 _sha1_round_add_79_U89  ( .A1(_sha1_round_n517 ), .A2(_sha1_round_f [3]), .ZN(_sha1_round_add_79_n26 ) );
OR2_X4 _sha1_round_add_79_U88  ( .A1(_sha1_round_f [24]), .A2(_sha1_round_add_79_n89 ), .ZN(_sha1_round_add_79_n25 ) );
AND2_X4 _sha1_round_add_79_U87  ( .A1(_sha1_round_add_79_n340 ), .A2(_sha1_round_add_79_n339 ), .ZN(_sha1_round_add_79_n23 ) );
AND2_X4 _sha1_round_add_79_U86  ( .A1(_sha1_round_add_79_n152 ), .A2(_sha1_round_add_79_n184 ), .ZN(_sha1_round_add_79_n22 ) );
AND2_X4 _sha1_round_add_79_U85  ( .A1(_sha1_round_add_79_n366 ), .A2(_sha1_round_add_79_n110 ), .ZN(_sha1_round_add_79_n21 ) );
OR2_X4 _sha1_round_add_79_U84  ( .A1(_sha1_round_add_79_n334 ), .A2(_sha1_round_add_79_n318 ), .ZN(_sha1_round_add_79_n20 ) );
OR2_X4 _sha1_round_add_79_U83  ( .A1(_sha1_round_add_79_n318 ), .A2(_sha1_round_add_79_n302 ), .ZN(_sha1_round_add_79_n19 ) );
OR2_X4 _sha1_round_add_79_U82  ( .A1(_sha1_round_add_79_n118 ), .A2(_sha1_round_add_79_n80 ), .ZN(_sha1_round_add_79_n18 ) );
OR2_X4 _sha1_round_add_79_U81  ( .A1(_sha1_round_add_79_n26 ), .A2(_sha1_round_add_79_n370 ), .ZN(_sha1_round_add_79_n17 ) );
OR2_X4 _sha1_round_add_79_U80  ( .A1(_sha1_round_add_79_n318 ), .A2(_sha1_round_add_79_n330 ), .ZN(_sha1_round_add_79_n16 ) );
AND2_X4 _sha1_round_add_79_U79  ( .A1(_sha1_round_add_79_n252 ), .A2(_sha1_round_add_79_n240 ), .ZN(_sha1_round_add_79_n15 ) );
AND2_X4 _sha1_round_add_79_U78  ( .A1(_sha1_round_add_79_n96 ), .A2(_sha1_round_add_79_n100 ), .ZN(_sha1_round_add_79_n14 ) );
OR2_X2 _sha1_round_add_79_U77  ( .A1(_sha1_round_add_79_n79 ), .A2(_sha1_round_add_79_n278 ), .ZN(_sha1_round_add_79_n12 ) );
AND2_X4 _sha1_round_add_79_U76  ( .A1(_sha1_round_add_79_n323 ), .A2(_sha1_round_add_79_n19 ), .ZN(_sha1_round_add_79_n11 ) );
INV_X1 _sha1_round_add_79_U75  ( .A(_sha1_round_k_27 ), .ZN(_sha1_round_add_79_n55 ) );
OR2_X4 _sha1_round_add_79_U74  ( .A1(_sha1_round_f [4]), .A2(_sha1_round_n2 ), .ZN(_sha1_round_add_79_n8 ) );
NAND2_X1 _sha1_round_add_79_U73  ( .A1(_sha1_round_add_79_n119 ), .A2(_sha1_round_add_79_n8 ), .ZN(_sha1_round_add_79_n126 ) );
NAND2_X1 _sha1_round_add_79_U72  ( .A1(_sha1_round_f [2]), .A2(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n371 ) );
NOR2_X2 _sha1_round_add_79_U71  ( .A1(_sha1_round_add_79_n26 ), .A2(_sha1_round_add_79_n371 ), .ZN(_sha1_round_add_79_n308 ) );
AND2_X2 _sha1_round_add_79_U70  ( .A1(_sha1_round_add_79_n302 ), .A2(_sha1_round_add_79_n303 ), .ZN(_sha1_round_add_79_n13 ) );
NAND2_X1 _sha1_round_add_79_U69  ( .A1(_sha1_round_add_79_n332 ), .A2(_sha1_round_add_79_n303 ), .ZN(_sha1_round_add_79_n331 ) );
NOR2_X2 _sha1_round_add_79_U68  ( .A1(_sha1_round_add_79_n67 ), .A2(_sha1_round_add_79_n331 ), .ZN(_sha1_round_add_79_n329 ) );
NAND2_X1 _sha1_round_add_79_U67  ( .A1(_sha1_round_f [14]), .A2(_sha1_round_k_30 ), .ZN(_sha1_round_add_79_n294 ) );
NOR2_X1 _sha1_round_add_79_U66  ( .A1(_sha1_round_add_79_n95 ), .A2(_sha1_round_add_79_n349 ), .ZN(_sha1_round_add_79_n94 ) );
INV_X1 _sha1_round_add_79_U65  ( .A(_sha1_round_add_79_n145 ), .ZN(_sha1_round_add_79_n185 ) );
NAND2_X1 _sha1_round_add_79_U64  ( .A1(_sha1_round_add_79_n106 ), .A2(_sha1_round_add_79_n107 ), .ZN(_sha1_round_add_79_n105 ) );
NOR2_X2 _sha1_round_add_79_U63  ( .A1(_sha1_round_add_79_n329 ), .A2(_sha1_round_add_79_n16 ), .ZN(_sha1_round_add_79_n324 ) );
NOR2_X2 _sha1_round_add_79_U62  ( .A1(_sha1_round_f [14]), .A2(_sha1_round_k_30 ), .ZN(_sha1_round_add_79_n317 ) );
NAND2_X2 _sha1_round_add_79_U61  ( .A1(_sha1_round_k_26 ), .A2(_sha1_round_f [20]), .ZN(_sha1_round_add_79_n258 ) );
NAND2_X2 _sha1_round_add_79_U60  ( .A1(_sha1_round_add_79_n109 ), .A2(_sha1_round_add_79_n110 ), .ZN(_sha1_round_add_79_n104 ) );
NOR2_X2 _sha1_round_add_79_U59  ( .A1(_sha1_round_f [1]), .A2(_sha1_round_n824 ), .ZN(_sha1_round_add_79_n168 ) );
NAND2_X2 _sha1_round_add_79_U58  ( .A1(_sha1_round_add_79_n293 ), .A2(_sha1_round_add_79_n233 ), .ZN(_sha1_round_add_79_n232 ) );
NAND2_X2 _sha1_round_add_79_U57  ( .A1(_sha1_round_add_79_n239 ), .A2(_sha1_round_add_79_n230 ), .ZN(_sha1_round_add_79_n224 ) );
NOR2_X2 _sha1_round_add_79_U56  ( .A1(_sha1_round_add_79_n190 ), .A2(_sha1_round_add_79_n183 ), .ZN(_sha1_round_add_79_n188 ) );
NAND3_X2 _sha1_round_add_79_U55  ( .A1(_sha1_round_f [18]), .A2(_sha1_round_add_79_n259 ), .A3(_sha1_round_add_79_n27 ), .ZN(_sha1_round_add_79_n251 ) );
INV_X4 _sha1_round_add_79_U54  ( .A(_sha1_round_add_79_n360 ), .ZN(_sha1_round_add_79_n41 ) );
NAND2_X2 _sha1_round_add_79_U53  ( .A1(_sha1_round_add_79_n364 ), .A2(_sha1_round_add_79_n365 ), .ZN(_sha1_round_add_79_n363 ) );
NOR2_X2 _sha1_round_add_79_U52  ( .A1(_sha1_round_add_79_n132 ), .A2(_sha1_round_add_79_n133 ), .ZN(_sha1_round_add_79_n130 ) );
NOR2_X2 _sha1_round_add_79_U51  ( .A1(_sha1_round_add_79_n130 ), .A2(_sha1_round_add_79_n131 ), .ZN(_sha1_round_add_79_n127 ) );
INV_X4 _sha1_round_add_79_U50  ( .A(_sha1_round_add_79_n349 ), .ZN(_sha1_round_add_79_n365 ) );
NOR2_X2 _sha1_round_add_79_U49  ( .A1(_sha1_round_f [7]), .A2(_sha1_round_k_27 ), .ZN(_sha1_round_add_79_n373 ) );
NAND3_X2 _sha1_round_add_79_U48  ( .A1(_sha1_round_add_79_n372 ), .A2(_sha1_round_add_79_n8 ), .A3(_sha1_round_add_79_n121 ), .ZN(_sha1_round_add_79_n108 ) );
NOR2_X2 _sha1_round_add_79_U47  ( .A1(_sha1_round_add_79_n379 ), .A2(_sha1_round_add_79_n373 ), .ZN(_sha1_round_add_79_n372 ) );
NOR2_X1 _sha1_round_add_79_U46  ( .A1(_sha1_round_add_79_n81 ), .A2(_sha1_round_add_79_n379 ), .ZN(_sha1_round_add_79_n116 ) );
INV_X4 _sha1_round_add_79_U45  ( .A(_sha1_round_add_79_n108 ), .ZN(_sha1_round_add_79_n106 ) );
NOR2_X4 _sha1_round_add_79_U44  ( .A1(_sha1_round_f [6]), .A2(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n379 ) );
INV_X2 _sha1_round_add_79_U43  ( .A(_sha1_round_add_79_n287 ), .ZN(_sha1_round_add_79_n286 ) );
NAND2_X1 _sha1_round_add_79_U42  ( .A1(_sha1_round_add_79_n287 ), .A2(_sha1_round_add_79_n293 ), .ZN(_sha1_round_add_79_n290 ) );
NOR2_X1 _sha1_round_add_79_U41  ( .A1(_sha1_round_n517 ), .A2(_sha1_round_f [3]), .ZN(_sha1_round_add_79_n84 ) );
NAND2_X4 _sha1_round_add_79_U40  ( .A1(_sha1_round_add_79_n285 ), .A2(_sha1_round_add_79_n284 ), .ZN(_sha1_round_add_79_n282 ) );
NAND2_X4 _sha1_round_add_79_U39  ( .A1(_sha1_round_add_79_n5 ), .A2(_sha1_round_add_79_n338 ), .ZN(_sha1_round_add_79_n336 ) );
NAND3_X4 _sha1_round_add_79_U38  ( .A1(_sha1_round_add_79_n240 ), .A2(_sha1_round_add_79_n241 ), .A3(_sha1_round_add_79_n242 ), .ZN(_sha1_round_add_79_n237 ) );
NOR3_X4 _sha1_round_add_79_U37  ( .A1(_sha1_round_add_79_n237 ), .A2(_sha1_round_add_79_n12 ), .A3(_sha1_round_add_79_n238 ), .ZN(_sha1_round_add_79_n234 ) );
NAND2_X1 _sha1_round_add_79_U36  ( .A1(_sha1_round_f [27]), .A2(_sha1_round_k_27 ), .ZN(_sha1_round_add_79_n152 ) );
NAND2_X1 _sha1_round_add_79_U35  ( .A1(_sha1_round_f [25]), .A2(_sha1_round_k_27 ), .ZN(_sha1_round_add_79_n198 ) );
OR2_X2 _sha1_round_add_79_U34  ( .A1(_sha1_round_add_79_n317 ), .A2(_sha1_round_add_79_n296 ), .ZN(_sha1_round_add_79_n24 ) );
NOR2_X1 _sha1_round_add_79_U33  ( .A1(_sha1_round_f [13]), .A2(_sha1_round_k[13] ), .ZN(_sha1_round_add_79_n318 ) );
OR2_X4 _sha1_round_add_79_U32  ( .A1(_sha1_round_f [19]), .A2(_sha1_round_k_26 ), .ZN(_sha1_round_add_79_n27 ) );
INV_X1 _sha1_round_add_79_U31  ( .A(_sha1_round_add_79_n340 ), .ZN(_sha1_round_add_79_n347 ) );
NAND2_X2 _sha1_round_add_79_U30  ( .A1(_sha1_round_add_79_n286 ), .A2(_sha1_round_add_79_n280 ), .ZN(_sha1_round_add_79_n285 ) );
NAND2_X2 _sha1_round_add_79_U29  ( .A1(_sha1_round_add_79_n358 ), .A2(_sha1_round_add_79_n357 ), .ZN(_sha1_round_add_79_n356 ) );
AND2_X4 _sha1_round_add_79_U28  ( .A1(_sha1_round_add_79_n100 ), .A2(_sha1_round_add_79_n99 ), .ZN(_sha1_round_add_79_n4 ) );
INV_X4 _sha1_round_add_79_U27  ( .A(_sha1_round_add_79_n281 ), .ZN(_sha1_round_N269 ) );
INV_X4 _sha1_round_add_79_U26  ( .A(_sha1_round_add_79_n321 ), .ZN(_sha1_round_add_79_n52 ) );
NAND2_X2 _sha1_round_add_79_U25  ( .A1(_sha1_round_add_79_n335 ), .A2(_sha1_round_add_79_n302 ), .ZN(_sha1_round_add_79_n333 ) );
NAND3_X2 _sha1_round_add_79_U24  ( .A1(_sha1_round_add_79_n225 ), .A2(_sha1_round_add_79_n229 ), .A3(_sha1_round_add_79_n224 ), .ZN(_sha1_round_add_79_n49 ) );
NAND2_X2 _sha1_round_add_79_U23  ( .A1(_sha1_round_add_79_n328 ), .A2(_sha1_round_add_79_n11 ), .ZN(_sha1_round_add_79_n325 ) );
NAND2_X2 _sha1_round_add_79_U22  ( .A1(_sha1_round_add_79_n367 ), .A2(_sha1_round_add_79_n368 ), .ZN(_sha1_round_add_79_n63 ) );
NAND2_X2 _sha1_round_add_79_U21  ( .A1(_sha1_round_add_79_n368 ), .A2(_sha1_round_add_79_n367 ), .ZN(_sha1_round_add_79_n107 ) );
NAND2_X2 _sha1_round_add_79_U20  ( .A1(_sha1_round_add_79_n359 ), .A2(_sha1_round_add_79_n340 ), .ZN(_sha1_round_add_79_n71 ) );
NOR2_X2 _sha1_round_add_79_U19  ( .A1(_sha1_round_add_79_n369 ), .A2(_sha1_round_add_79_n62 ), .ZN(_sha1_round_add_79_n368 ) );
NAND2_X2 _sha1_round_add_79_U18  ( .A1(_sha1_round_add_79_n366 ), .A2(_sha1_round_add_79_n106 ), .ZN(_sha1_round_add_79_n60 ) );
NAND2_X2 _sha1_round_add_79_U17  ( .A1(_sha1_round_add_79_n288 ), .A2(_sha1_round_add_79_n289 ), .ZN(_sha1_round_add_79_n293 ) );
NAND2_X2 _sha1_round_add_79_U16  ( .A1(_sha1_round_f [0]), .A2(_sha1_round_k_23 ), .ZN(_sha1_round_add_79_n312 ) );
NAND3_X4 _sha1_round_add_79_U15  ( .A1(_sha1_round_add_79_n274 ), .A2(_sha1_round_add_79_n275 ), .A3(_sha1_round_add_79_n276 ), .ZN(_sha1_round_add_79_n250 ) );
NOR2_X4 _sha1_round_add_79_U14  ( .A1(_sha1_round_add_79_n114 ), .A2(_sha1_round_add_79_n81 ), .ZN(_sha1_round_add_79_n112 ) );
INV_X2 _sha1_round_add_79_U13  ( .A(_sha1_round_add_79_n31 ), .ZN(_sha1_round_add_79_n319 ) );
NAND2_X4 _sha1_round_add_79_U12  ( .A1(_sha1_round_add_79_n363 ), .A2(_sha1_round_add_79_n96 ), .ZN(_sha1_round_add_79_n360 ) );
NOR3_X2 _sha1_round_add_79_U11  ( .A1(_sha1_round_add_79_n378 ), .A2(_sha1_round_add_79_n379 ), .A3(_sha1_round_add_79_n380 ), .ZN(_sha1_round_add_79_n377 ) );
NAND2_X1 _sha1_round_add_79_U10  ( .A1(_sha1_round_add_79_n8 ), .A2(_sha1_round_add_79_n63 ), .ZN(_sha1_round_add_79_n125 ) );
AND3_X4 _sha1_round_add_79_U9  ( .A1(_sha1_round_add_79_n107 ), .A2(_sha1_round_add_79_n31 ), .A3(_sha1_round_add_79_n106 ), .ZN(_sha1_round_add_79_n67 ) );
INV_X8 _sha1_round_add_79_U8  ( .A(_sha1_round_add_79_n351 ), .ZN(_sha1_round_N263 ) );
CLKBUF_X2 _sha1_round_add_79_U7  ( .A(_sha1_round_f [6]), .Z(_sha1_round_add_79_n2 ) );
NOR2_X2 _sha1_round_add_79_U6  ( .A1(_sha1_round_add_79_n17 ), .A2(_sha1_round_add_79_n132 ), .ZN(_sha1_round_add_79_n62 ) );
AND2_X2 _sha1_round_add_79_U5  ( .A1(_sha1_round_add_79_n303 ), .A2(_sha1_round_add_79_n332 ), .ZN(_sha1_round_add_79_n5 ) );
AND2_X4 _sha1_round_add_79_U4  ( .A1(_sha1_round_add_79_n205 ), .A2(_sha1_round_add_79_n193 ), .ZN(_sha1_round_add_79_n1 ) );
NOR2_X4 _sha1_round_add_79_U3  ( .A1(_sha1_round_f [2]), .A2(_sha1_round_add_79_n87 ), .ZN(_sha1_round_add_79_n132 ) );
NAND2_X2 _sha1_round_add_79_U2  ( .A1(_sha1_round_add_79_n356 ), .A2(_sha1_round_add_79_n344 ), .ZN(_sha1_round_add_79_n352 ) );
NAND2_X2 _sha1_round_add_79_2_U405  ( .A1(w[0]), .A2(rnd_q[0]), .ZN(_sha1_round_add_79_2_n223 ) );
INV_X4 _sha1_round_add_79_2_U404  ( .A(_sha1_round_add_79_2_n223 ), .ZN(_sha1_round_add_79_2_n299 ) );
NAND2_X2 _sha1_round_add_79_2_U403  ( .A1(w[9]), .A2(rnd_q[9]), .ZN(_sha1_round_add_79_2_n349 ) );
INV_X4 _sha1_round_add_79_2_U402  ( .A(_sha1_round_add_79_2_n349 ), .ZN(_sha1_round_add_79_2_n40 ) );
INV_X4 _sha1_round_add_79_2_U401  ( .A(_sha1_round_add_79_2_n83 ), .ZN(_sha1_round_add_79_2_n298 ) );
NAND2_X2 _sha1_round_add_79_2_U400  ( .A1(rnd_q[2]), .A2(w[2]), .ZN(_sha1_round_add_79_2_n374 ) );
INV_X4 _sha1_round_add_79_2_U399  ( .A(_sha1_round_add_79_2_n107 ), .ZN(_sha1_round_add_79_2_n370 ) );
NAND2_X2 _sha1_round_add_79_2_U398  ( .A1(w[3]), .A2(rnd_q[3]), .ZN(_sha1_round_add_79_2_n72 ) );
NAND2_X2 _sha1_round_add_79_2_U397  ( .A1(w[0]), .A2(rnd_q[0]), .ZN(_sha1_round_add_79_2_n372 ) );
NAND2_X2 _sha1_round_add_79_2_U396  ( .A1(w[1]), .A2(rnd_q[1]), .ZN(_sha1_round_add_79_2_n373 ) );
NAND2_X2 _sha1_round_add_79_2_U395  ( .A1(_sha1_round_add_79_2_n372 ), .A2(_sha1_round_add_79_2_n373 ), .ZN(_sha1_round_add_79_2_n369 ) );
INV_X4 _sha1_round_add_79_2_U394  ( .A(_sha1_round_add_79_2_n61 ), .ZN(_sha1_round_add_79_2_n363 ) );
INV_X4 _sha1_round_add_79_2_U393  ( .A(w[4]), .ZN(_sha1_round_add_79_2_n366 ) );
INV_X4 _sha1_round_add_79_2_U392  ( .A(rnd_q[4]), .ZN(_sha1_round_add_79_2_n367 ) );
NAND2_X2 _sha1_round_add_79_2_U391  ( .A1(_sha1_round_add_79_2_n366 ), .A2(_sha1_round_add_79_2_n367 ), .ZN(_sha1_round_add_79_2_n71 ) );
INV_X4 _sha1_round_add_79_2_U390  ( .A(_sha1_round_add_79_2_n262 ), .ZN(_sha1_round_add_79_2_n56 ) );
NAND2_X2 _sha1_round_add_79_2_U389  ( .A1(rnd_q[6]), .A2(w[6]), .ZN(_sha1_round_add_79_2_n362 ) );
INV_X4 _sha1_round_add_79_2_U388  ( .A(_sha1_round_add_79_2_n276 ), .ZN(_sha1_round_add_79_2_n358 ) );
NAND2_X2 _sha1_round_add_79_2_U387  ( .A1(w[7]), .A2(rnd_q[7]), .ZN(_sha1_round_add_79_2_n269 ) );
NAND2_X2 _sha1_round_add_79_2_U386  ( .A1(w[4]), .A2(rnd_q[4]), .ZN(_sha1_round_add_79_2_n81 ) );
NAND2_X2 _sha1_round_add_79_2_U385  ( .A1(w[5]), .A2(rnd_q[5]), .ZN(_sha1_round_add_79_2_n69 ) );
NAND2_X2 _sha1_round_add_79_2_U384  ( .A1(_sha1_round_add_79_2_n81 ), .A2(_sha1_round_add_79_2_n69 ), .ZN(_sha1_round_add_79_2_n360 ) );
INV_X4 _sha1_round_add_79_2_U383  ( .A(_sha1_round_add_79_2_n47 ), .ZN(_sha1_round_add_79_2_n321 ) );
NAND2_X2 _sha1_round_add_79_2_U382  ( .A1(w[8]), .A2(rnd_q[8]), .ZN(_sha1_round_add_79_2_n52 ) );
NAND2_X2 _sha1_round_add_79_2_U381  ( .A1(_sha1_round_add_79_2_n321 ), .A2(_sha1_round_add_79_2_n52 ), .ZN(_sha1_round_add_79_2_n357 ) );
XNOR2_X2 _sha1_round_add_79_2_U380  ( .A(_sha1_round_add_79_2_n352 ), .B(_sha1_round_add_79_2_n353 ), .ZN(_sha1_round_N294 ) );
INV_X4 _sha1_round_add_79_2_U379  ( .A(_sha1_round_add_79_2_n285 ), .ZN(_sha1_round_add_79_2_n340 ) );
XNOR2_X2 _sha1_round_add_79_2_U378  ( .A(_sha1_round_add_79_2_n344 ), .B(_sha1_round_add_79_2_n345 ), .ZN(_sha1_round_N295 ) );
INV_X4 _sha1_round_add_79_2_U377  ( .A(w[12]), .ZN(_sha1_round_add_79_2_n342 ) );
INV_X4 _sha1_round_add_79_2_U376  ( .A(rnd_q[12]), .ZN(_sha1_round_add_79_2_n343 ) );
NAND2_X2 _sha1_round_add_79_2_U375  ( .A1(_sha1_round_add_79_2_n342 ), .A2(_sha1_round_add_79_2_n343 ), .ZN(_sha1_round_add_79_2_n301 ) );
NAND2_X2 _sha1_round_add_79_2_U374  ( .A1(w[12]), .A2(rnd_q[12]), .ZN(_sha1_round_add_79_2_n292 ) );
NAND2_X2 _sha1_round_add_79_2_U373  ( .A1(_sha1_round_add_79_2_n301 ), .A2(_sha1_round_add_79_2_n292 ), .ZN(_sha1_round_add_79_2_n329 ) );
INV_X4 _sha1_round_add_79_2_U372  ( .A(_sha1_round_add_79_2_n44 ), .ZN(_sha1_round_add_79_2_n338 ) );
INV_X4 _sha1_round_add_79_2_U371  ( .A(_sha1_round_add_79_2_n264 ), .ZN(_sha1_round_add_79_2_n268 ) );
NAND2_X2 _sha1_round_add_79_2_U370  ( .A1(_sha1_round_add_79_2_n268 ), .A2(_sha1_round_add_79_2_n47 ), .ZN(_sha1_round_add_79_2_n330 ) );
INV_X4 _sha1_round_add_79_2_U369  ( .A(_sha1_round_add_79_2_n41 ), .ZN(_sha1_round_add_79_2_n336 ) );
INV_X4 _sha1_round_add_79_2_U368  ( .A(_sha1_round_add_79_2_n335 ), .ZN(_sha1_round_add_79_2_n337 ) );
NAND4_X2 _sha1_round_add_79_2_U367  ( .A1(w[8]), .A2(rnd_q[8]), .A3(_sha1_round_add_79_2_n336 ), .A4(_sha1_round_add_79_2_n337 ), .ZN(_sha1_round_add_79_2_n332 ) );
NAND2_X2 _sha1_round_add_79_2_U366  ( .A1(_sha1_round_add_79_2_n286 ), .A2(_sha1_round_add_79_2_n285 ), .ZN(_sha1_round_add_79_2_n322 ) );
INV_X4 _sha1_round_add_79_2_U365  ( .A(_sha1_round_add_79_2_n49 ), .ZN(_sha1_round_add_79_2_n273 ) );
NAND2_X2 _sha1_round_add_79_2_U364  ( .A1(_sha1_round_add_79_2_n273 ), .A2(_sha1_round_add_79_2_n268 ), .ZN(_sha1_round_add_79_2_n331 ) );
XNOR2_X2 _sha1_round_add_79_2_U363  ( .A(_sha1_round_add_79_2_n329 ), .B(_sha1_round_add_79_2_n328 ), .ZN(_sha1_round_N296 ) );
NAND2_X2 _sha1_round_add_79_2_U362  ( .A1(_sha1_round_add_79_2_n328 ), .A2(_sha1_round_add_79_2_n301 ), .ZN(_sha1_round_add_79_2_n327 ) );
NAND2_X2 _sha1_round_add_79_2_U361  ( .A1(_sha1_round_add_79_2_n327 ), .A2(_sha1_round_add_79_2_n292 ), .ZN(_sha1_round_add_79_2_n323 ) );
NAND2_X2 _sha1_round_add_79_2_U360  ( .A1(w[13]), .A2(rnd_q[13]), .ZN(_sha1_round_add_79_2_n279 ) );
INV_X4 _sha1_round_add_79_2_U359  ( .A(w[13]), .ZN(_sha1_round_add_79_2_n325 ) );
INV_X4 _sha1_round_add_79_2_U358  ( .A(rnd_q[13]), .ZN(_sha1_round_add_79_2_n326 ) );
NAND2_X2 _sha1_round_add_79_2_U357  ( .A1(_sha1_round_add_79_2_n325 ), .A2(_sha1_round_add_79_2_n326 ), .ZN(_sha1_round_add_79_2_n300 ) );
NAND2_X2 _sha1_round_add_79_2_U356  ( .A1(_sha1_round_add_79_2_n279 ), .A2(_sha1_round_add_79_2_n300 ), .ZN(_sha1_round_add_79_2_n324 ) );
XNOR2_X2 _sha1_round_add_79_2_U355  ( .A(_sha1_round_add_79_2_n323 ), .B(_sha1_round_add_79_2_n324 ), .ZN(_sha1_round_N297 ) );
INV_X4 _sha1_round_add_79_2_U354  ( .A(_sha1_round_add_79_2_n322 ), .ZN(_sha1_round_add_79_2_n319 ) );
INV_X4 _sha1_round_add_79_2_U353  ( .A(_sha1_round_add_79_2_n76 ), .ZN(_sha1_round_add_79_2_n275 ) );
NAND2_X2 _sha1_round_add_79_2_U352  ( .A1(_sha1_round_add_79_2_n317 ), .A2(_sha1_round_add_79_2_n318 ), .ZN(_sha1_round_add_79_2_n316 ) );
NAND2_X2 _sha1_round_add_79_2_U351  ( .A1(_sha1_round_add_79_2_n315 ), .A2(_sha1_round_add_79_2_n316 ), .ZN(_sha1_round_add_79_2_n314 ) );
NAND2_X2 _sha1_round_add_79_2_U350  ( .A1(_sha1_round_add_79_2_n314 ), .A2(_sha1_round_add_79_2_n301 ), .ZN(_sha1_round_add_79_2_n307 ) );
NAND2_X2 _sha1_round_add_79_2_U349  ( .A1(_sha1_round_add_79_2_n307 ), .A2(_sha1_round_add_79_2_n292 ), .ZN(_sha1_round_add_79_2_n313 ) );
NAND2_X2 _sha1_round_add_79_2_U348  ( .A1(_sha1_round_add_79_2_n313 ), .A2(_sha1_round_add_79_2_n300 ), .ZN(_sha1_round_add_79_2_n312 ) );
NAND2_X2 _sha1_round_add_79_2_U347  ( .A1(_sha1_round_add_79_2_n279 ), .A2(_sha1_round_add_79_2_n312 ), .ZN(_sha1_round_add_79_2_n308 ) );
INV_X4 _sha1_round_add_79_2_U346  ( .A(w[14]), .ZN(_sha1_round_add_79_2_n310 ) );
INV_X4 _sha1_round_add_79_2_U345  ( .A(rnd_q[14]), .ZN(_sha1_round_add_79_2_n311 ) );
NAND2_X2 _sha1_round_add_79_2_U344  ( .A1(_sha1_round_add_79_2_n310 ), .A2(_sha1_round_add_79_2_n311 ), .ZN(_sha1_round_add_79_2_n281 ) );
NAND2_X2 _sha1_round_add_79_2_U343  ( .A1(w[14]), .A2(rnd_q[14]), .ZN(_sha1_round_add_79_2_n280 ) );
NAND2_X2 _sha1_round_add_79_2_U342  ( .A1(_sha1_round_add_79_2_n281 ), .A2(_sha1_round_add_79_2_n280 ), .ZN(_sha1_round_add_79_2_n309 ) );
XNOR2_X2 _sha1_round_add_79_2_U341  ( .A(_sha1_round_add_79_2_n308 ), .B(_sha1_round_add_79_2_n309 ), .ZN(_sha1_round_N298 ) );
INV_X4 _sha1_round_add_79_2_U340  ( .A(_sha1_round_add_79_2_n280 ), .ZN(_sha1_round_add_79_2_n306 ) );
NAND2_X2 _sha1_round_add_79_2_U339  ( .A1(w[15]), .A2(rnd_q[15]), .ZN(_sha1_round_add_79_2_n284 ) );
INV_X4 _sha1_round_add_79_2_U338  ( .A(w[15]), .ZN(_sha1_round_add_79_2_n303 ) );
INV_X4 _sha1_round_add_79_2_U337  ( .A(rnd_q[15]), .ZN(_sha1_round_add_79_2_n304 ) );
NAND2_X2 _sha1_round_add_79_2_U336  ( .A1(_sha1_round_add_79_2_n303 ), .A2(_sha1_round_add_79_2_n304 ), .ZN(_sha1_round_add_79_2_n282 ) );
NAND2_X2 _sha1_round_add_79_2_U335  ( .A1(_sha1_round_add_79_2_n284 ), .A2(_sha1_round_add_79_2_n282 ), .ZN(_sha1_round_add_79_2_n302 ) );
NAND2_X2 _sha1_round_add_79_2_U334  ( .A1(w[16]), .A2(rnd_q[16]), .ZN(_sha1_round_add_79_2_n251 ) );
NAND2_X2 _sha1_round_add_79_2_U333  ( .A1(_sha1_round_add_79_2_n251 ), .A2(_sha1_round_add_79_2_n253 ), .ZN(_sha1_round_add_79_2_n254 ) );
NAND2_X2 _sha1_round_add_79_2_U332  ( .A1(_sha1_round_add_79_2_n261 ), .A2(_sha1_round_add_79_2_n268 ), .ZN(_sha1_round_add_79_2_n294 ) );
NAND2_X2 _sha1_round_add_79_2_U331  ( .A1(w[1]), .A2(rnd_q[1]), .ZN(_sha1_round_add_79_2_n108 ) );
INV_X4 _sha1_round_add_79_2_U330  ( .A(_sha1_round_add_79_2_n108 ), .ZN(_sha1_round_add_79_2_n222 ) );
NAND2_X2 _sha1_round_add_79_2_U329  ( .A1(_sha1_round_add_79_2_n296 ), .A2(_sha1_round_add_79_2_n273 ), .ZN(_sha1_round_add_79_2_n295 ) );
NAND3_X2 _sha1_round_add_79_2_U328  ( .A1(_sha1_round_add_79_2_n261 ), .A2(_sha1_round_add_79_2_n273 ), .A3(_sha1_round_add_79_2_n293 ), .ZN(_sha1_round_add_79_2_n289 ) );
INV_X4 _sha1_round_add_79_2_U327  ( .A(_sha1_round_add_79_2_n292 ), .ZN(_sha1_round_add_79_2_n291 ) );
NAND2_X2 _sha1_round_add_79_2_U326  ( .A1(_sha1_round_add_79_2_n291 ), .A2(_sha1_round_add_79_2_n261 ), .ZN(_sha1_round_add_79_2_n290 ) );
NAND2_X2 _sha1_round_add_79_2_U325  ( .A1(_sha1_round_add_79_2_n289 ), .A2(_sha1_round_add_79_2_n290 ), .ZN(_sha1_round_add_79_2_n288 ) );
NAND2_X2 _sha1_round_add_79_2_U324  ( .A1(_sha1_round_add_79_2_n279 ), .A2(_sha1_round_add_79_2_n280 ), .ZN(_sha1_round_add_79_2_n278 ) );
NAND2_X2 _sha1_round_add_79_2_U323  ( .A1(_sha1_round_add_79_2_n277 ), .A2(_sha1_round_add_79_2_n278 ), .ZN(_sha1_round_add_79_2_n270 ) );
NAND3_X2 _sha1_round_add_79_2_U322  ( .A1(_sha1_round_add_79_2_n276 ), .A2(_sha1_round_add_79_2_n261 ), .A3(_sha1_round_add_79_2_n268 ), .ZN(_sha1_round_add_79_2_n271 ) );
NAND3_X2 _sha1_round_add_79_2_U321  ( .A1(_sha1_round_add_79_2_n261 ), .A2(_sha1_round_add_79_2_n273 ), .A3(_sha1_round_add_79_2_n274 ), .ZN(_sha1_round_add_79_2_n272 ) );
NAND3_X2 _sha1_round_add_79_2_U320  ( .A1(_sha1_round_add_79_2_n270 ), .A2(_sha1_round_add_79_2_n271 ), .A3(_sha1_round_add_79_2_n272 ), .ZN(_sha1_round_add_79_2_n257 ) );
INV_X4 _sha1_round_add_79_2_U319  ( .A(_sha1_round_add_79_2_n269 ), .ZN(_sha1_round_add_79_2_n57 ) );
NAND3_X2 _sha1_round_add_79_2_U318  ( .A1(_sha1_round_add_79_2_n57 ), .A2(_sha1_round_add_79_2_n261 ), .A3(_sha1_round_add_79_2_n268 ), .ZN(_sha1_round_add_79_2_n259 ) );
NAND2_X2 _sha1_round_add_79_2_U317  ( .A1(_sha1_round_add_79_2_n81 ), .A2(_sha1_round_add_79_2_n69 ), .ZN(_sha1_round_add_79_2_n267 ) );
NAND2_X2 _sha1_round_add_79_2_U316  ( .A1(_sha1_round_add_79_2_n266 ), .A2(_sha1_round_add_79_2_n267 ), .ZN(_sha1_round_add_79_2_n265 ) );
NAND2_X2 _sha1_round_add_79_2_U315  ( .A1(_sha1_round_add_79_2_n259 ), .A2(_sha1_round_add_79_2_n260 ), .ZN(_sha1_round_add_79_2_n258 ) );
NOR2_X2 _sha1_round_add_79_2_U314  ( .A1(_sha1_round_add_79_2_n257 ), .A2(_sha1_round_add_79_2_n258 ), .ZN(_sha1_round_add_79_2_n256 ) );
XNOR2_X2 _sha1_round_add_79_2_U313  ( .A(_sha1_round_add_79_2_n254 ), .B(_sha1_round_add_79_2_n118 ), .ZN(_sha1_round_N300 ) );
INV_X4 _sha1_round_add_79_2_U312  ( .A(_sha1_round_add_79_2_n231 ), .ZN(_sha1_round_add_79_2_n253 ) );
NAND2_X2 _sha1_round_add_79_2_U311  ( .A1(_sha1_round_add_79_2_n118 ), .A2(_sha1_round_add_79_2_n253 ), .ZN(_sha1_round_add_79_2_n252 ) );
NAND2_X2 _sha1_round_add_79_2_U310  ( .A1(_sha1_round_add_79_2_n251 ), .A2(_sha1_round_add_79_2_n252 ), .ZN(_sha1_round_add_79_2_n246 ) );
INV_X4 _sha1_round_add_79_2_U309  ( .A(w[17]), .ZN(_sha1_round_add_79_2_n249 ) );
INV_X4 _sha1_round_add_79_2_U308  ( .A(rnd_q[17]), .ZN(_sha1_round_add_79_2_n250 ) );
NAND2_X2 _sha1_round_add_79_2_U307  ( .A1(_sha1_round_add_79_2_n249 ), .A2(_sha1_round_add_79_2_n250 ), .ZN(_sha1_round_add_79_2_n244 ) );
INV_X4 _sha1_round_add_79_2_U306  ( .A(_sha1_round_add_79_2_n244 ), .ZN(_sha1_round_add_79_2_n233 ) );
NAND2_X2 _sha1_round_add_79_2_U305  ( .A1(w[17]), .A2(rnd_q[17]), .ZN(_sha1_round_add_79_2_n243 ) );
INV_X4 _sha1_round_add_79_2_U304  ( .A(_sha1_round_add_79_2_n243 ), .ZN(_sha1_round_add_79_2_n248 ) );
INV_X4 _sha1_round_add_79_2_U303  ( .A(_sha1_round_add_79_2_n118 ), .ZN(_sha1_round_add_79_2_n245 ) );
NAND2_X2 _sha1_round_add_79_2_U302  ( .A1(_sha1_round_add_79_2_n242 ), .A2(_sha1_round_add_79_2_n243 ), .ZN(_sha1_round_add_79_2_n237 ) );
NAND2_X2 _sha1_round_add_79_2_U301  ( .A1(w[18]), .A2(rnd_q[18]), .ZN(_sha1_round_add_79_2_n236 ) );
INV_X4 _sha1_round_add_79_2_U300  ( .A(w[18]), .ZN(_sha1_round_add_79_2_n239 ) );
INV_X4 _sha1_round_add_79_2_U299  ( .A(rnd_q[18]), .ZN(_sha1_round_add_79_2_n240 ) );
NAND2_X2 _sha1_round_add_79_2_U298  ( .A1(_sha1_round_add_79_2_n239 ), .A2(_sha1_round_add_79_2_n240 ), .ZN(_sha1_round_add_79_2_n234 ) );
NAND2_X2 _sha1_round_add_79_2_U297  ( .A1(_sha1_round_add_79_2_n236 ), .A2(_sha1_round_add_79_2_n234 ), .ZN(_sha1_round_add_79_2_n238 ) );
NAND2_X2 _sha1_round_add_79_2_U296  ( .A1(_sha1_round_add_79_2_n237 ), .A2(_sha1_round_add_79_2_n234 ), .ZN(_sha1_round_add_79_2_n235 ) );
NAND2_X2 _sha1_round_add_79_2_U295  ( .A1(_sha1_round_add_79_2_n235 ), .A2(_sha1_round_add_79_2_n236 ), .ZN(_sha1_round_add_79_2_n185 ) );
INV_X4 _sha1_round_add_79_2_U294  ( .A(_sha1_round_add_79_2_n185 ), .ZN(_sha1_round_add_79_2_n229 ) );
INV_X4 _sha1_round_add_79_2_U293  ( .A(_sha1_round_add_79_2_n234 ), .ZN(_sha1_round_add_79_2_n232 ) );
NAND2_X2 _sha1_round_add_79_2_U292  ( .A1(_sha1_round_add_79_2_n219 ), .A2(_sha1_round_add_79_2_n118 ), .ZN(_sha1_round_add_79_2_n230 ) );
NAND2_X2 _sha1_round_add_79_2_U291  ( .A1(_sha1_round_add_79_2_n229 ), .A2(_sha1_round_add_79_2_n230 ), .ZN(_sha1_round_add_79_2_n225 ) );
INV_X4 _sha1_round_add_79_2_U290  ( .A(w[19]), .ZN(_sha1_round_add_79_2_n227 ) );
INV_X4 _sha1_round_add_79_2_U289  ( .A(rnd_q[19]), .ZN(_sha1_round_add_79_2_n228 ) );
NAND2_X2 _sha1_round_add_79_2_U288  ( .A1(_sha1_round_add_79_2_n227 ), .A2(_sha1_round_add_79_2_n228 ), .ZN(_sha1_round_add_79_2_n186 ) );
NAND2_X2 _sha1_round_add_79_2_U287  ( .A1(w[19]), .A2(rnd_q[19]), .ZN(_sha1_round_add_79_2_n220 ) );
NAND2_X2 _sha1_round_add_79_2_U286  ( .A1(_sha1_round_add_79_2_n186 ), .A2(_sha1_round_add_79_2_n220 ), .ZN(_sha1_round_add_79_2_n226 ) );
XNOR2_X2 _sha1_round_add_79_2_U285  ( .A(_sha1_round_add_79_2_n225 ), .B(_sha1_round_add_79_2_n226 ), .ZN(_sha1_round_N303 ) );
XNOR2_X2 _sha1_round_add_79_2_U284  ( .A(_sha1_round_add_79_2_n223 ), .B(_sha1_round_add_79_2_n221 ), .ZN(_sha1_round_N285 ) );
INV_X4 _sha1_round_add_79_2_U283  ( .A(_sha1_round_add_79_2_n220 ), .ZN(_sha1_round_add_79_2_n119 ) );
NAND2_X2 _sha1_round_add_79_2_U282  ( .A1(_sha1_round_add_79_2_n217 ), .A2(_sha1_round_add_79_2_n218 ), .ZN(_sha1_round_add_79_2_n205 ) );
INV_X4 _sha1_round_add_79_2_U281  ( .A(_sha1_round_add_79_2_n205 ), .ZN(_sha1_round_add_79_2_n197 ) );
XNOR2_X2 _sha1_round_add_79_2_U280  ( .A(_sha1_round_add_79_2_n197 ), .B(_sha1_round_add_79_2_n216 ), .ZN(_sha1_round_N304 ) );
NAND2_X2 _sha1_round_add_79_2_U279  ( .A1(w[21]), .A2(rnd_q[21]), .ZN(_sha1_round_add_79_2_n209 ) );
INV_X4 _sha1_round_add_79_2_U278  ( .A(_sha1_round_add_79_2_n209 ), .ZN(_sha1_round_add_79_2_n212 ) );
XNOR2_X2 _sha1_round_add_79_2_U277  ( .A(_sha1_round_add_79_2_n210 ), .B(_sha1_round_add_79_2_n211 ), .ZN(_sha1_round_N305 ) );
NAND2_X2 _sha1_round_add_79_2_U276  ( .A1(_sha1_round_add_79_2_n208 ), .A2(_sha1_round_add_79_2_n209 ), .ZN(_sha1_round_add_79_2_n195 ) );
INV_X4 _sha1_round_add_79_2_U275  ( .A(_sha1_round_add_79_2_n195 ), .ZN(_sha1_round_add_79_2_n203 ) );
NAND2_X2 _sha1_round_add_79_2_U274  ( .A1(_sha1_round_add_79_2_n198 ), .A2(_sha1_round_add_79_2_n205 ), .ZN(_sha1_round_add_79_2_n204 ) );
NAND2_X2 _sha1_round_add_79_2_U273  ( .A1(_sha1_round_add_79_2_n203 ), .A2(_sha1_round_add_79_2_n204 ), .ZN(_sha1_round_add_79_2_n199 ) );
NAND2_X2 _sha1_round_add_79_2_U272  ( .A1(w[22]), .A2(rnd_q[22]), .ZN(_sha1_round_add_79_2_n194 ) );
INV_X4 _sha1_round_add_79_2_U271  ( .A(w[22]), .ZN(_sha1_round_add_79_2_n201 ) );
INV_X4 _sha1_round_add_79_2_U270  ( .A(rnd_q[22]), .ZN(_sha1_round_add_79_2_n202 ) );
NAND2_X2 _sha1_round_add_79_2_U269  ( .A1(_sha1_round_add_79_2_n201 ), .A2(_sha1_round_add_79_2_n202 ), .ZN(_sha1_round_add_79_2_n196 ) );
NAND2_X2 _sha1_round_add_79_2_U268  ( .A1(_sha1_round_add_79_2_n194 ), .A2(_sha1_round_add_79_2_n196 ), .ZN(_sha1_round_add_79_2_n200 ) );
XNOR2_X2 _sha1_round_add_79_2_U267  ( .A(_sha1_round_add_79_2_n199 ), .B(_sha1_round_add_79_2_n200 ), .ZN(_sha1_round_N306 ) );
NAND2_X2 _sha1_round_add_79_2_U266  ( .A1(_sha1_round_add_79_2_n198 ), .A2(_sha1_round_add_79_2_n196 ), .ZN(_sha1_round_add_79_2_n188 ) );
NAND2_X2 _sha1_round_add_79_2_U265  ( .A1(_sha1_round_add_79_2_n195 ), .A2(_sha1_round_add_79_2_n196 ), .ZN(_sha1_round_add_79_2_n193 ) );
NAND2_X2 _sha1_round_add_79_2_U264  ( .A1(_sha1_round_add_79_2_n193 ), .A2(_sha1_round_add_79_2_n194 ), .ZN(_sha1_round_add_79_2_n183 ) );
INV_X4 _sha1_round_add_79_2_U263  ( .A(w[23]), .ZN(_sha1_round_add_79_2_n190 ) );
INV_X4 _sha1_round_add_79_2_U262  ( .A(rnd_q[23]), .ZN(_sha1_round_add_79_2_n191 ) );
NAND2_X2 _sha1_round_add_79_2_U261  ( .A1(_sha1_round_add_79_2_n190 ), .A2(_sha1_round_add_79_2_n191 ), .ZN(_sha1_round_add_79_2_n184 ) );
NAND2_X2 _sha1_round_add_79_2_U260  ( .A1(w[23]), .A2(rnd_q[23]), .ZN(_sha1_round_add_79_2_n129 ) );
NAND2_X2 _sha1_round_add_79_2_U259  ( .A1(_sha1_round_add_79_2_n184 ), .A2(_sha1_round_add_79_2_n129 ), .ZN(_sha1_round_add_79_2_n189 ) );
INV_X4 _sha1_round_add_79_2_U258  ( .A(_sha1_round_add_79_2_n188 ), .ZN(_sha1_round_add_79_2_n187 ) );
NAND2_X2 _sha1_round_add_79_2_U257  ( .A1(_sha1_round_add_79_2_n119 ), .A2(_sha1_round_add_79_2_n2 ), .ZN(_sha1_round_add_79_2_n170 ) );
NAND2_X2 _sha1_round_add_79_2_U256  ( .A1(_sha1_round_add_79_2_n169 ), .A2(_sha1_round_add_79_2_n170 ), .ZN(_sha1_round_add_79_2_n181 ) );
NAND2_X2 _sha1_round_add_79_2_U255  ( .A1(_sha1_round_add_79_2_n183 ), .A2(_sha1_round_add_79_2_n184 ), .ZN(_sha1_round_add_79_2_n122 ) );
NAND2_X2 _sha1_round_add_79_2_U254  ( .A1(_sha1_round_add_79_2_n122 ), .A2(_sha1_round_add_79_2_n129 ), .ZN(_sha1_round_add_79_2_n182 ) );
NOR2_X2 _sha1_round_add_79_2_U253  ( .A1(_sha1_round_add_79_2_n181 ), .A2(_sha1_round_add_79_2_n182 ), .ZN(_sha1_round_add_79_2_n180 ) );
NAND2_X2 _sha1_round_add_79_2_U252  ( .A1(w[24]), .A2(rnd_q[24]), .ZN(_sha1_round_add_79_2_n175 ) );
INV_X4 _sha1_round_add_79_2_U251  ( .A(_sha1_round_add_79_2_n175 ), .ZN(_sha1_round_add_79_2_n166 ) );
NAND2_X2 _sha1_round_add_79_2_U250  ( .A1(_sha1_round_add_79_2_n169 ), .A2(_sha1_round_add_79_2_n170 ), .ZN(_sha1_round_add_79_2_n177 ) );
NAND2_X2 _sha1_round_add_79_2_U249  ( .A1(_sha1_round_add_79_2_n122 ), .A2(_sha1_round_add_79_2_n129 ), .ZN(_sha1_round_add_79_2_n178 ) );
NOR2_X2 _sha1_round_add_79_2_U248  ( .A1(_sha1_round_add_79_2_n177 ), .A2(_sha1_round_add_79_2_n178 ), .ZN(_sha1_round_add_79_2_n176 ) );
NAND2_X2 _sha1_round_add_79_2_U247  ( .A1(_sha1_round_add_79_2_n174 ), .A2(_sha1_round_add_79_2_n175 ), .ZN(_sha1_round_add_79_2_n172 ) );
INV_X4 _sha1_round_add_79_2_U246  ( .A(_sha1_round_add_79_2_n171 ), .ZN(_sha1_round_add_79_2_n167 ) );
NAND4_X2 _sha1_round_add_79_2_U245  ( .A1(_sha1_round_add_79_2_n122 ), .A2(_sha1_round_add_79_2_n129 ), .A3(_sha1_round_add_79_2_n169 ), .A4(_sha1_round_add_79_2_n170 ), .ZN(_sha1_round_add_79_2_n168 ) );
NAND2_X2 _sha1_round_add_79_2_U244  ( .A1(w[26]), .A2(rnd_q[26]), .ZN(_sha1_round_add_79_2_n140 ) );
INV_X4 _sha1_round_add_79_2_U243  ( .A(w[26]), .ZN(_sha1_round_add_79_2_n160 ) );
INV_X4 _sha1_round_add_79_2_U242  ( .A(rnd_q[26]), .ZN(_sha1_round_add_79_2_n161 ) );
NAND2_X2 _sha1_round_add_79_2_U241  ( .A1(_sha1_round_add_79_2_n160 ), .A2(_sha1_round_add_79_2_n161 ), .ZN(_sha1_round_add_79_2_n158 ) );
NAND2_X2 _sha1_round_add_79_2_U240  ( .A1(_sha1_round_add_79_2_n140 ), .A2(_sha1_round_add_79_2_n158 ), .ZN(_sha1_round_add_79_2_n159 ) );
INV_X4 _sha1_round_add_79_2_U239  ( .A(_sha1_round_add_79_2_n140 ), .ZN(_sha1_round_add_79_2_n151 ) );
INV_X4 _sha1_round_add_79_2_U238  ( .A(_sha1_round_add_79_2_n158 ), .ZN(_sha1_round_add_79_2_n149 ) );
NAND2_X2 _sha1_round_add_79_2_U237  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(_sha1_round_add_79_2_n155 ) );
NAND2_X2 _sha1_round_add_79_2_U236  ( .A1(w[24]), .A2(rnd_q[24]), .ZN(_sha1_round_add_79_2_n156 ) );
NAND2_X2 _sha1_round_add_79_2_U235  ( .A1(_sha1_round_add_79_2_n155 ), .A2(_sha1_round_add_79_2_n156 ), .ZN(_sha1_round_add_79_2_n154 ) );
NAND2_X2 _sha1_round_add_79_2_U234  ( .A1(_sha1_round_add_79_2_n153 ), .A2(_sha1_round_add_79_2_n154 ), .ZN(_sha1_round_add_79_2_n139 ) );
INV_X4 _sha1_round_add_79_2_U233  ( .A(_sha1_round_add_79_2_n139 ), .ZN(_sha1_round_add_79_2_n152 ) );
NAND2_X2 _sha1_round_add_79_2_U232  ( .A1(_sha1_round_add_79_2_n141 ), .A2(_sha1_round_add_79_2_n131 ), .ZN(_sha1_round_add_79_2_n147 ) );
NAND2_X2 _sha1_round_add_79_2_U231  ( .A1(_sha1_round_add_79_2_n146 ), .A2(_sha1_round_add_79_2_n147 ), .ZN(_sha1_round_add_79_2_n142 ) );
INV_X4 _sha1_round_add_79_2_U230  ( .A(w[27]), .ZN(_sha1_round_add_79_2_n144 ) );
INV_X4 _sha1_round_add_79_2_U229  ( .A(rnd_q[27]), .ZN(_sha1_round_add_79_2_n145 ) );
NAND2_X2 _sha1_round_add_79_2_U228  ( .A1(_sha1_round_add_79_2_n144 ), .A2(_sha1_round_add_79_2_n145 ), .ZN(_sha1_round_add_79_2_n130 ) );
NAND2_X2 _sha1_round_add_79_2_U227  ( .A1(w[27]), .A2(rnd_q[27]), .ZN(_sha1_round_add_79_2_n137 ) );
NAND2_X2 _sha1_round_add_79_2_U226  ( .A1(_sha1_round_add_79_2_n130 ), .A2(_sha1_round_add_79_2_n137 ), .ZN(_sha1_round_add_79_2_n143 ) );
XNOR2_X2 _sha1_round_add_79_2_U225  ( .A(_sha1_round_add_79_2_n142 ), .B(_sha1_round_add_79_2_n143 ), .ZN(_sha1_round_N311 ) );
NAND2_X2 _sha1_round_add_79_2_U224  ( .A1(_sha1_round_add_79_2_n139 ), .A2(_sha1_round_add_79_2_n140 ), .ZN(_sha1_round_add_79_2_n138 ) );
NAND2_X2 _sha1_round_add_79_2_U223  ( .A1(_sha1_round_add_79_2_n138 ), .A2(_sha1_round_add_79_2_n130 ), .ZN(_sha1_round_add_79_2_n136 ) );
NAND2_X2 _sha1_round_add_79_2_U222  ( .A1(_sha1_round_add_79_2_n136 ), .A2(_sha1_round_add_79_2_n137 ), .ZN(_sha1_round_add_79_2_n125 ) );
INV_X4 _sha1_round_add_79_2_U221  ( .A(w[28]), .ZN(_sha1_round_add_79_2_n134 ) );
INV_X4 _sha1_round_add_79_2_U220  ( .A(rnd_q[28]), .ZN(_sha1_round_add_79_2_n135 ) );
NAND2_X2 _sha1_round_add_79_2_U219  ( .A1(_sha1_round_add_79_2_n134 ), .A2(_sha1_round_add_79_2_n135 ), .ZN(_sha1_round_add_79_2_n126 ) );
NAND2_X2 _sha1_round_add_79_2_U218  ( .A1(w[28]), .A2(rnd_q[28]), .ZN(_sha1_round_add_79_2_n132 ) );
NAND2_X2 _sha1_round_add_79_2_U217  ( .A1(_sha1_round_add_79_2_n126 ), .A2(_sha1_round_add_79_2_n132 ), .ZN(_sha1_round_add_79_2_n133 ) );
INV_X4 _sha1_round_add_79_2_U216  ( .A(_sha1_round_add_79_2_n132 ), .ZN(_sha1_round_add_79_2_n127 ) );
NAND2_X2 _sha1_round_add_79_2_U215  ( .A1(_sha1_round_add_79_2_n125 ), .A2(_sha1_round_add_79_2_n126 ), .ZN(_sha1_round_add_79_2_n124 ) );
NAND2_X2 _sha1_round_add_79_2_U214  ( .A1(_sha1_round_add_79_2_n123 ), .A2(_sha1_round_add_79_2_n124 ), .ZN(_sha1_round_add_79_2_n97 ) );
INV_X4 _sha1_round_add_79_2_U213  ( .A(_sha1_round_add_79_2_n122 ), .ZN(_sha1_round_add_79_2_n120 ) );
INV_X4 _sha1_round_add_79_2_U212  ( .A(_sha1_round_add_79_2_n121 ), .ZN(_sha1_round_add_79_2_n115 ) );
NAND2_X2 _sha1_round_add_79_2_U211  ( .A1(_sha1_round_add_79_2_n116 ), .A2(_sha1_round_add_79_2_n117 ), .ZN(_sha1_round_add_79_2_n94 ) );
NAND2_X2 _sha1_round_add_79_2_U210  ( .A1(_sha1_round_add_79_2_n94 ), .A2(_sha1_round_add_79_2_n3 ), .ZN(_sha1_round_add_79_2_n114 ) );
NAND2_X2 _sha1_round_add_79_2_U209  ( .A1(_sha1_round_add_79_2_n113 ), .A2(_sha1_round_add_79_2_n114 ), .ZN(_sha1_round_add_79_2_n109 ) );
NAND2_X2 _sha1_round_add_79_2_U208  ( .A1(w[29]), .A2(rnd_q[29]), .ZN(_sha1_round_add_79_2_n96 ) );
INV_X4 _sha1_round_add_79_2_U207  ( .A(w[29]), .ZN(_sha1_round_add_79_2_n111 ) );
INV_X4 _sha1_round_add_79_2_U206  ( .A(rnd_q[29]), .ZN(_sha1_round_add_79_2_n112 ) );
NAND2_X2 _sha1_round_add_79_2_U205  ( .A1(_sha1_round_add_79_2_n111 ), .A2(_sha1_round_add_79_2_n112 ), .ZN(_sha1_round_add_79_2_n99 ) );
NAND2_X2 _sha1_round_add_79_2_U204  ( .A1(_sha1_round_add_79_2_n96 ), .A2(_sha1_round_add_79_2_n99 ), .ZN(_sha1_round_add_79_2_n110 ) );
XNOR2_X2 _sha1_round_add_79_2_U203  ( .A(_sha1_round_add_79_2_n109 ), .B(_sha1_round_add_79_2_n110 ), .ZN(_sha1_round_N313 ) );
XNOR2_X2 _sha1_round_add_79_2_U202  ( .A(_sha1_round_add_79_2_n86 ), .B(_sha1_round_add_79_2_n106 ), .ZN(_sha1_round_N286 ) );
NAND2_X2 _sha1_round_add_79_2_U201  ( .A1(_sha1_round_add_79_2_n97 ), .A2(_sha1_round_add_79_2_n99 ), .ZN(_sha1_round_add_79_2_n103 ) );
NAND2_X2 _sha1_round_add_79_2_U200  ( .A1(_sha1_round_add_79_2_n1 ), .A2(_sha1_round_add_79_2_n99 ), .ZN(_sha1_round_add_79_2_n104 ) );
NAND4_X2 _sha1_round_add_79_2_U199  ( .A1(_sha1_round_add_79_2_n103 ), .A2(_sha1_round_add_79_2_n96 ), .A3(_sha1_round_add_79_2_n104 ), .A4(_sha1_round_add_79_2_n105 ), .ZN(_sha1_round_add_79_2_n100 ) );
INV_X4 _sha1_round_add_79_2_U198  ( .A(w[30]), .ZN(_sha1_round_add_79_2_n101 ) );
INV_X4 _sha1_round_add_79_2_U197  ( .A(rnd_q[30]), .ZN(_sha1_round_add_79_2_n102 ) );
INV_X4 _sha1_round_add_79_2_U196  ( .A(_sha1_round_add_79_2_n99 ), .ZN(_sha1_round_add_79_2_n98 ) );
NAND2_X2 _sha1_round_add_79_2_U195  ( .A1(_sha1_round_add_79_2_n93 ), .A2(_sha1_round_add_79_2_n97 ), .ZN(_sha1_round_add_79_2_n89 ) );
NAND2_X2 _sha1_round_add_79_2_U194  ( .A1(_sha1_round_add_79_2_n93 ), .A2(_sha1_round_add_79_2_n1 ), .ZN(_sha1_round_add_79_2_n91 ) );
NAND4_X2 _sha1_round_add_79_2_U193  ( .A1(_sha1_round_add_79_2_n89 ), .A2(_sha1_round_add_79_2_n90 ), .A3(_sha1_round_add_79_2_n91 ), .A4(_sha1_round_add_79_2_n92 ), .ZN(_sha1_round_add_79_2_n87 ) );
XNOR2_X2 _sha1_round_add_79_2_U192  ( .A(w[31]), .B(rnd_q[31]), .ZN(_sha1_round_add_79_2_n88 ) );
XNOR2_X2 _sha1_round_add_79_2_U191  ( .A(_sha1_round_add_79_2_n87 ), .B(_sha1_round_add_79_2_n88 ), .ZN(_sha1_round_N315 ) );
NAND2_X2 _sha1_round_add_79_2_U190  ( .A1(_sha1_round_add_79_2_n72 ), .A2(_sha1_round_add_79_2_n83 ), .ZN(_sha1_round_add_79_2_n82 ) );
INV_X4 _sha1_round_add_79_2_U189  ( .A(_sha1_round_add_79_2_n71 ), .ZN(_sha1_round_add_79_2_n64 ) );
INV_X4 _sha1_round_add_79_2_U188  ( .A(_sha1_round_add_79_2_n81 ), .ZN(_sha1_round_add_79_2_n75 ) );
XNOR2_X2 _sha1_round_add_79_2_U187  ( .A(_sha1_round_add_79_2_n48 ), .B(_sha1_round_add_79_2_n80 ), .ZN(_sha1_round_N288 ) );
INV_X4 _sha1_round_add_79_2_U186  ( .A(_sha1_round_add_79_2_n69 ), .ZN(_sha1_round_add_79_2_n62 ) );
XNOR2_X2 _sha1_round_add_79_2_U185  ( .A(_sha1_round_add_79_2_n77 ), .B(_sha1_round_add_79_2_n78 ), .ZN(_sha1_round_N289 ) );
INV_X4 _sha1_round_add_79_2_U184  ( .A(_sha1_round_add_79_2_n60 ), .ZN(_sha1_round_add_79_2_n70 ) );
NAND2_X2 _sha1_round_add_79_2_U183  ( .A1(_sha1_round_add_79_2_n68 ), .A2(_sha1_round_add_79_2_n69 ), .ZN(_sha1_round_add_79_2_n67 ) );
INV_X4 _sha1_round_add_79_2_U182  ( .A(_sha1_round_add_79_2_n66 ), .ZN(_sha1_round_add_79_2_n65 ) );
XNOR2_X2 _sha1_round_add_79_2_U181  ( .A(_sha1_round_add_79_2_n54 ), .B(_sha1_round_add_79_2_n55 ), .ZN(_sha1_round_N291 ) );
INV_X4 _sha1_round_add_79_2_U180  ( .A(_sha1_round_add_79_2_n52 ), .ZN(_sha1_round_add_79_2_n43 ) );
XNOR2_X2 _sha1_round_add_79_2_U179  ( .A(_sha1_round_add_79_2_n50 ), .B(_sha1_round_add_79_2_n51 ), .ZN(_sha1_round_N292 ) );
XNOR2_X2 _sha1_round_add_79_2_U178  ( .A(_sha1_round_add_79_2_n38 ), .B(_sha1_round_add_79_2_n39 ), .ZN(_sha1_round_N293 ) );
NAND2_X2 _sha1_round_add_79_2_U177  ( .A1(_sha1_round_add_79_2_n72 ), .A2(_sha1_round_add_79_2_n73 ), .ZN(_sha1_round_add_79_2_n368 ) );
AND2_X2 _sha1_round_add_79_2_U176  ( .A1(w[11]), .A2(rnd_q[11]), .ZN(_sha1_round_add_79_2_n37 ) );
AND2_X2 _sha1_round_add_79_2_U175  ( .A1(w[2]), .A2(rnd_q[2]), .ZN(_sha1_round_add_79_2_n36 ) );
AND2_X2 _sha1_round_add_79_2_U174  ( .A1(w[6]), .A2(rnd_q[6]), .ZN(_sha1_round_add_79_2_n35 ) );
NOR2_X2 _sha1_round_add_79_2_U173  ( .A1(rnd_q[20]), .A2(w[20]), .ZN(_sha1_round_add_79_2_n207 ) );
NOR2_X2 _sha1_round_add_79_2_U172  ( .A1(rnd_q[21]), .A2(w[21]), .ZN(_sha1_round_add_79_2_n206 ) );
NOR2_X2 _sha1_round_add_79_2_U171  ( .A1(_sha1_round_add_79_2_n206 ), .A2(_sha1_round_add_79_2_n207 ), .ZN(_sha1_round_add_79_2_n198 ) );
NOR2_X2 _sha1_round_add_79_2_U170  ( .A1(rnd_q[10]), .A2(w[10]), .ZN(_sha1_round_add_79_2_n341 ) );
AND2_X2 _sha1_round_add_79_2_U169  ( .A1(w[10]), .A2(rnd_q[10]), .ZN(_sha1_round_add_79_2_n34 ) );
OR2_X2 _sha1_round_add_79_2_U168  ( .A1(w[3]), .A2(rnd_q[3]), .ZN(_sha1_round_add_79_2_n83 ) );
NOR2_X2 _sha1_round_add_79_2_U167  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(_sha1_round_add_79_2_n157 ) );
NOR2_X2 _sha1_round_add_79_2_U166  ( .A1(_sha1_round_add_79_2_n149 ), .A2(_sha1_round_add_79_2_n157 ), .ZN(_sha1_round_add_79_2_n153 ) );
NAND3_X2 _sha1_round_add_79_2_U165  ( .A1(rnd_q[20]), .A2(_sha1_round_add_79_2_n11 ), .A3(w[20]), .ZN(_sha1_round_add_79_2_n208 ) );
NAND3_X2 _sha1_round_add_79_2_U164  ( .A1(rnd_q[16]), .A2(w[16]), .A3(_sha1_round_add_79_2_n244 ), .ZN(_sha1_round_add_79_2_n242 ) );
NOR2_X2 _sha1_round_add_79_2_U163  ( .A1(rnd_q[20]), .A2(w[20]), .ZN(_sha1_round_add_79_2_n215 ) );
NOR2_X2 _sha1_round_add_79_2_U162  ( .A1(rnd_q[5]), .A2(w[5]), .ZN(_sha1_round_add_79_2_n365 ) );
NOR2_X2 _sha1_round_add_79_2_U161  ( .A1(_sha1_round_add_79_2_n56 ), .A2(_sha1_round_add_79_2_n365 ), .ZN(_sha1_round_add_79_2_n364 ) );
NOR2_X2 _sha1_round_add_79_2_U160  ( .A1(_sha1_round_add_79_2_n9 ), .A2(_sha1_round_add_79_2_n95 ), .ZN(_sha1_round_add_79_2_n90 ) );
NOR2_X2 _sha1_round_add_79_2_U159  ( .A1(_sha1_round_add_79_2_n298 ), .A2(_sha1_round_add_79_2_n374 ), .ZN(_sha1_round_add_79_2_n76 ) );
NOR2_X2 _sha1_round_add_79_2_U158  ( .A1(rnd_q[0]), .A2(w[0]), .ZN(_sha1_round_add_79_2_n224 ) );
NOR2_X2 _sha1_round_add_79_2_U157  ( .A1(_sha1_round_add_79_2_n299 ), .A2(_sha1_round_add_79_2_n224 ), .ZN(_sha1_round_N284 ) );
NOR2_X2 _sha1_round_add_79_2_U156  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(_sha1_round_add_79_2_n164 ) );
NAND3_X2 _sha1_round_add_79_2_U155  ( .A1(rnd_q[9]), .A2(w[9]), .A3(_sha1_round_add_79_2_n337 ), .ZN(_sha1_round_add_79_2_n333 ) );
NOR2_X2 _sha1_round_add_79_2_U154  ( .A1(_sha1_round_add_79_2_n34 ), .A2(_sha1_round_add_79_2_n37 ), .ZN(_sha1_round_add_79_2_n334 ) );
NAND3_X2 _sha1_round_add_79_2_U153  ( .A1(_sha1_round_add_79_2_n332 ), .A2(_sha1_round_add_79_2_n333 ), .A3(_sha1_round_add_79_2_n334 ), .ZN(_sha1_round_add_79_2_n286 ) );
NOR2_X2 _sha1_round_add_79_2_U152  ( .A1(rnd_q[10]), .A2(w[10]), .ZN(_sha1_round_add_79_2_n335 ) );
NOR2_X2 _sha1_round_add_79_2_U151  ( .A1(rnd_q[21]), .A2(w[21]), .ZN(_sha1_round_add_79_2_n213 ) );
NOR2_X2 _sha1_round_add_79_2_U150  ( .A1(_sha1_round_add_79_2_n214 ), .A2(_sha1_round_add_79_2_n7 ), .ZN(_sha1_round_add_79_2_n210 ) );
NOR2_X2 _sha1_round_add_79_2_U149  ( .A1(_sha1_round_add_79_2_n212 ), .A2(_sha1_round_add_79_2_n213 ), .ZN(_sha1_round_add_79_2_n211 ) );
NOR2_X2 _sha1_round_add_79_2_U148  ( .A1(rnd_q[9]), .A2(w[9]), .ZN(_sha1_round_add_79_2_n41 ) );
NOR2_X2 _sha1_round_add_79_2_U147  ( .A1(rnd_q[8]), .A2(w[8]), .ZN(_sha1_round_add_79_2_n44 ) );
NOR2_X2 _sha1_round_add_79_2_U146  ( .A1(rnd_q[16]), .A2(w[16]), .ZN(_sha1_round_add_79_2_n231 ) );
OR2_X2 _sha1_round_add_79_2_U145  ( .A1(w[11]), .A2(rnd_q[11]), .ZN(_sha1_round_add_79_2_n285 ) );
NOR2_X2 _sha1_round_add_79_2_U144  ( .A1(rnd_q[24]), .A2(w[24]), .ZN(_sha1_round_add_79_2_n148 ) );
NOR2_X2 _sha1_round_add_79_2_U143  ( .A1(rnd_q[1]), .A2(w[1]), .ZN(_sha1_round_add_79_2_n107 ) );
NOR2_X2 _sha1_round_add_79_2_U142  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(_sha1_round_add_79_2_n150 ) );
NOR3_X2 _sha1_round_add_79_2_U141  ( .A1(_sha1_round_add_79_2_n148 ), .A2(_sha1_round_add_79_2_n149 ), .A3(_sha1_round_add_79_2_n150 ), .ZN(_sha1_round_add_79_2_n131 ) );
NOR2_X2 _sha1_round_add_79_2_U140  ( .A1(rnd_q[2]), .A2(w[2]), .ZN(_sha1_round_add_79_2_n85 ) );
NOR2_X2 _sha1_round_add_79_2_U139  ( .A1(rnd_q[6]), .A2(w[6]), .ZN(_sha1_round_add_79_2_n61 ) );
NOR2_X2 _sha1_round_add_79_2_U138  ( .A1(rnd_q[5]), .A2(w[5]), .ZN(_sha1_round_add_79_2_n60 ) );
OR2_X2 _sha1_round_add_79_2_U137  ( .A1(w[7]), .A2(rnd_q[7]), .ZN(_sha1_round_add_79_2_n262 ) );
NOR2_X2 _sha1_round_add_79_2_U136  ( .A1(_sha1_round_add_79_2_n4 ), .A2(_sha1_round_add_79_2_n96 ), .ZN(_sha1_round_add_79_2_n95 ) );
NOR2_X2 _sha1_round_add_79_2_U135  ( .A1(_sha1_round_add_79_2_n4 ), .A2(_sha1_round_add_79_2_n98 ), .ZN(_sha1_round_add_79_2_n93 ) );
OR2_X2 _sha1_round_add_79_2_U134  ( .A1(_sha1_round_add_79_2_n60 ), .A2(_sha1_round_add_79_2_n61 ), .ZN(_sha1_round_add_79_2_n33 ) );
AND3_X2 _sha1_round_add_79_2_U133  ( .A1(_sha1_round_add_79_2_n131 ), .A2(_sha1_round_add_79_2_n130 ), .A3(_sha1_round_add_79_2_n141 ), .ZN(_sha1_round_add_79_2_n32 ) );
OR2_X2 _sha1_round_add_79_2_U132  ( .A1(_sha1_round_add_79_2_n44 ), .A2(_sha1_round_add_79_2_n41 ), .ZN(_sha1_round_add_79_2_n31 ) );
AND2_X2 _sha1_round_add_79_2_U131  ( .A1(_sha1_round_add_79_2_n282 ), .A2(_sha1_round_add_79_2_n281 ), .ZN(_sha1_round_add_79_2_n277 ) );
NOR2_X2 _sha1_round_add_79_2_U130  ( .A1(_sha1_round_add_79_2_n340 ), .A2(_sha1_round_add_79_2_n341 ), .ZN(_sha1_round_add_79_2_n339 ) );
NAND3_X2 _sha1_round_add_79_2_U129  ( .A1(_sha1_round_add_79_2_n336 ), .A2(_sha1_round_add_79_2_n338 ), .A3(_sha1_round_add_79_2_n339 ), .ZN(_sha1_round_add_79_2_n264 ) );
NAND3_X2 _sha1_round_add_79_2_U128  ( .A1(_sha1_round_add_79_2_n70 ), .A2(_sha1_round_add_79_2_n71 ), .A3(_sha1_round_add_79_2_n66 ), .ZN(_sha1_round_add_79_2_n68 ) );
NAND3_X2 _sha1_round_add_79_2_U127  ( .A1(_sha1_round_add_79_2_n3 ), .A2(_sha1_round_add_79_2_n99 ), .A3(_sha1_round_add_79_2_n94 ), .ZN(_sha1_round_add_79_2_n105 ) );
NOR2_X2 _sha1_round_add_79_2_U126  ( .A1(_sha1_round_add_79_2_n222 ), .A2(_sha1_round_add_79_2_n107 ), .ZN(_sha1_round_add_79_2_n221 ) );
NOR2_X2 _sha1_round_add_79_2_U125  ( .A1(_sha1_round_add_79_2_n61 ), .A2(_sha1_round_add_79_2_n60 ), .ZN(_sha1_round_add_79_2_n266 ) );
NOR2_X2 _sha1_round_add_79_2_U124  ( .A1(_sha1_round_add_79_2_n48 ), .A2(_sha1_round_add_79_2_n49 ), .ZN(_sha1_round_add_79_2_n356 ) );
NOR2_X2 _sha1_round_add_79_2_U123  ( .A1(_sha1_round_add_79_2_n356 ), .A2(_sha1_round_add_79_2_n357 ), .ZN(_sha1_round_add_79_2_n355 ) );
NOR2_X2 _sha1_round_add_79_2_U122  ( .A1(_sha1_round_add_79_2_n48 ), .A2(_sha1_round_add_79_2_n49 ), .ZN(_sha1_round_add_79_2_n350 ) );
NAND3_X2 _sha1_round_add_79_2_U121  ( .A1(_sha1_round_add_79_2_n52 ), .A2(_sha1_round_add_79_2_n349 ), .A3(_sha1_round_add_79_2_n321 ), .ZN(_sha1_round_add_79_2_n351 ) );
NOR2_X2 _sha1_round_add_79_2_U120  ( .A1(_sha1_round_add_79_2_n350 ), .A2(_sha1_round_add_79_2_n351 ), .ZN(_sha1_round_add_79_2_n347 ) );
NOR2_X2 _sha1_round_add_79_2_U119  ( .A1(_sha1_round_add_79_2_n48 ), .A2(_sha1_round_add_79_2_n49 ), .ZN(_sha1_round_add_79_2_n46 ) );
NOR2_X2 _sha1_round_add_79_2_U118  ( .A1(_sha1_round_add_79_2_n46 ), .A2(_sha1_round_add_79_2_n47 ), .ZN(_sha1_round_add_79_2_n45 ) );
NAND3_X2 _sha1_round_add_79_2_U117  ( .A1(_sha1_round_add_79_2_n73 ), .A2(_sha1_round_add_79_2_n72 ), .A3(_sha1_round_add_79_2_n275 ), .ZN(_sha1_round_add_79_2_n318 ) );
NOR4_X2 _sha1_round_add_79_2_U116  ( .A1(_sha1_round_add_79_2_n297 ), .A2(_sha1_round_add_79_2_n298 ), .A3(_sha1_round_add_79_2_n85 ), .A4(_sha1_round_add_79_2_n107 ), .ZN(_sha1_round_add_79_2_n296 ) );
NOR2_X2 _sha1_round_add_79_2_U115  ( .A1(_sha1_round_add_79_2_n294 ), .A2(_sha1_round_add_79_2_n295 ), .ZN(_sha1_round_add_79_2_n287 ) );
NOR2_X2 _sha1_round_add_79_2_U114  ( .A1(_sha1_round_add_79_2_n121 ), .A2(_sha1_round_add_79_2_n129 ), .ZN(_sha1_round_add_79_2_n128 ) );
NOR2_X2 _sha1_round_add_79_2_U113  ( .A1(_sha1_round_add_79_2_n151 ), .A2(_sha1_round_add_79_2_n152 ), .ZN(_sha1_round_add_79_2_n146 ) );
NOR2_X2 _sha1_round_add_79_2_U112  ( .A1(_sha1_round_add_79_2_n166 ), .A2(_sha1_round_add_79_2_n6 ), .ZN(_sha1_round_add_79_2_n165 ) );
NOR2_X2 _sha1_round_add_79_2_U111  ( .A1(_sha1_round_add_79_2_n164 ), .A2(_sha1_round_add_79_2_n165 ), .ZN(_sha1_round_add_79_2_n163 ) );
NOR2_X2 _sha1_round_add_79_2_U110  ( .A1(_sha1_round_add_79_2_n85 ), .A2(_sha1_round_add_79_2_n86 ), .ZN(_sha1_round_add_79_2_n84 ) );
NAND3_X2 _sha1_round_add_79_2_U109  ( .A1(_sha1_round_add_79_2_n185 ), .A2(_sha1_round_add_79_2_n186 ), .A3(_sha1_round_add_79_2_n2 ), .ZN(_sha1_round_add_79_2_n169 ) );
NOR2_X2 _sha1_round_add_79_2_U108  ( .A1(_sha1_round_add_79_2_n75 ), .A2(_sha1_round_add_79_2_n76 ), .ZN(_sha1_round_add_79_2_n74 ) );
NAND3_X2 _sha1_round_add_79_2_U107  ( .A1(_sha1_round_add_79_2_n73 ), .A2(_sha1_round_add_79_2_n74 ), .A3(_sha1_round_add_79_2_n72 ), .ZN(_sha1_round_add_79_2_n66 ) );
NOR2_X2 _sha1_round_add_79_2_U106  ( .A1(_sha1_round_add_79_2_n298 ), .A2(_sha1_round_add_79_2_n85 ), .ZN(_sha1_round_add_79_2_n371 ) );
NAND3_X2 _sha1_round_add_79_2_U105  ( .A1(_sha1_round_add_79_2_n369 ), .A2(_sha1_round_add_79_2_n370 ), .A3(_sha1_round_add_79_2_n371 ), .ZN(_sha1_round_add_79_2_n73 ) );
NAND3_X2 _sha1_round_add_79_2_U104  ( .A1(_sha1_round_add_79_2_n358 ), .A2(_sha1_round_add_79_2_n269 ), .A3(_sha1_round_add_79_2_n359 ), .ZN(_sha1_round_add_79_2_n47 ) );
AND2_X4 _sha1_round_add_79_2_U103  ( .A1(_sha1_round_add_79_2_n31 ), .A2(_sha1_round_add_79_2_n349 ), .ZN(_sha1_round_add_79_2_n29 ) );
OR2_X2 _sha1_round_add_79_2_U102  ( .A1(_sha1_round_add_79_2_n29 ), .A2(_sha1_round_add_79_2_n335 ), .ZN(_sha1_round_add_79_2_n348 ) );
NAND3_X2 _sha1_round_add_79_2_U101  ( .A1(_sha1_round_add_79_2_n130 ), .A2(_sha1_round_add_79_2_n126 ), .A3(_sha1_round_add_79_2_n131 ), .ZN(_sha1_round_add_79_2_n121 ) );
NOR3_X2 _sha1_round_add_79_2_U100  ( .A1(_sha1_round_add_79_2_n245 ), .A2(_sha1_round_add_79_2_n233 ), .A3(_sha1_round_add_79_2_n231 ), .ZN(_sha1_round_add_79_2_n241 ) );
NOR2_X2 _sha1_round_add_79_2_U99  ( .A1(_sha1_round_add_79_2_n60 ), .A2(_sha1_round_add_79_2_n61 ), .ZN(_sha1_round_add_79_2_n361 ) );
OR2_X4 _sha1_round_add_79_2_U98  ( .A1(_sha1_round_add_79_2_n107 ), .A2(_sha1_round_add_79_2_n223 ), .ZN(_sha1_round_add_79_2_n28 ) );
AND2_X2 _sha1_round_add_79_2_U97  ( .A1(_sha1_round_add_79_2_n108 ), .A2(_sha1_round_add_79_2_n28 ), .ZN(_sha1_round_add_79_2_n86 ) );
NOR3_X2 _sha1_round_add_79_2_U96  ( .A1(_sha1_round_add_79_2_n231 ), .A2(_sha1_round_add_79_2_n232 ), .A3(_sha1_round_add_79_2_n233 ), .ZN(_sha1_round_add_79_2_n219 ) );
OR2_X4 _sha1_round_add_79_2_U95  ( .A1(_sha1_round_add_79_2_n4 ), .A2(_sha1_round_add_79_2_n9 ), .ZN(_sha1_round_add_79_2_n27 ) );
XNOR2_X2 _sha1_round_add_79_2_U94  ( .A(_sha1_round_add_79_2_n100 ), .B(_sha1_round_add_79_2_n27 ), .ZN(_sha1_round_N314 ) );
NOR2_X2 _sha1_round_add_79_2_U93  ( .A1(_sha1_round_add_79_2_n319 ), .A2(_sha1_round_add_79_2_n320 ), .ZN(_sha1_round_add_79_2_n315 ) );
NOR2_X2 _sha1_round_add_79_2_U92  ( .A1(_sha1_round_add_79_2_n127 ), .A2(_sha1_round_add_79_2_n128 ), .ZN(_sha1_round_add_79_2_n123 ) );
NOR2_X2 _sha1_round_add_79_2_U91  ( .A1(_sha1_round_add_79_2_n164 ), .A2(_sha1_round_add_79_2_n6 ), .ZN(_sha1_round_add_79_2_n173 ) );
XOR2_X2 _sha1_round_add_79_2_U90  ( .A(_sha1_round_add_79_2_n172 ), .B(_sha1_round_add_79_2_n173 ), .Z(_sha1_round_N309 ) );
NOR2_X2 _sha1_round_add_79_2_U89  ( .A1(_sha1_round_add_79_2_n355 ), .A2(_sha1_round_add_79_2_n31 ), .ZN(_sha1_round_add_79_2_n354 ) );
NOR2_X2 _sha1_round_add_79_2_U88  ( .A1(_sha1_round_add_79_2_n40 ), .A2(_sha1_round_add_79_2_n354 ), .ZN(_sha1_round_add_79_2_n352 ) );
NOR2_X2 _sha1_round_add_79_2_U87  ( .A1(_sha1_round_add_79_2_n34 ), .A2(_sha1_round_add_79_2_n335 ), .ZN(_sha1_round_add_79_2_n353 ) );
NOR2_X2 _sha1_round_add_79_2_U86  ( .A1(_sha1_round_add_79_2_n97 ), .A2(_sha1_round_add_79_2_n1 ), .ZN(_sha1_round_add_79_2_n113 ) );
NOR2_X2 _sha1_round_add_79_2_U85  ( .A1(_sha1_round_add_79_2_n233 ), .A2(_sha1_round_add_79_2_n248 ), .ZN(_sha1_round_add_79_2_n247 ) );
XOR2_X2 _sha1_round_add_79_2_U84  ( .A(_sha1_round_add_79_2_n246 ), .B(_sha1_round_add_79_2_n247 ), .Z(_sha1_round_N301 ) );
OR2_X4 _sha1_round_add_79_2_U83  ( .A1(_sha1_round_add_79_2_n32 ), .A2(_sha1_round_add_79_2_n125 ), .ZN(_sha1_round_add_79_2_n25 ) );
XNOR2_X2 _sha1_round_add_79_2_U82  ( .A(_sha1_round_add_79_2_n25 ), .B(_sha1_round_add_79_2_n133 ), .ZN(_sha1_round_N312 ) );
NOR2_X2 _sha1_round_add_79_2_U81  ( .A1(_sha1_round_add_79_2_n148 ), .A2(_sha1_round_add_79_2_n166 ), .ZN(_sha1_round_add_79_2_n179 ) );
XOR2_X2 _sha1_round_add_79_2_U80  ( .A(_sha1_round_add_79_2_n141 ), .B(_sha1_round_add_79_2_n179 ), .Z(_sha1_round_N308 ) );
NOR2_X2 _sha1_round_add_79_2_U79  ( .A1(_sha1_round_add_79_2_n48 ), .A2(_sha1_round_add_79_2_n49 ), .ZN(_sha1_round_add_79_2_n53 ) );
NOR2_X2 _sha1_round_add_79_2_U78  ( .A1(_sha1_round_add_79_2_n53 ), .A2(_sha1_round_add_79_2_n47 ), .ZN(_sha1_round_add_79_2_n50 ) );
NOR2_X2 _sha1_round_add_79_2_U77  ( .A1(_sha1_round_add_79_2_n44 ), .A2(_sha1_round_add_79_2_n43 ), .ZN(_sha1_round_add_79_2_n51 ) );
NOR2_X2 _sha1_round_add_79_2_U76  ( .A1(_sha1_round_add_79_2_n44 ), .A2(_sha1_round_add_79_2_n45 ), .ZN(_sha1_round_add_79_2_n42 ) );
NOR2_X2 _sha1_round_add_79_2_U75  ( .A1(_sha1_round_add_79_2_n42 ), .A2(_sha1_round_add_79_2_n43 ), .ZN(_sha1_round_add_79_2_n38 ) );
NOR2_X2 _sha1_round_add_79_2_U74  ( .A1(_sha1_round_add_79_2_n40 ), .A2(_sha1_round_add_79_2_n41 ), .ZN(_sha1_round_add_79_2_n39 ) );
NOR2_X2 _sha1_round_add_79_2_U73  ( .A1(_sha1_round_add_79_2_n347 ), .A2(_sha1_round_add_79_2_n348 ), .ZN(_sha1_round_add_79_2_n346 ) );
NOR2_X2 _sha1_round_add_79_2_U72  ( .A1(_sha1_round_add_79_2_n346 ), .A2(_sha1_round_add_79_2_n34 ), .ZN(_sha1_round_add_79_2_n344 ) );
NOR2_X2 _sha1_round_add_79_2_U71  ( .A1(_sha1_round_add_79_2_n7 ), .A2(_sha1_round_add_79_2_n215 ), .ZN(_sha1_round_add_79_2_n216 ) );
NOR2_X2 _sha1_round_add_79_2_U70  ( .A1(_sha1_round_add_79_2_n59 ), .A2(_sha1_round_add_79_2_n33 ), .ZN(_sha1_round_add_79_2_n58 ) );
NOR2_X2 _sha1_round_add_79_2_U69  ( .A1(_sha1_round_add_79_2_n58 ), .A2(_sha1_round_add_79_2_n35 ), .ZN(_sha1_round_add_79_2_n54 ) );
AND3_X4 _sha1_round_add_79_2_U68  ( .A1(_sha1_round_add_79_2_n281 ), .A2(_sha1_round_add_79_2_n282 ), .A3(_sha1_round_add_79_2_n300 ), .ZN(_sha1_round_add_79_2_n24 ) );
AND2_X2 _sha1_round_add_79_2_U67  ( .A1(_sha1_round_add_79_2_n301 ), .A2(_sha1_round_add_79_2_n24 ), .ZN(_sha1_round_add_79_2_n261 ) );
NOR2_X2 _sha1_round_add_79_2_U66  ( .A1(_sha1_round_add_79_2_n76 ), .A2(_sha1_round_add_79_2_n368 ), .ZN(_sha1_round_add_79_2_n48 ) );
NOR2_X2 _sha1_round_add_79_2_U65  ( .A1(_sha1_round_add_79_2_n48 ), .A2(_sha1_round_add_79_2_n64 ), .ZN(_sha1_round_add_79_2_n79 ) );
NOR2_X2 _sha1_round_add_79_2_U64  ( .A1(_sha1_round_add_79_2_n79 ), .A2(_sha1_round_add_79_2_n75 ), .ZN(_sha1_round_add_79_2_n77 ) );
NOR2_X2 _sha1_round_add_79_2_U63  ( .A1(_sha1_round_add_79_2_n62 ), .A2(_sha1_round_add_79_2_n60 ), .ZN(_sha1_round_add_79_2_n78 ) );
NOR2_X2 _sha1_round_add_79_2_U62  ( .A1(_sha1_round_add_79_2_n36 ), .A2(_sha1_round_add_79_2_n85 ), .ZN(_sha1_round_add_79_2_n106 ) );
NAND3_X2 _sha1_round_add_79_2_U61  ( .A1(_sha1_round_add_79_2_n93 ), .A2(_sha1_round_add_79_2_n3 ), .A3(_sha1_round_add_79_2_n94 ), .ZN(_sha1_round_add_79_2_n92 ) );
NAND3_X2 _sha1_round_add_79_2_U60  ( .A1(_sha1_round_add_79_2_n330 ), .A2(_sha1_round_add_79_2_n322 ), .A3(_sha1_round_add_79_2_n10 ), .ZN(_sha1_round_add_79_2_n328 ) );
NAND3_X2 _sha1_round_add_79_2_U59  ( .A1(_sha1_round_add_79_2_n5 ), .A2(_sha1_round_add_79_2_n2 ), .A3(_sha1_round_add_79_2_n118 ), .ZN(_sha1_round_add_79_2_n171 ) );
NOR2_X2 _sha1_round_add_79_2_U58  ( .A1(_sha1_round_add_79_2_n64 ), .A2(_sha1_round_add_79_2_n65 ), .ZN(_sha1_round_add_79_2_n63 ) );
NOR2_X2 _sha1_round_add_79_2_U57  ( .A1(_sha1_round_add_79_2_n62 ), .A2(_sha1_round_add_79_2_n63 ), .ZN(_sha1_round_add_79_2_n59 ) );
NOR2_X2 _sha1_round_add_79_2_U56  ( .A1(_sha1_round_add_79_2_n197 ), .A2(_sha1_round_add_79_2_n188 ), .ZN(_sha1_round_add_79_2_n192 ) );
NOR2_X2 _sha1_round_add_79_2_U55  ( .A1(_sha1_round_add_79_2_n222 ), .A2(_sha1_round_add_79_2_n299 ), .ZN(_sha1_round_add_79_2_n297 ) );
NOR2_X2 _sha1_round_add_79_2_U54  ( .A1(_sha1_round_add_79_2_n119 ), .A2(_sha1_round_add_79_2_n8 ), .ZN(_sha1_round_add_79_2_n217 ) );
NOR2_X2 _sha1_round_add_79_2_U53  ( .A1(_sha1_round_add_79_2_n287 ), .A2(_sha1_round_add_79_2_n288 ), .ZN(_sha1_round_add_79_2_n255 ) );
NAND3_X2 _sha1_round_add_79_2_U52  ( .A1(_sha1_round_add_79_2_n255 ), .A2(_sha1_round_add_79_2_n12 ), .A3(_sha1_round_add_79_2_n256 ), .ZN(_sha1_round_add_79_2_n118 ) );
NOR2_X2 _sha1_round_add_79_2_U51  ( .A1(_sha1_round_add_79_2_n119 ), .A2(_sha1_round_add_79_2_n8 ), .ZN(_sha1_round_add_79_2_n116 ) );
NOR2_X2 _sha1_round_add_79_2_U50  ( .A1(_sha1_round_add_79_2_n64 ), .A2(_sha1_round_add_79_2_n75 ), .ZN(_sha1_round_add_79_2_n80 ) );
NOR2_X1 _sha1_round_add_79_2_U49  ( .A1(_sha1_round_add_79_2_n56 ), .A2(_sha1_round_add_79_2_n362 ), .ZN(_sha1_round_add_79_2_n276 ) );
OR2_X4 _sha1_round_add_79_2_U48  ( .A1(_sha1_round_add_79_2_n164 ), .A2(_sha1_round_add_79_2_n148 ), .ZN(_sha1_round_add_79_2_n23 ) );
NOR2_X2 _sha1_round_add_79_2_U47  ( .A1(_sha1_round_add_79_2_n167 ), .A2(_sha1_round_add_79_2_n168 ), .ZN(_sha1_round_add_79_2_n22 ) );
NOR2_X2 _sha1_round_add_79_2_U46  ( .A1(_sha1_round_add_79_2_n22 ), .A2(_sha1_round_add_79_2_n23 ), .ZN(_sha1_round_add_79_2_n162 ) );
AND2_X2 _sha1_round_add_79_2_U45  ( .A1(_sha1_round_add_79_2_n171 ), .A2(_sha1_round_add_79_2_n176 ), .ZN(_sha1_round_add_79_2_n21 ) );
OR2_X2 _sha1_round_add_79_2_U44  ( .A1(_sha1_round_add_79_2_n21 ), .A2(_sha1_round_add_79_2_n148 ), .ZN(_sha1_round_add_79_2_n174 ) );
NAND2_X2 _sha1_round_add_79_2_U43  ( .A1(_sha1_round_add_79_2_n300 ), .A2(_sha1_round_add_79_2_n281 ), .ZN(_sha1_round_add_79_2_n20 ) );
AND3_X4 _sha1_round_add_79_2_U42  ( .A1(_sha1_round_add_79_2_n292 ), .A2(_sha1_round_add_79_2_n279 ), .A3(_sha1_round_add_79_2_n307 ), .ZN(_sha1_round_add_79_2_n19 ) );
NOR2_X2 _sha1_round_add_79_2_U41  ( .A1(_sha1_round_add_79_2_n19 ), .A2(_sha1_round_add_79_2_n20 ), .ZN(_sha1_round_add_79_2_n305 ) );
NAND3_X1 _sha1_round_add_79_2_U40  ( .A1(_sha1_round_add_79_2_n261 ), .A2(_sha1_round_add_79_2_n285 ), .A3(_sha1_round_add_79_2_n286 ), .ZN(_sha1_round_add_79_2_n283 ) );
NOR2_X2 _sha1_round_add_79_2_U39  ( .A1(_sha1_round_add_79_2_n35 ), .A2(_sha1_round_add_79_2_n61 ), .ZN(_sha1_round_add_79_2_n18 ) );
XOR2_X2 _sha1_round_add_79_2_U38  ( .A(_sha1_round_add_79_2_n67 ), .B(_sha1_round_add_79_2_n18 ), .Z(_sha1_round_N290 ) );
NOR2_X1 _sha1_round_add_79_2_U37  ( .A1(_sha1_round_add_79_2_n215 ), .A2(_sha1_round_add_79_2_n197 ), .ZN(_sha1_round_add_79_2_n214 ) );
NOR2_X1 _sha1_round_add_79_2_U36  ( .A1(_sha1_round_add_79_2_n264 ), .A2(_sha1_round_add_79_2_n49 ), .ZN(_sha1_round_add_79_2_n317 ) );
NOR2_X1 _sha1_round_add_79_2_U35  ( .A1(_sha1_round_add_79_2_n264 ), .A2(_sha1_round_add_79_2_n72 ), .ZN(_sha1_round_add_79_2_n293 ) );
NAND3_X1 _sha1_round_add_79_2_U34  ( .A1(_sha1_round_add_79_2_n261 ), .A2(_sha1_round_add_79_2_n262 ), .A3(_sha1_round_add_79_2_n263 ), .ZN(_sha1_round_add_79_2_n260 ) );
NOR2_X1 _sha1_round_add_79_2_U33  ( .A1(_sha1_round_add_79_2_n264 ), .A2(_sha1_round_add_79_2_n265 ), .ZN(_sha1_round_add_79_2_n263 ) );
NOR2_X2 _sha1_round_add_79_2_U32  ( .A1(_sha1_round_add_79_2_n162 ), .A2(_sha1_round_add_79_2_n163 ), .ZN(_sha1_round_add_79_2_n17 ) );
XOR2_X2 _sha1_round_add_79_2_U31  ( .A(_sha1_round_add_79_2_n17 ), .B(_sha1_round_add_79_2_n159 ), .Z(_sha1_round_N310 ) );
NAND2_X1 _sha1_round_add_79_2_U30  ( .A1(_sha1_round_add_79_2_n171 ), .A2(_sha1_round_add_79_2_n180 ), .ZN(_sha1_round_add_79_2_n141 ) );
NOR2_X2 _sha1_round_add_79_2_U29  ( .A1(_sha1_round_add_79_2_n192 ), .A2(_sha1_round_add_79_2_n183 ), .ZN(_sha1_round_add_79_2_n16 ) );
XOR2_X2 _sha1_round_add_79_2_U28  ( .A(_sha1_round_add_79_2_n16 ), .B(_sha1_round_add_79_2_n189 ), .Z(_sha1_round_N307 ) );
NOR2_X2 _sha1_round_add_79_2_U27  ( .A1(_sha1_round_add_79_2_n84 ), .A2(_sha1_round_add_79_2_n36 ), .ZN(_sha1_round_add_79_2_n15 ) );
XOR2_X2 _sha1_round_add_79_2_U26  ( .A(_sha1_round_add_79_2_n15 ), .B(_sha1_round_add_79_2_n82 ), .Z(_sha1_round_N287 ) );
NOR2_X2 _sha1_round_add_79_2_U25  ( .A1(_sha1_round_add_79_2_n305 ), .A2(_sha1_round_add_79_2_n306 ), .ZN(_sha1_round_add_79_2_n14 ) );
XOR2_X2 _sha1_round_add_79_2_U24  ( .A(_sha1_round_add_79_2_n14 ), .B(_sha1_round_add_79_2_n302 ), .Z(_sha1_round_N299 ) );
NOR2_X1 _sha1_round_add_79_2_U23  ( .A1(_sha1_round_add_79_2_n340 ), .A2(_sha1_round_add_79_2_n37 ), .ZN(_sha1_round_add_79_2_n345 ) );
NOR2_X2 _sha1_round_add_79_2_U22  ( .A1(_sha1_round_add_79_2_n241 ), .A2(_sha1_round_add_79_2_n237 ), .ZN(_sha1_round_add_79_2_n13 ) );
XOR2_X2 _sha1_round_add_79_2_U21  ( .A(_sha1_round_add_79_2_n13 ), .B(_sha1_round_add_79_2_n238 ), .Z(_sha1_round_N302 ) );
NAND3_X1 _sha1_round_add_79_2_U20  ( .A1(_sha1_round_add_79_2_n360 ), .A2(_sha1_round_add_79_2_n262 ), .A3(_sha1_round_add_79_2_n361 ), .ZN(_sha1_round_add_79_2_n359 ) );
NOR2_X1 _sha1_round_add_79_2_U19  ( .A1(_sha1_round_add_79_2_n56 ), .A2(_sha1_round_add_79_2_n57 ), .ZN(_sha1_round_add_79_2_n55 ) );
NOR2_X1 _sha1_round_add_79_2_U18  ( .A1(_sha1_round_add_79_2_n321 ), .A2(_sha1_round_add_79_2_n264 ), .ZN(_sha1_round_add_79_2_n320 ) );
NOR2_X1 _sha1_round_add_79_2_U17  ( .A1(_sha1_round_add_79_2_n264 ), .A2(_sha1_round_add_79_2_n275 ), .ZN(_sha1_round_add_79_2_n274 ) );
NAND2_X1 _sha1_round_add_79_2_U16  ( .A1(_sha1_round_add_79_2_n5 ), .A2(_sha1_round_add_79_2_n118 ), .ZN(_sha1_round_add_79_2_n218 ) );
NAND2_X1 _sha1_round_add_79_2_U15  ( .A1(_sha1_round_add_79_2_n5 ), .A2(_sha1_round_add_79_2_n118 ), .ZN(_sha1_round_add_79_2_n117 ) );
NAND3_X2 _sha1_round_add_79_2_U14  ( .A1(_sha1_round_add_79_2_n363 ), .A2(_sha1_round_add_79_2_n71 ), .A3(_sha1_round_add_79_2_n364 ), .ZN(_sha1_round_add_79_2_n49 ) );
AND2_X4 _sha1_round_add_79_2_U13  ( .A1(_sha1_round_add_79_2_n283 ), .A2(_sha1_round_add_79_2_n284 ), .ZN(_sha1_round_add_79_2_n12 ) );
OR2_X4 _sha1_round_add_79_2_U12  ( .A1(rnd_q[21]), .A2(w[21]), .ZN(_sha1_round_add_79_2_n11 ) );
OR2_X4 _sha1_round_add_79_2_U11  ( .A1(_sha1_round_add_79_2_n48 ), .A2(_sha1_round_add_79_2_n331 ), .ZN(_sha1_round_add_79_2_n10 ) );
AND2_X4 _sha1_round_add_79_2_U10  ( .A1(w[30]), .A2(rnd_q[30]), .ZN(_sha1_round_add_79_2_n9 ) );
AND2_X4 _sha1_round_add_79_2_U9  ( .A1(_sha1_round_add_79_2_n185 ), .A2(_sha1_round_add_79_2_n186 ), .ZN(_sha1_round_add_79_2_n8 ) );
AND2_X4 _sha1_round_add_79_2_U8  ( .A1(w[20]), .A2(rnd_q[20]), .ZN(_sha1_round_add_79_2_n7 ) );
AND2_X4 _sha1_round_add_79_2_U7  ( .A1(w[25]), .A2(rnd_q[25]), .ZN(_sha1_round_add_79_2_n6 ) );
AND2_X4 _sha1_round_add_79_2_U6  ( .A1(_sha1_round_add_79_2_n219 ), .A2(_sha1_round_add_79_2_n186 ), .ZN(_sha1_round_add_79_2_n5 ) );
AND2_X4 _sha1_round_add_79_2_U5  ( .A1(_sha1_round_add_79_2_n101 ), .A2(_sha1_round_add_79_2_n102 ), .ZN(_sha1_round_add_79_2_n4 ) );
AND2_X4 _sha1_round_add_79_2_U4  ( .A1(_sha1_round_add_79_2_n2 ), .A2(_sha1_round_add_79_2_n115 ), .ZN(_sha1_round_add_79_2_n3 ) );
AND2_X4 _sha1_round_add_79_2_U3  ( .A1(_sha1_round_add_79_2_n187 ), .A2(_sha1_round_add_79_2_n184 ), .ZN(_sha1_round_add_79_2_n2 ) );
AND2_X4 _sha1_round_add_79_2_U2  ( .A1(_sha1_round_add_79_2_n120 ), .A2(_sha1_round_add_79_2_n115 ), .ZN(_sha1_round_add_79_2_n1 ) );
AND2_X2 _rnd_cnt_reg_U15  ( .A1(rnd_cnt_d[6]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N9 ) );
AND2_X2 _rnd_cnt_reg_U14  ( .A1(rnd_cnt_d[5]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N8 ) );
AND2_X2 _rnd_cnt_reg_U13  ( .A1(rnd_cnt_d[4]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N7 ) );
AND2_X2 _rnd_cnt_reg_U12  ( .A1(rnd_cnt_d[3]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N6 ) );
INV_X4 _rnd_cnt_reg_U11  ( .A(_rnd_cnt_reg_n70 ), .ZN(rnd_cnt_q[2]) );
INV_X4 _rnd_cnt_reg_U10  ( .A(_rnd_cnt_reg_n40 ), .ZN(rnd_cnt_q[3]) );
INV_X1 _rnd_cnt_reg_U7  ( .A(n7117), .ZN(_rnd_cnt_reg_n12 ) );
AND2_X4 _rnd_cnt_reg_U6  ( .A1(rnd_cnt_d[2]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N5 ) );
INV_X4 _rnd_cnt_reg_U5  ( .A(_rnd_cnt_reg_n60 ), .ZN(rnd_cnt_q[5]) );
INV_X4 _rnd_cnt_reg_U4  ( .A(_rnd_cnt_reg_n2 ), .ZN(rnd_cnt_q[6]) );
INV_X8 _rnd_cnt_reg_U3  ( .A(_rnd_cnt_reg_n10 ), .ZN(rnd_cnt_q[4]) );
DFF_X2 _rnd_cnt_reg_q_reg_5_  ( .D(_rnd_cnt_reg_N8 ), .CK(clk), .Q(), .QN(_rnd_cnt_reg_n60 ) );
DFF_X2 _rnd_cnt_reg_q_reg_4_  ( .D(_rnd_cnt_reg_N7 ), .CK(clk), .Q(), .QN(_rnd_cnt_reg_n10 ) );
DFF_X1 _rnd_cnt_reg_q_reg_6_  ( .D(_rnd_cnt_reg_N9 ), .CK(clk), .Q(), .QN(_rnd_cnt_reg_n2 ) );
DFF_X2 _rnd_cnt_reg_q_reg_2_  ( .D(_rnd_cnt_reg_N5 ), .CK(clk), .Q(), .QN(_rnd_cnt_reg_n70 ) );
AND2_X2 _rnd_cnt_reg_U9  ( .A1(rnd_cnt_d[0]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N3 ) );
AND2_X2 _rnd_cnt_reg_U8  ( .A1(rnd_cnt_d[1]), .A2(_rnd_cnt_reg_n12 ), .ZN(_rnd_cnt_reg_N4 ) );
DFF_X2 _rnd_cnt_reg_q_reg_0_  ( .D(_rnd_cnt_reg_N3 ), .CK(clk), .Q(rnd_cnt_q[0]), .QN() );
DFF_X2 _rnd_cnt_reg_q_reg_1_  ( .D(_rnd_cnt_reg_N4 ), .CK(clk), .Q(rnd_cnt_q[1]), .QN() );
DFF_X2 _rnd_cnt_reg_q_reg_3_  ( .D(_rnd_cnt_reg_N6 ), .CK(clk), .Q(), .QN(_rnd_cnt_reg_n40 ) );
INV_X4 _state_reg_U5  ( .A(n7117), .ZN(_state_reg_n2 ) );
AND2_X4 _state_reg_U3  ( .A1(next_state[1]), .A2(_state_reg_n2 ), .ZN(_state_reg_N4 ) );
AND2_X2 _state_reg_U4  ( .A1(next_state[0]), .A2(_state_reg_n2 ), .ZN(_state_reg_N3 ) );
DFF_X2 _state_reg_q_reg_0_  ( .D(_state_reg_N3 ), .CK(clk), .Q(state[0]),.QN() );
DFF_X2 _state_reg_q_reg_1_  ( .D(_state_reg_N4 ), .CK(clk), .Q(state[1]),.QN() );
AND2_X2 _w_reg_U562  ( .A1(w_d[497]), .A2(_w_reg_n610 ), .ZN(_w_reg_N500 ));
AND2_X2 _w_reg_U561  ( .A1(w_d[496]), .A2(_w_reg_n610 ), .ZN(_w_reg_N499 ));
AND2_X2 _w_reg_U560  ( .A1(w_d[495]), .A2(_w_reg_n610 ), .ZN(_w_reg_N498 ));
AND2_X2 _w_reg_U559  ( .A1(w_d[494]), .A2(_w_reg_n610 ), .ZN(_w_reg_N497 ));
AND2_X2 _w_reg_U558  ( .A1(w_d[493]), .A2(_w_reg_n610 ), .ZN(_w_reg_N496 ));
AND2_X2 _w_reg_U557  ( .A1(w_d[492]), .A2(_w_reg_n610 ), .ZN(_w_reg_N495 ));
AND2_X2 _w_reg_U556  ( .A1(w_d[491]), .A2(_w_reg_n610 ), .ZN(_w_reg_N494 ));
AND2_X2 _w_reg_U555  ( .A1(w_d[490]), .A2(_w_reg_n600 ), .ZN(_w_reg_N493 ));
AND2_X2 _w_reg_U554  ( .A1(w_d[489]), .A2(_w_reg_n600 ), .ZN(_w_reg_N492 ));
AND2_X2 _w_reg_U553  ( .A1(w_d[488]), .A2(_w_reg_n600 ), .ZN(_w_reg_N491 ));
AND2_X2 _w_reg_U552  ( .A1(w_d[487]), .A2(_w_reg_n600 ), .ZN(_w_reg_N490 ));
AND2_X2 _w_reg_U551  ( .A1(w_d[486]), .A2(_w_reg_n600 ), .ZN(_w_reg_N489 ));
AND2_X2 _w_reg_U550  ( .A1(w_d[485]), .A2(_w_reg_n600 ), .ZN(_w_reg_N488 ));
AND2_X2 _w_reg_U549  ( .A1(w_d[484]), .A2(_w_reg_n600 ), .ZN(_w_reg_N487 ));
AND2_X2 _w_reg_U548  ( .A1(w_d[483]), .A2(_w_reg_n600 ), .ZN(_w_reg_N486 ));
AND2_X2 _w_reg_U547  ( .A1(w_d[482]), .A2(_w_reg_n600 ), .ZN(_w_reg_N485 ));
AND2_X2 _w_reg_U546  ( .A1(w_d[481]), .A2(_w_reg_n600 ), .ZN(_w_reg_N484 ));
AND2_X2 _w_reg_U545  ( .A1(w_d[480]), .A2(_w_reg_n600 ), .ZN(_w_reg_N483 ));
INV_X4 _w_reg_U544  ( .A(reset), .ZN(_w_reg_n1070 ) );
BUF_X4 _w_reg_U543  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1060 ) );
BUF_X4 _w_reg_U542  ( .A(_w_reg_n1070 ), .Z(_w_reg_n660 ) );
BUF_X4 _w_reg_U541  ( .A(_w_reg_n1070 ), .Z(_w_reg_n670 ) );
BUF_X4 _w_reg_U540  ( .A(_w_reg_n1070 ), .Z(_w_reg_n610 ) );
BUF_X4 _w_reg_U539  ( .A(_w_reg_n1070 ), .Z(_w_reg_n600 ) );
BUF_X4 _w_reg_U538  ( .A(_w_reg_n1070 ), .Z(_w_reg_n680 ) );
BUF_X4 _w_reg_U537  ( .A(_w_reg_n1070 ), .Z(_w_reg_n690 ) );
BUF_X4 _w_reg_U536  ( .A(_w_reg_n1070 ), .Z(_w_reg_n700 ) );
BUF_X4 _w_reg_U535  ( .A(_w_reg_n1070 ), .Z(_w_reg_n710 ) );
BUF_X4 _w_reg_U534  ( .A(_w_reg_n1070 ), .Z(_w_reg_n720 ) );
BUF_X4 _w_reg_U533  ( .A(_w_reg_n1070 ), .Z(_w_reg_n730 ) );
BUF_X4 _w_reg_U532  ( .A(_w_reg_n1070 ), .Z(_w_reg_n740 ) );
BUF_X4 _w_reg_U531  ( .A(_w_reg_n1070 ), .Z(_w_reg_n750 ) );
BUF_X4 _w_reg_U530  ( .A(_w_reg_n1070 ), .Z(_w_reg_n760 ) );
BUF_X4 _w_reg_U529  ( .A(_w_reg_n1070 ), .Z(_w_reg_n770 ) );
BUF_X4 _w_reg_U528  ( .A(_w_reg_n1070 ), .Z(_w_reg_n780 ) );
BUF_X4 _w_reg_U527  ( .A(_w_reg_n1070 ), .Z(_w_reg_n790 ) );
BUF_X4 _w_reg_U526  ( .A(_w_reg_n1070 ), .Z(_w_reg_n800 ) );
BUF_X4 _w_reg_U525  ( .A(_w_reg_n1070 ), .Z(_w_reg_n810 ) );
BUF_X4 _w_reg_U524  ( .A(_w_reg_n1070 ), .Z(_w_reg_n820 ) );
BUF_X4 _w_reg_U523  ( .A(_w_reg_n1070 ), .Z(_w_reg_n830 ) );
BUF_X4 _w_reg_U522  ( .A(_w_reg_n1070 ), .Z(_w_reg_n840 ) );
BUF_X4 _w_reg_U521  ( .A(_w_reg_n1070 ), .Z(_w_reg_n850 ) );
BUF_X4 _w_reg_U520  ( .A(_w_reg_n1070 ), .Z(_w_reg_n860 ) );
BUF_X4 _w_reg_U519  ( .A(_w_reg_n1070 ), .Z(_w_reg_n870 ) );
BUF_X4 _w_reg_U518  ( .A(_w_reg_n1070 ), .Z(_w_reg_n880 ) );
BUF_X4 _w_reg_U517  ( .A(_w_reg_n1070 ), .Z(_w_reg_n890 ) );
BUF_X4 _w_reg_U516  ( .A(_w_reg_n1070 ), .Z(_w_reg_n900 ) );
BUF_X4 _w_reg_U515  ( .A(_w_reg_n1070 ), .Z(_w_reg_n910 ) );
BUF_X4 _w_reg_U514  ( .A(_w_reg_n1070 ), .Z(_w_reg_n920 ) );
BUF_X4 _w_reg_U503  ( .A(_w_reg_n1070 ), .Z(_w_reg_n930 ) );
BUF_X4 _w_reg_U492  ( .A(_w_reg_n1070 ), .Z(_w_reg_n940 ) );
BUF_X4 _w_reg_U481  ( .A(_w_reg_n1070 ), .Z(_w_reg_n950 ) );
BUF_X4 _w_reg_U470  ( .A(_w_reg_n1070 ), .Z(_w_reg_n960 ) );
BUF_X4 _w_reg_U459  ( .A(_w_reg_n1070 ), .Z(_w_reg_n970 ) );
BUF_X4 _w_reg_U448  ( .A(_w_reg_n1070 ), .Z(_w_reg_n980 ) );
BUF_X4 _w_reg_U437  ( .A(_w_reg_n1070 ), .Z(_w_reg_n990 ) );
BUF_X4 _w_reg_U426  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1000 ) );
BUF_X4 _w_reg_U415  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1010 ) );
BUF_X4 _w_reg_U404  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1020 ) );
BUF_X4 _w_reg_U393  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1030 ) );
BUF_X4 _w_reg_U382  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1040 ) );
BUF_X4 _w_reg_U371  ( .A(_w_reg_n1070 ), .Z(_w_reg_n1050 ) );
BUF_X4 _w_reg_U360  ( .A(_w_reg_n1070 ), .Z(_w_reg_n620 ) );
BUF_X4 _w_reg_U349  ( .A(_w_reg_n1070 ), .Z(_w_reg_n630 ) );
BUF_X4 _w_reg_U338  ( .A(_w_reg_n1070 ), .Z(_w_reg_n640 ) );
BUF_X4 _w_reg_U327  ( .A(_w_reg_n1070 ), .Z(_w_reg_n650 ) );
AND2_X1 _w_reg_U316  ( .A1(w_d[31]), .A2(_w_reg_n820 ), .ZN(_w_reg_N34 ) );
AND2_X1 _w_reg_U305  ( .A1(w_d[30]), .A2(_w_reg_n830 ), .ZN(_w_reg_N33 ) );
AND2_X1 _w_reg_U294  ( .A1(w_d[29]), .A2(_w_reg_n840 ), .ZN(_w_reg_N32 ) );
AND2_X1 _w_reg_U293  ( .A1(w_d[28]), .A2(_w_reg_n850 ), .ZN(_w_reg_N31 ) );
AND2_X1 _w_reg_U282  ( .A1(w_d[27]), .A2(_w_reg_n860 ), .ZN(_w_reg_N30 ) );
AND2_X1 _w_reg_U271  ( .A1(w_d[26]), .A2(_w_reg_n870 ), .ZN(_w_reg_N29 ) );
AND2_X1 _w_reg_U260  ( .A1(w_d[25]), .A2(_w_reg_n880 ), .ZN(_w_reg_N28 ) );
AND2_X1 _w_reg_U249  ( .A1(w_d[24]), .A2(_w_reg_n890 ), .ZN(_w_reg_N27 ) );
AND2_X1 _w_reg_U183  ( .A1(w_d[23]), .A2(_w_reg_n900 ), .ZN(_w_reg_N26 ) );
AND2_X1 _w_reg_U90  ( .A1(w_d[22]), .A2(_w_reg_n910 ), .ZN(_w_reg_N25 ) );
AND2_X1 _w_reg_U89  ( .A1(w_d[21]), .A2(_w_reg_n920 ), .ZN(_w_reg_N24 ) );
AND2_X1 _w_reg_U88  ( .A1(w_d[20]), .A2(_w_reg_n930 ), .ZN(_w_reg_N23 ) );
AND2_X1 _w_reg_U87  ( .A1(w_d[19]), .A2(_w_reg_n940 ), .ZN(_w_reg_N22 ) );
AND2_X1 _w_reg_U86  ( .A1(w_d[18]), .A2(_w_reg_n950 ), .ZN(_w_reg_N21 ) );
AND2_X1 _w_reg_U85  ( .A1(w_d[17]), .A2(_w_reg_n960 ), .ZN(_w_reg_N20 ) );
AND2_X1 _w_reg_U84  ( .A1(w_d[16]), .A2(_w_reg_n970 ), .ZN(_w_reg_N19 ) );
AND2_X1 _w_reg_U82  ( .A1(w_d[15]), .A2(_w_reg_n980 ), .ZN(_w_reg_N18 ) );
AND2_X1 _w_reg_U81  ( .A1(w_d[14]), .A2(_w_reg_n990 ), .ZN(_w_reg_N17 ) );
AND2_X1 _w_reg_U80  ( .A1(w_d[13]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N16 ) );
AND2_X1 _w_reg_U79  ( .A1(w_d[12]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N15 ) );
AND2_X1 _w_reg_U78  ( .A1(w_d[11]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N14 ) );
AND2_X1 _w_reg_U77  ( .A1(w_d[10]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N13 ) );
AND2_X1 _w_reg_U76  ( .A1(w_d[9]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N12 ) );
AND2_X1 _w_reg_U75  ( .A1(w_d[8]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N11 ) );
AND2_X1 _w_reg_U74  ( .A1(w_d[7]), .A2(_w_reg_n1060 ), .ZN(_w_reg_N10 ) );
AND2_X1 _w_reg_U73  ( .A1(w_d[6]), .A2(_w_reg_n620 ), .ZN(_w_reg_N9 ) );
AND2_X1 _w_reg_U72  ( .A1(w_d[5]), .A2(_w_reg_n630 ), .ZN(_w_reg_N8 ) );
AND2_X1 _w_reg_U70  ( .A1(w_d[4]), .A2(_w_reg_n640 ), .ZN(_w_reg_N7 ) );
AND2_X1 _w_reg_U46  ( .A1(w_d[3]), .A2(_w_reg_n650 ), .ZN(_w_reg_N6 ) );
AND2_X1 _w_reg_U35  ( .A1(w_d[2]), .A2(_w_reg_n670 ), .ZN(_w_reg_N5 ) );
AND2_X1 _w_reg_U24  ( .A1(w_d[1]), .A2(_w_reg_n760 ), .ZN(_w_reg_N4 ) );
AND2_X1 _w_reg_U13  ( .A1(w_d[0]), .A2(_w_reg_n860 ), .ZN(_w_reg_N3 ) );
AND2_X2 _w_reg_U513  ( .A1(w_d[97]), .A2(_w_reg_n1060 ), .ZN(_w_reg_N100 ));
AND2_X2 _w_reg_U512  ( .A1(w_d[98]), .A2(_w_reg_n1060 ), .ZN(_w_reg_N101 ));
AND2_X2 _w_reg_U511  ( .A1(w_d[99]), .A2(_w_reg_n1060 ), .ZN(_w_reg_N102 ));
AND2_X2 _w_reg_U510  ( .A1(w_d[100]), .A2(_w_reg_n1060 ), .ZN(_w_reg_N103 ));
AND2_X2 _w_reg_U509  ( .A1(w_d[101]), .A2(_w_reg_n1060 ), .ZN(_w_reg_N104 ));
AND2_X2 _w_reg_U508  ( .A1(w_d[102]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N105 ));
AND2_X2 _w_reg_U507  ( .A1(w_d[103]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N106 ));
AND2_X2 _w_reg_U506  ( .A1(w_d[104]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N107 ));
AND2_X2 _w_reg_U505  ( .A1(w_d[105]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N108 ));
AND2_X2 _w_reg_U504  ( .A1(w_d[106]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N109 ));
AND2_X2 _w_reg_U502  ( .A1(w_d[107]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N110 ));
AND2_X2 _w_reg_U501  ( .A1(w_d[108]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N111 ));
AND2_X2 _w_reg_U500  ( .A1(w_d[109]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N112 ));
AND2_X2 _w_reg_U499  ( .A1(w_d[110]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N113 ));
AND2_X2 _w_reg_U498  ( .A1(w_d[111]), .A2(_w_reg_n1050 ), .ZN(_w_reg_N114 ));
AND2_X2 _w_reg_U497  ( .A1(w_d[112]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N115 ));
AND2_X2 _w_reg_U496  ( .A1(w_d[113]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N116 ));
AND2_X2 _w_reg_U495  ( .A1(w_d[114]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N117 ));
AND2_X2 _w_reg_U494  ( .A1(w_d[115]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N118 ));
AND2_X2 _w_reg_U493  ( .A1(w_d[116]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N119 ));
AND2_X2 _w_reg_U491  ( .A1(w_d[117]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N120 ));
AND2_X2 _w_reg_U490  ( .A1(w_d[118]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N121 ));
AND2_X2 _w_reg_U489  ( .A1(w_d[119]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N122 ));
AND2_X2 _w_reg_U488  ( .A1(w_d[120]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N123 ));
AND2_X2 _w_reg_U487  ( .A1(w_d[121]), .A2(_w_reg_n1040 ), .ZN(_w_reg_N124 ));
AND2_X2 _w_reg_U486  ( .A1(w_d[122]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N125 ));
AND2_X2 _w_reg_U485  ( .A1(w_d[123]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N126 ));
AND2_X2 _w_reg_U484  ( .A1(w_d[124]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N127 ));
AND2_X2 _w_reg_U483  ( .A1(w_d[125]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N128 ));
AND2_X2 _w_reg_U482  ( .A1(w_d[126]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N129 ));
AND2_X2 _w_reg_U480  ( .A1(w_d[127]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N130 ));
AND2_X2 _w_reg_U479  ( .A1(w_d[128]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N131 ));
AND2_X2 _w_reg_U478  ( .A1(w_d[129]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N132 ));
AND2_X2 _w_reg_U477  ( .A1(w_d[130]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N133 ));
AND2_X2 _w_reg_U476  ( .A1(w_d[131]), .A2(_w_reg_n1030 ), .ZN(_w_reg_N134 ));
AND2_X2 _w_reg_U475  ( .A1(w_d[132]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N135 ));
AND2_X2 _w_reg_U474  ( .A1(w_d[133]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N136 ));
AND2_X2 _w_reg_U473  ( .A1(w_d[134]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N137 ));
AND2_X2 _w_reg_U472  ( .A1(w_d[135]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N138 ));
AND2_X2 _w_reg_U471  ( .A1(w_d[136]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N139 ));
AND2_X2 _w_reg_U469  ( .A1(w_d[137]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N140 ));
AND2_X2 _w_reg_U468  ( .A1(w_d[138]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N141 ));
AND2_X2 _w_reg_U467  ( .A1(w_d[139]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N142 ));
AND2_X2 _w_reg_U466  ( .A1(w_d[140]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N143 ));
AND2_X2 _w_reg_U465  ( .A1(w_d[141]), .A2(_w_reg_n1020 ), .ZN(_w_reg_N144 ));
AND2_X2 _w_reg_U464  ( .A1(w_d[142]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N145 ));
AND2_X2 _w_reg_U463  ( .A1(w_d[143]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N146 ));
AND2_X2 _w_reg_U462  ( .A1(w_d[144]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N147 ));
AND2_X2 _w_reg_U461  ( .A1(w_d[145]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N148 ));
AND2_X2 _w_reg_U460  ( .A1(w_d[146]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N149 ));
AND2_X2 _w_reg_U458  ( .A1(w_d[147]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N150 ));
AND2_X2 _w_reg_U457  ( .A1(w_d[148]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N151 ));
AND2_X2 _w_reg_U456  ( .A1(w_d[149]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N152 ));
AND2_X2 _w_reg_U455  ( .A1(w_d[150]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N153 ));
AND2_X2 _w_reg_U454  ( .A1(w_d[151]), .A2(_w_reg_n1010 ), .ZN(_w_reg_N154 ));
AND2_X2 _w_reg_U453  ( .A1(w_d[152]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N155 ));
AND2_X2 _w_reg_U452  ( .A1(w_d[153]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N156 ));
AND2_X2 _w_reg_U451  ( .A1(w_d[154]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N157 ));
AND2_X2 _w_reg_U450  ( .A1(w_d[155]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N158 ));
AND2_X2 _w_reg_U449  ( .A1(w_d[156]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N159 ));
AND2_X2 _w_reg_U447  ( .A1(w_d[157]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N160 ));
AND2_X2 _w_reg_U446  ( .A1(w_d[158]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N161 ));
AND2_X2 _w_reg_U445  ( .A1(w_d[159]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N162 ));
AND2_X2 _w_reg_U444  ( .A1(w_d[160]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N163 ));
AND2_X2 _w_reg_U443  ( .A1(w_d[161]), .A2(_w_reg_n1000 ), .ZN(_w_reg_N164 ));
AND2_X2 _w_reg_U442  ( .A1(w_d[162]), .A2(_w_reg_n990 ), .ZN(_w_reg_N165 ));
AND2_X2 _w_reg_U441  ( .A1(w_d[163]), .A2(_w_reg_n990 ), .ZN(_w_reg_N166 ));
AND2_X2 _w_reg_U440  ( .A1(w_d[164]), .A2(_w_reg_n990 ), .ZN(_w_reg_N167 ));
AND2_X2 _w_reg_U439  ( .A1(w_d[165]), .A2(_w_reg_n990 ), .ZN(_w_reg_N168 ));
AND2_X2 _w_reg_U438  ( .A1(w_d[166]), .A2(_w_reg_n990 ), .ZN(_w_reg_N169 ));
AND2_X2 _w_reg_U436  ( .A1(w_d[167]), .A2(_w_reg_n990 ), .ZN(_w_reg_N170 ));
AND2_X2 _w_reg_U435  ( .A1(w_d[168]), .A2(_w_reg_n990 ), .ZN(_w_reg_N171 ));
AND2_X2 _w_reg_U434  ( .A1(w_d[169]), .A2(_w_reg_n990 ), .ZN(_w_reg_N172 ));
AND2_X2 _w_reg_U433  ( .A1(w_d[170]), .A2(_w_reg_n990 ), .ZN(_w_reg_N173 ));
AND2_X2 _w_reg_U432  ( .A1(w_d[171]), .A2(_w_reg_n990 ), .ZN(_w_reg_N174 ));
AND2_X2 _w_reg_U431  ( .A1(w_d[172]), .A2(_w_reg_n980 ), .ZN(_w_reg_N175 ));
AND2_X2 _w_reg_U430  ( .A1(w_d[173]), .A2(_w_reg_n980 ), .ZN(_w_reg_N176 ));
AND2_X2 _w_reg_U429  ( .A1(w_d[174]), .A2(_w_reg_n980 ), .ZN(_w_reg_N177 ));
AND2_X2 _w_reg_U428  ( .A1(w_d[175]), .A2(_w_reg_n980 ), .ZN(_w_reg_N178 ));
AND2_X2 _w_reg_U427  ( .A1(w_d[176]), .A2(_w_reg_n980 ), .ZN(_w_reg_N179 ));
AND2_X2 _w_reg_U425  ( .A1(w_d[177]), .A2(_w_reg_n980 ), .ZN(_w_reg_N180 ));
AND2_X2 _w_reg_U424  ( .A1(w_d[178]), .A2(_w_reg_n980 ), .ZN(_w_reg_N181 ));
AND2_X2 _w_reg_U423  ( .A1(w_d[179]), .A2(_w_reg_n980 ), .ZN(_w_reg_N182 ));
AND2_X2 _w_reg_U422  ( .A1(w_d[180]), .A2(_w_reg_n980 ), .ZN(_w_reg_N183 ));
AND2_X2 _w_reg_U421  ( .A1(w_d[181]), .A2(_w_reg_n980 ), .ZN(_w_reg_N184 ));
AND2_X2 _w_reg_U420  ( .A1(w_d[182]), .A2(_w_reg_n970 ), .ZN(_w_reg_N185 ));
AND2_X2 _w_reg_U419  ( .A1(w_d[183]), .A2(_w_reg_n970 ), .ZN(_w_reg_N186 ));
AND2_X2 _w_reg_U418  ( .A1(w_d[184]), .A2(_w_reg_n970 ), .ZN(_w_reg_N187 ));
AND2_X2 _w_reg_U417  ( .A1(w_d[185]), .A2(_w_reg_n970 ), .ZN(_w_reg_N188 ));
AND2_X2 _w_reg_U416  ( .A1(w_d[186]), .A2(_w_reg_n970 ), .ZN(_w_reg_N189 ));
AND2_X2 _w_reg_U414  ( .A1(w_d[187]), .A2(_w_reg_n970 ), .ZN(_w_reg_N190 ));
AND2_X2 _w_reg_U413  ( .A1(w_d[188]), .A2(_w_reg_n970 ), .ZN(_w_reg_N191 ));
AND2_X2 _w_reg_U412  ( .A1(w_d[189]), .A2(_w_reg_n970 ), .ZN(_w_reg_N192 ));
AND2_X2 _w_reg_U411  ( .A1(w_d[190]), .A2(_w_reg_n970 ), .ZN(_w_reg_N193 ));
AND2_X2 _w_reg_U410  ( .A1(w_d[191]), .A2(_w_reg_n970 ), .ZN(_w_reg_N194 ));
AND2_X2 _w_reg_U409  ( .A1(w_d[192]), .A2(_w_reg_n960 ), .ZN(_w_reg_N195 ));
AND2_X2 _w_reg_U408  ( .A1(w_d[193]), .A2(_w_reg_n960 ), .ZN(_w_reg_N196 ));
AND2_X2 _w_reg_U407  ( .A1(w_d[194]), .A2(_w_reg_n960 ), .ZN(_w_reg_N197 ));
AND2_X2 _w_reg_U406  ( .A1(w_d[195]), .A2(_w_reg_n960 ), .ZN(_w_reg_N198 ));
AND2_X2 _w_reg_U405  ( .A1(w_d[196]), .A2(_w_reg_n960 ), .ZN(_w_reg_N199 ));
AND2_X2 _w_reg_U403  ( .A1(w_d[197]), .A2(_w_reg_n960 ), .ZN(_w_reg_N200 ));
AND2_X2 _w_reg_U402  ( .A1(w_d[198]), .A2(_w_reg_n960 ), .ZN(_w_reg_N201 ));
AND2_X2 _w_reg_U401  ( .A1(w_d[199]), .A2(_w_reg_n960 ), .ZN(_w_reg_N202 ));
AND2_X2 _w_reg_U400  ( .A1(w_d[200]), .A2(_w_reg_n960 ), .ZN(_w_reg_N203 ));
AND2_X2 _w_reg_U399  ( .A1(w_d[201]), .A2(_w_reg_n960 ), .ZN(_w_reg_N204 ));
AND2_X2 _w_reg_U398  ( .A1(w_d[202]), .A2(_w_reg_n950 ), .ZN(_w_reg_N205 ));
AND2_X2 _w_reg_U397  ( .A1(w_d[203]), .A2(_w_reg_n950 ), .ZN(_w_reg_N206 ));
AND2_X2 _w_reg_U396  ( .A1(w_d[204]), .A2(_w_reg_n950 ), .ZN(_w_reg_N207 ));
AND2_X2 _w_reg_U395  ( .A1(w_d[205]), .A2(_w_reg_n950 ), .ZN(_w_reg_N208 ));
AND2_X2 _w_reg_U394  ( .A1(w_d[206]), .A2(_w_reg_n950 ), .ZN(_w_reg_N209 ));
AND2_X2 _w_reg_U392  ( .A1(w_d[207]), .A2(_w_reg_n950 ), .ZN(_w_reg_N210 ));
AND2_X2 _w_reg_U391  ( .A1(w_d[208]), .A2(_w_reg_n950 ), .ZN(_w_reg_N211 ));
AND2_X2 _w_reg_U390  ( .A1(w_d[209]), .A2(_w_reg_n950 ), .ZN(_w_reg_N212 ));
AND2_X2 _w_reg_U389  ( .A1(w_d[210]), .A2(_w_reg_n950 ), .ZN(_w_reg_N213 ));
AND2_X2 _w_reg_U388  ( .A1(w_d[211]), .A2(_w_reg_n950 ), .ZN(_w_reg_N214 ));
AND2_X2 _w_reg_U387  ( .A1(w_d[212]), .A2(_w_reg_n940 ), .ZN(_w_reg_N215 ));
AND2_X2 _w_reg_U386  ( .A1(w_d[213]), .A2(_w_reg_n940 ), .ZN(_w_reg_N216 ));
AND2_X2 _w_reg_U385  ( .A1(w_d[214]), .A2(_w_reg_n940 ), .ZN(_w_reg_N217 ));
AND2_X2 _w_reg_U384  ( .A1(w_d[215]), .A2(_w_reg_n940 ), .ZN(_w_reg_N218 ));
AND2_X2 _w_reg_U383  ( .A1(w_d[216]), .A2(_w_reg_n940 ), .ZN(_w_reg_N219 ));
AND2_X2 _w_reg_U381  ( .A1(w_d[217]), .A2(_w_reg_n940 ), .ZN(_w_reg_N220 ));
AND2_X2 _w_reg_U380  ( .A1(w_d[218]), .A2(_w_reg_n940 ), .ZN(_w_reg_N221 ));
AND2_X2 _w_reg_U379  ( .A1(w_d[219]), .A2(_w_reg_n940 ), .ZN(_w_reg_N222 ));
AND2_X2 _w_reg_U378  ( .A1(w_d[220]), .A2(_w_reg_n940 ), .ZN(_w_reg_N223 ));
AND2_X2 _w_reg_U377  ( .A1(w_d[221]), .A2(_w_reg_n940 ), .ZN(_w_reg_N224 ));
AND2_X2 _w_reg_U376  ( .A1(w_d[222]), .A2(_w_reg_n930 ), .ZN(_w_reg_N225 ));
AND2_X2 _w_reg_U375  ( .A1(w_d[223]), .A2(_w_reg_n930 ), .ZN(_w_reg_N226 ));
AND2_X2 _w_reg_U374  ( .A1(w_d[224]), .A2(_w_reg_n930 ), .ZN(_w_reg_N227 ));
AND2_X2 _w_reg_U373  ( .A1(w_d[225]), .A2(_w_reg_n930 ), .ZN(_w_reg_N228 ));
AND2_X2 _w_reg_U372  ( .A1(w_d[226]), .A2(_w_reg_n930 ), .ZN(_w_reg_N229 ));
AND2_X2 _w_reg_U370  ( .A1(w_d[227]), .A2(_w_reg_n930 ), .ZN(_w_reg_N230 ));
AND2_X2 _w_reg_U369  ( .A1(w_d[228]), .A2(_w_reg_n930 ), .ZN(_w_reg_N231 ));
AND2_X2 _w_reg_U368  ( .A1(w_d[229]), .A2(_w_reg_n930 ), .ZN(_w_reg_N232 ));
AND2_X2 _w_reg_U367  ( .A1(w_d[230]), .A2(_w_reg_n930 ), .ZN(_w_reg_N233 ));
AND2_X2 _w_reg_U366  ( .A1(w_d[231]), .A2(_w_reg_n930 ), .ZN(_w_reg_N234 ));
AND2_X2 _w_reg_U365  ( .A1(w_d[232]), .A2(_w_reg_n920 ), .ZN(_w_reg_N235 ));
AND2_X2 _w_reg_U364  ( .A1(w_d[233]), .A2(_w_reg_n920 ), .ZN(_w_reg_N236 ));
AND2_X2 _w_reg_U363  ( .A1(w_d[234]), .A2(_w_reg_n920 ), .ZN(_w_reg_N237 ));
AND2_X2 _w_reg_U362  ( .A1(w_d[235]), .A2(_w_reg_n920 ), .ZN(_w_reg_N238 ));
AND2_X2 _w_reg_U361  ( .A1(w_d[236]), .A2(_w_reg_n920 ), .ZN(_w_reg_N239 ));
AND2_X2 _w_reg_U359  ( .A1(w_d[237]), .A2(_w_reg_n920 ), .ZN(_w_reg_N240 ));
AND2_X2 _w_reg_U358  ( .A1(w_d[238]), .A2(_w_reg_n920 ), .ZN(_w_reg_N241 ));
AND2_X2 _w_reg_U357  ( .A1(w_d[239]), .A2(_w_reg_n920 ), .ZN(_w_reg_N242 ));
AND2_X2 _w_reg_U356  ( .A1(w_d[240]), .A2(_w_reg_n920 ), .ZN(_w_reg_N243 ));
AND2_X2 _w_reg_U355  ( .A1(w_d[241]), .A2(_w_reg_n920 ), .ZN(_w_reg_N244 ));
AND2_X2 _w_reg_U354  ( .A1(w_d[242]), .A2(_w_reg_n910 ), .ZN(_w_reg_N245 ));
AND2_X2 _w_reg_U353  ( .A1(w_d[243]), .A2(_w_reg_n910 ), .ZN(_w_reg_N246 ));
AND2_X2 _w_reg_U352  ( .A1(w_d[244]), .A2(_w_reg_n910 ), .ZN(_w_reg_N247 ));
AND2_X2 _w_reg_U351  ( .A1(w_d[245]), .A2(_w_reg_n910 ), .ZN(_w_reg_N248 ));
AND2_X2 _w_reg_U350  ( .A1(w_d[246]), .A2(_w_reg_n910 ), .ZN(_w_reg_N249 ));
AND2_X2 _w_reg_U348  ( .A1(w_d[247]), .A2(_w_reg_n910 ), .ZN(_w_reg_N250 ));
AND2_X2 _w_reg_U347  ( .A1(w_d[248]), .A2(_w_reg_n910 ), .ZN(_w_reg_N251 ));
AND2_X2 _w_reg_U346  ( .A1(w_d[249]), .A2(_w_reg_n910 ), .ZN(_w_reg_N252 ));
AND2_X2 _w_reg_U345  ( .A1(w_d[250]), .A2(_w_reg_n910 ), .ZN(_w_reg_N253 ));
AND2_X2 _w_reg_U344  ( .A1(w_d[251]), .A2(_w_reg_n910 ), .ZN(_w_reg_N254 ));
AND2_X2 _w_reg_U343  ( .A1(w_d[252]), .A2(_w_reg_n900 ), .ZN(_w_reg_N255 ));
AND2_X2 _w_reg_U342  ( .A1(w_d[253]), .A2(_w_reg_n900 ), .ZN(_w_reg_N256 ));
AND2_X2 _w_reg_U341  ( .A1(w_d[254]), .A2(_w_reg_n900 ), .ZN(_w_reg_N257 ));
AND2_X2 _w_reg_U340  ( .A1(w_d[255]), .A2(_w_reg_n900 ), .ZN(_w_reg_N258 ));
AND2_X2 _w_reg_U339  ( .A1(w_d[256]), .A2(_w_reg_n900 ), .ZN(_w_reg_N259 ));
AND2_X2 _w_reg_U337  ( .A1(w_d[257]), .A2(_w_reg_n900 ), .ZN(_w_reg_N260 ));
AND2_X2 _w_reg_U336  ( .A1(w_d[258]), .A2(_w_reg_n900 ), .ZN(_w_reg_N261 ));
AND2_X2 _w_reg_U335  ( .A1(w_d[259]), .A2(_w_reg_n900 ), .ZN(_w_reg_N262 ));
AND2_X2 _w_reg_U334  ( .A1(w_d[260]), .A2(_w_reg_n900 ), .ZN(_w_reg_N263 ));
AND2_X2 _w_reg_U333  ( .A1(w_d[261]), .A2(_w_reg_n900 ), .ZN(_w_reg_N264 ));
AND2_X2 _w_reg_U332  ( .A1(w_d[262]), .A2(_w_reg_n890 ), .ZN(_w_reg_N265 ));
AND2_X2 _w_reg_U331  ( .A1(w_d[263]), .A2(_w_reg_n890 ), .ZN(_w_reg_N266 ));
AND2_X2 _w_reg_U330  ( .A1(w_d[264]), .A2(_w_reg_n890 ), .ZN(_w_reg_N267 ));
AND2_X2 _w_reg_U329  ( .A1(w_d[265]), .A2(_w_reg_n890 ), .ZN(_w_reg_N268 ));
AND2_X2 _w_reg_U328  ( .A1(w_d[266]), .A2(_w_reg_n890 ), .ZN(_w_reg_N269 ));
AND2_X2 _w_reg_U326  ( .A1(w_d[267]), .A2(_w_reg_n890 ), .ZN(_w_reg_N270 ));
AND2_X2 _w_reg_U325  ( .A1(w_d[268]), .A2(_w_reg_n890 ), .ZN(_w_reg_N271 ));
AND2_X2 _w_reg_U324  ( .A1(w_d[269]), .A2(_w_reg_n890 ), .ZN(_w_reg_N272 ));
AND2_X2 _w_reg_U323  ( .A1(w_d[270]), .A2(_w_reg_n890 ), .ZN(_w_reg_N273 ));
AND2_X2 _w_reg_U322  ( .A1(w_d[271]), .A2(_w_reg_n890 ), .ZN(_w_reg_N274 ));
AND2_X2 _w_reg_U321  ( .A1(w_d[272]), .A2(_w_reg_n880 ), .ZN(_w_reg_N275 ));
AND2_X2 _w_reg_U320  ( .A1(w_d[273]), .A2(_w_reg_n880 ), .ZN(_w_reg_N276 ));
AND2_X2 _w_reg_U319  ( .A1(w_d[274]), .A2(_w_reg_n880 ), .ZN(_w_reg_N277 ));
AND2_X2 _w_reg_U318  ( .A1(w_d[275]), .A2(_w_reg_n880 ), .ZN(_w_reg_N278 ));
AND2_X2 _w_reg_U317  ( .A1(w_d[276]), .A2(_w_reg_n880 ), .ZN(_w_reg_N279 ));
AND2_X2 _w_reg_U315  ( .A1(w_d[277]), .A2(_w_reg_n880 ), .ZN(_w_reg_N280 ));
AND2_X2 _w_reg_U314  ( .A1(w_d[278]), .A2(_w_reg_n880 ), .ZN(_w_reg_N281 ));
AND2_X2 _w_reg_U313  ( .A1(w_d[279]), .A2(_w_reg_n880 ), .ZN(_w_reg_N282 ));
AND2_X2 _w_reg_U312  ( .A1(w_d[280]), .A2(_w_reg_n880 ), .ZN(_w_reg_N283 ));
AND2_X2 _w_reg_U311  ( .A1(w_d[281]), .A2(_w_reg_n880 ), .ZN(_w_reg_N284 ));
AND2_X2 _w_reg_U310  ( .A1(w_d[282]), .A2(_w_reg_n870 ), .ZN(_w_reg_N285 ));
AND2_X2 _w_reg_U309  ( .A1(w_d[283]), .A2(_w_reg_n870 ), .ZN(_w_reg_N286 ));
AND2_X2 _w_reg_U308  ( .A1(w_d[284]), .A2(_w_reg_n870 ), .ZN(_w_reg_N287 ));
AND2_X2 _w_reg_U307  ( .A1(w_d[285]), .A2(_w_reg_n870 ), .ZN(_w_reg_N288 ));
AND2_X2 _w_reg_U306  ( .A1(w_d[286]), .A2(_w_reg_n870 ), .ZN(_w_reg_N289 ));
AND2_X2 _w_reg_U304  ( .A1(w_d[287]), .A2(_w_reg_n870 ), .ZN(_w_reg_N290 ));
AND2_X2 _w_reg_U303  ( .A1(w_d[288]), .A2(_w_reg_n870 ), .ZN(_w_reg_N291 ));
AND2_X2 _w_reg_U302  ( .A1(w_d[289]), .A2(_w_reg_n870 ), .ZN(_w_reg_N292 ));
AND2_X2 _w_reg_U301  ( .A1(w_d[290]), .A2(_w_reg_n870 ), .ZN(_w_reg_N293 ));
AND2_X2 _w_reg_U300  ( .A1(w_d[291]), .A2(_w_reg_n870 ), .ZN(_w_reg_N294 ));
AND2_X2 _w_reg_U299  ( .A1(w_d[292]), .A2(_w_reg_n860 ), .ZN(_w_reg_N295 ));
AND2_X2 _w_reg_U298  ( .A1(w_d[293]), .A2(_w_reg_n860 ), .ZN(_w_reg_N296 ));
AND2_X2 _w_reg_U297  ( .A1(w_d[294]), .A2(_w_reg_n860 ), .ZN(_w_reg_N297 ));
AND2_X2 _w_reg_U296  ( .A1(w_d[295]), .A2(_w_reg_n860 ), .ZN(_w_reg_N298 ));
AND2_X2 _w_reg_U295  ( .A1(w_d[296]), .A2(_w_reg_n860 ), .ZN(_w_reg_N299 ));
AND2_X2 _w_reg_U292  ( .A1(w_d[297]), .A2(_w_reg_n860 ), .ZN(_w_reg_N300 ));
AND2_X2 _w_reg_U291  ( .A1(w_d[298]), .A2(_w_reg_n860 ), .ZN(_w_reg_N301 ));
AND2_X2 _w_reg_U290  ( .A1(w_d[299]), .A2(_w_reg_n860 ), .ZN(_w_reg_N302 ));
AND2_X2 _w_reg_U289  ( .A1(w_d[300]), .A2(_w_reg_n860 ), .ZN(_w_reg_N303 ));
AND2_X2 _w_reg_U288  ( .A1(w_d[301]), .A2(_w_reg_n850 ), .ZN(_w_reg_N304 ));
AND2_X2 _w_reg_U287  ( .A1(w_d[302]), .A2(_w_reg_n850 ), .ZN(_w_reg_N305 ));
AND2_X2 _w_reg_U286  ( .A1(w_d[303]), .A2(_w_reg_n850 ), .ZN(_w_reg_N306 ));
AND2_X2 _w_reg_U285  ( .A1(w_d[304]), .A2(_w_reg_n850 ), .ZN(_w_reg_N307 ));
AND2_X2 _w_reg_U284  ( .A1(w_d[305]), .A2(_w_reg_n850 ), .ZN(_w_reg_N308 ));
AND2_X2 _w_reg_U283  ( .A1(w_d[306]), .A2(_w_reg_n850 ), .ZN(_w_reg_N309 ));
AND2_X2 _w_reg_U281  ( .A1(w_d[307]), .A2(_w_reg_n850 ), .ZN(_w_reg_N310 ));
AND2_X2 _w_reg_U280  ( .A1(w_d[308]), .A2(_w_reg_n850 ), .ZN(_w_reg_N311 ));
AND2_X2 _w_reg_U279  ( .A1(w_d[309]), .A2(_w_reg_n850 ), .ZN(_w_reg_N312 ));
AND2_X2 _w_reg_U278  ( .A1(w_d[310]), .A2(_w_reg_n850 ), .ZN(_w_reg_N313 ));
AND2_X2 _w_reg_U277  ( .A1(w_d[311]), .A2(_w_reg_n840 ), .ZN(_w_reg_N314 ));
AND2_X2 _w_reg_U276  ( .A1(w_d[312]), .A2(_w_reg_n840 ), .ZN(_w_reg_N315 ));
AND2_X2 _w_reg_U275  ( .A1(w_d[313]), .A2(_w_reg_n840 ), .ZN(_w_reg_N316 ));
AND2_X2 _w_reg_U274  ( .A1(w_d[314]), .A2(_w_reg_n840 ), .ZN(_w_reg_N317 ));
AND2_X2 _w_reg_U273  ( .A1(w_d[315]), .A2(_w_reg_n840 ), .ZN(_w_reg_N318 ));
AND2_X2 _w_reg_U272  ( .A1(w_d[316]), .A2(_w_reg_n840 ), .ZN(_w_reg_N319 ));
AND2_X2 _w_reg_U270  ( .A1(w_d[317]), .A2(_w_reg_n840 ), .ZN(_w_reg_N320 ));
AND2_X2 _w_reg_U269  ( .A1(w_d[318]), .A2(_w_reg_n840 ), .ZN(_w_reg_N321 ));
AND2_X2 _w_reg_U268  ( .A1(w_d[319]), .A2(_w_reg_n840 ), .ZN(_w_reg_N322 ));
AND2_X2 _w_reg_U267  ( .A1(w_d[320]), .A2(_w_reg_n840 ), .ZN(_w_reg_N323 ));
AND2_X2 _w_reg_U266  ( .A1(w_d[321]), .A2(_w_reg_n830 ), .ZN(_w_reg_N324 ));
AND2_X2 _w_reg_U265  ( .A1(w_d[322]), .A2(_w_reg_n830 ), .ZN(_w_reg_N325 ));
AND2_X2 _w_reg_U264  ( .A1(w_d[323]), .A2(_w_reg_n830 ), .ZN(_w_reg_N326 ));
AND2_X2 _w_reg_U263  ( .A1(w_d[324]), .A2(_w_reg_n830 ), .ZN(_w_reg_N327 ));
AND2_X2 _w_reg_U262  ( .A1(w_d[325]), .A2(_w_reg_n830 ), .ZN(_w_reg_N328 ));
AND2_X2 _w_reg_U261  ( .A1(w_d[326]), .A2(_w_reg_n830 ), .ZN(_w_reg_N329 ));
AND2_X2 _w_reg_U259  ( .A1(w_d[327]), .A2(_w_reg_n830 ), .ZN(_w_reg_N330 ));
AND2_X2 _w_reg_U258  ( .A1(w_d[328]), .A2(_w_reg_n830 ), .ZN(_w_reg_N331 ));
AND2_X2 _w_reg_U257  ( .A1(w_d[329]), .A2(_w_reg_n830 ), .ZN(_w_reg_N332 ));
AND2_X2 _w_reg_U256  ( .A1(w_d[330]), .A2(_w_reg_n830 ), .ZN(_w_reg_N333 ));
AND2_X2 _w_reg_U255  ( .A1(w_d[331]), .A2(_w_reg_n820 ), .ZN(_w_reg_N334 ));
AND2_X2 _w_reg_U254  ( .A1(w_d[332]), .A2(_w_reg_n820 ), .ZN(_w_reg_N335 ));
AND2_X2 _w_reg_U253  ( .A1(w_d[333]), .A2(_w_reg_n820 ), .ZN(_w_reg_N336 ));
AND2_X2 _w_reg_U252  ( .A1(w_d[334]), .A2(_w_reg_n820 ), .ZN(_w_reg_N337 ));
AND2_X2 _w_reg_U251  ( .A1(w_d[335]), .A2(_w_reg_n820 ), .ZN(_w_reg_N338 ));
AND2_X2 _w_reg_U250  ( .A1(w_d[336]), .A2(_w_reg_n820 ), .ZN(_w_reg_N339 ));
AND2_X2 _w_reg_U248  ( .A1(w_d[337]), .A2(_w_reg_n820 ), .ZN(_w_reg_N340 ));
AND2_X2 _w_reg_U247  ( .A1(w_d[338]), .A2(_w_reg_n820 ), .ZN(_w_reg_N341 ));
AND2_X2 _w_reg_U246  ( .A1(w_d[339]), .A2(_w_reg_n820 ), .ZN(_w_reg_N342 ));
AND2_X2 _w_reg_U245  ( .A1(w_d[340]), .A2(_w_reg_n820 ), .ZN(_w_reg_N343 ));
AND2_X2 _w_reg_U244  ( .A1(w_d[341]), .A2(_w_reg_n810 ), .ZN(_w_reg_N344 ));
AND2_X2 _w_reg_U243  ( .A1(w_d[342]), .A2(_w_reg_n810 ), .ZN(_w_reg_N345 ));
AND2_X2 _w_reg_U242  ( .A1(w_d[343]), .A2(_w_reg_n810 ), .ZN(_w_reg_N346 ));
AND2_X2 _w_reg_U241  ( .A1(w_d[344]), .A2(_w_reg_n810 ), .ZN(_w_reg_N347 ));
AND2_X2 _w_reg_U240  ( .A1(w_d[345]), .A2(_w_reg_n810 ), .ZN(_w_reg_N348 ));
AND2_X2 _w_reg_U239  ( .A1(w_d[346]), .A2(_w_reg_n810 ), .ZN(_w_reg_N349 ));
AND2_X2 _w_reg_U238  ( .A1(w_d[32]), .A2(_w_reg_n810 ), .ZN(_w_reg_N35 ) );
AND2_X2 _w_reg_U237  ( .A1(w_d[347]), .A2(_w_reg_n810 ), .ZN(_w_reg_N350 ));
AND2_X2 _w_reg_U236  ( .A1(w_d[348]), .A2(_w_reg_n810 ), .ZN(_w_reg_N351 ));
AND2_X2 _w_reg_U235  ( .A1(w_d[349]), .A2(_w_reg_n810 ), .ZN(_w_reg_N352 ));
AND2_X2 _w_reg_U234  ( .A1(w_d[350]), .A2(_w_reg_n810 ), .ZN(_w_reg_N353 ));
AND2_X2 _w_reg_U233  ( .A1(w_d[351]), .A2(_w_reg_n800 ), .ZN(_w_reg_N354 ));
AND2_X2 _w_reg_U232  ( .A1(w_d[352]), .A2(_w_reg_n800 ), .ZN(_w_reg_N355 ));
AND2_X2 _w_reg_U231  ( .A1(w_d[353]), .A2(_w_reg_n800 ), .ZN(_w_reg_N356 ));
AND2_X2 _w_reg_U230  ( .A1(w_d[354]), .A2(_w_reg_n800 ), .ZN(_w_reg_N357 ));
AND2_X2 _w_reg_U229  ( .A1(w_d[355]), .A2(_w_reg_n800 ), .ZN(_w_reg_N358 ));
AND2_X2 _w_reg_U228  ( .A1(w_d[356]), .A2(_w_reg_n800 ), .ZN(_w_reg_N359 ));
AND2_X2 _w_reg_U227  ( .A1(w_d[33]), .A2(_w_reg_n800 ), .ZN(_w_reg_N36 ) );
AND2_X2 _w_reg_U226  ( .A1(w_d[357]), .A2(_w_reg_n800 ), .ZN(_w_reg_N360 ));
AND2_X2 _w_reg_U225  ( .A1(w_d[358]), .A2(_w_reg_n800 ), .ZN(_w_reg_N361 ));
AND2_X2 _w_reg_U224  ( .A1(w_d[359]), .A2(_w_reg_n800 ), .ZN(_w_reg_N362 ));
AND2_X2 _w_reg_U223  ( .A1(w_d[360]), .A2(_w_reg_n800 ), .ZN(_w_reg_N363 ));
AND2_X2 _w_reg_U222  ( .A1(w_d[361]), .A2(_w_reg_n790 ), .ZN(_w_reg_N364 ));
AND2_X2 _w_reg_U221  ( .A1(w_d[362]), .A2(_w_reg_n790 ), .ZN(_w_reg_N365 ));
AND2_X2 _w_reg_U220  ( .A1(w_d[363]), .A2(_w_reg_n790 ), .ZN(_w_reg_N366 ));
AND2_X2 _w_reg_U219  ( .A1(w_d[364]), .A2(_w_reg_n790 ), .ZN(_w_reg_N367 ));
AND2_X2 _w_reg_U218  ( .A1(w_d[365]), .A2(_w_reg_n790 ), .ZN(_w_reg_N368 ));
AND2_X2 _w_reg_U217  ( .A1(w_d[366]), .A2(_w_reg_n790 ), .ZN(_w_reg_N369 ));
AND2_X2 _w_reg_U216  ( .A1(w_d[34]), .A2(_w_reg_n790 ), .ZN(_w_reg_N37 ) );
AND2_X2 _w_reg_U215  ( .A1(w_d[367]), .A2(_w_reg_n790 ), .ZN(_w_reg_N370 ));
AND2_X2 _w_reg_U214  ( .A1(w_d[368]), .A2(_w_reg_n790 ), .ZN(_w_reg_N371 ));
AND2_X2 _w_reg_U213  ( .A1(w_d[369]), .A2(_w_reg_n790 ), .ZN(_w_reg_N372 ));
AND2_X2 _w_reg_U212  ( .A1(w_d[370]), .A2(_w_reg_n790 ), .ZN(_w_reg_N373 ));
AND2_X2 _w_reg_U211  ( .A1(w_d[371]), .A2(_w_reg_n780 ), .ZN(_w_reg_N374 ));
AND2_X2 _w_reg_U210  ( .A1(w_d[372]), .A2(_w_reg_n780 ), .ZN(_w_reg_N375 ));
AND2_X2 _w_reg_U209  ( .A1(w_d[373]), .A2(_w_reg_n780 ), .ZN(_w_reg_N376 ));
AND2_X2 _w_reg_U208  ( .A1(w_d[374]), .A2(_w_reg_n780 ), .ZN(_w_reg_N377 ));
AND2_X2 _w_reg_U207  ( .A1(w_d[375]), .A2(_w_reg_n780 ), .ZN(_w_reg_N378 ));
AND2_X2 _w_reg_U206  ( .A1(w_d[376]), .A2(_w_reg_n780 ), .ZN(_w_reg_N379 ));
AND2_X2 _w_reg_U205  ( .A1(w_d[35]), .A2(_w_reg_n780 ), .ZN(_w_reg_N38 ) );
AND2_X2 _w_reg_U204  ( .A1(w_d[377]), .A2(_w_reg_n780 ), .ZN(_w_reg_N380 ));
AND2_X2 _w_reg_U203  ( .A1(w_d[378]), .A2(_w_reg_n780 ), .ZN(_w_reg_N381 ));
AND2_X2 _w_reg_U202  ( .A1(w_d[379]), .A2(_w_reg_n780 ), .ZN(_w_reg_N382 ));
AND2_X2 _w_reg_U201  ( .A1(w_d[380]), .A2(_w_reg_n780 ), .ZN(_w_reg_N383 ));
AND2_X2 _w_reg_U200  ( .A1(w_d[381]), .A2(_w_reg_n770 ), .ZN(_w_reg_N384 ));
AND2_X2 _w_reg_U199  ( .A1(w_d[382]), .A2(_w_reg_n770 ), .ZN(_w_reg_N385 ));
AND2_X2 _w_reg_U198  ( .A1(w_d[383]), .A2(_w_reg_n770 ), .ZN(_w_reg_N386 ));
AND2_X2 _w_reg_U197  ( .A1(w_d[384]), .A2(_w_reg_n770 ), .ZN(_w_reg_N387 ));
AND2_X2 _w_reg_U196  ( .A1(w_d[385]), .A2(_w_reg_n770 ), .ZN(_w_reg_N388 ));
AND2_X2 _w_reg_U195  ( .A1(w_d[386]), .A2(_w_reg_n770 ), .ZN(_w_reg_N389 ));
AND2_X2 _w_reg_U194  ( .A1(w_d[36]), .A2(_w_reg_n770 ), .ZN(_w_reg_N39 ) );
AND2_X2 _w_reg_U193  ( .A1(w_d[387]), .A2(_w_reg_n770 ), .ZN(_w_reg_N390 ));
AND2_X2 _w_reg_U192  ( .A1(w_d[388]), .A2(_w_reg_n770 ), .ZN(_w_reg_N391 ));
AND2_X2 _w_reg_U191  ( .A1(w_d[389]), .A2(_w_reg_n770 ), .ZN(_w_reg_N392 ));
AND2_X2 _w_reg_U190  ( .A1(w_d[390]), .A2(_w_reg_n770 ), .ZN(_w_reg_N393 ));
AND2_X2 _w_reg_U189  ( .A1(w_d[391]), .A2(_w_reg_n760 ), .ZN(_w_reg_N394 ));
AND2_X2 _w_reg_U188  ( .A1(w_d[392]), .A2(_w_reg_n760 ), .ZN(_w_reg_N395 ));
AND2_X2 _w_reg_U187  ( .A1(w_d[393]), .A2(_w_reg_n760 ), .ZN(_w_reg_N396 ));
AND2_X2 _w_reg_U186  ( .A1(w_d[394]), .A2(_w_reg_n760 ), .ZN(_w_reg_N397 ));
AND2_X2 _w_reg_U185  ( .A1(w_d[395]), .A2(_w_reg_n760 ), .ZN(_w_reg_N398 ));
AND2_X2 _w_reg_U184  ( .A1(w_d[396]), .A2(_w_reg_n760 ), .ZN(_w_reg_N399 ));
AND2_X2 _w_reg_U182  ( .A1(w_d[37]), .A2(_w_reg_n760 ), .ZN(_w_reg_N40 ) );
AND2_X2 _w_reg_U181  ( .A1(w_d[397]), .A2(_w_reg_n760 ), .ZN(_w_reg_N400 ));
AND2_X2 _w_reg_U180  ( .A1(w_d[398]), .A2(_w_reg_n760 ), .ZN(_w_reg_N401 ));
AND2_X2 _w_reg_U179  ( .A1(w_d[399]), .A2(_w_reg_n760 ), .ZN(_w_reg_N402 ));
AND2_X2 _w_reg_U178  ( .A1(w_d[400]), .A2(_w_reg_n750 ), .ZN(_w_reg_N403 ));
AND2_X2 _w_reg_U177  ( .A1(w_d[401]), .A2(_w_reg_n750 ), .ZN(_w_reg_N404 ));
AND2_X2 _w_reg_U176  ( .A1(w_d[402]), .A2(_w_reg_n750 ), .ZN(_w_reg_N405 ));
AND2_X2 _w_reg_U175  ( .A1(w_d[403]), .A2(_w_reg_n750 ), .ZN(_w_reg_N406 ));
AND2_X2 _w_reg_U174  ( .A1(w_d[404]), .A2(_w_reg_n750 ), .ZN(_w_reg_N407 ));
AND2_X2 _w_reg_U173  ( .A1(w_d[405]), .A2(_w_reg_n750 ), .ZN(_w_reg_N408 ));
AND2_X2 _w_reg_U172  ( .A1(w_d[406]), .A2(_w_reg_n750 ), .ZN(_w_reg_N409 ));
AND2_X2 _w_reg_U171  ( .A1(w_d[38]), .A2(_w_reg_n750 ), .ZN(_w_reg_N41 ) );
AND2_X2 _w_reg_U170  ( .A1(w_d[407]), .A2(_w_reg_n750 ), .ZN(_w_reg_N410 ));
AND2_X2 _w_reg_U169  ( .A1(w_d[408]), .A2(_w_reg_n750 ), .ZN(_w_reg_N411 ));
AND2_X2 _w_reg_U168  ( .A1(w_d[409]), .A2(_w_reg_n750 ), .ZN(_w_reg_N412 ));
AND2_X2 _w_reg_U167  ( .A1(w_d[410]), .A2(_w_reg_n740 ), .ZN(_w_reg_N413 ));
AND2_X2 _w_reg_U166  ( .A1(w_d[411]), .A2(_w_reg_n740 ), .ZN(_w_reg_N414 ));
AND2_X2 _w_reg_U165  ( .A1(w_d[412]), .A2(_w_reg_n740 ), .ZN(_w_reg_N415 ));
AND2_X2 _w_reg_U164  ( .A1(w_d[413]), .A2(_w_reg_n740 ), .ZN(_w_reg_N416 ));
AND2_X2 _w_reg_U163  ( .A1(w_d[414]), .A2(_w_reg_n740 ), .ZN(_w_reg_N417 ));
AND2_X2 _w_reg_U162  ( .A1(w_d[415]), .A2(_w_reg_n740 ), .ZN(_w_reg_N418 ));
AND2_X2 _w_reg_U161  ( .A1(w_d[416]), .A2(_w_reg_n740 ), .ZN(_w_reg_N419 ));
AND2_X2 _w_reg_U160  ( .A1(w_d[39]), .A2(_w_reg_n740 ), .ZN(_w_reg_N42 ) );
AND2_X2 _w_reg_U159  ( .A1(w_d[417]), .A2(_w_reg_n740 ), .ZN(_w_reg_N420 ));
AND2_X2 _w_reg_U158  ( .A1(w_d[418]), .A2(_w_reg_n740 ), .ZN(_w_reg_N421 ));
AND2_X2 _w_reg_U157  ( .A1(w_d[419]), .A2(_w_reg_n740 ), .ZN(_w_reg_N422 ));
AND2_X2 _w_reg_U156  ( .A1(w_d[420]), .A2(_w_reg_n730 ), .ZN(_w_reg_N423 ));
AND2_X2 _w_reg_U155  ( .A1(w_d[421]), .A2(_w_reg_n730 ), .ZN(_w_reg_N424 ));
AND2_X2 _w_reg_U154  ( .A1(w_d[422]), .A2(_w_reg_n730 ), .ZN(_w_reg_N425 ));
AND2_X2 _w_reg_U153  ( .A1(w_d[423]), .A2(_w_reg_n730 ), .ZN(_w_reg_N426 ));
AND2_X2 _w_reg_U152  ( .A1(w_d[424]), .A2(_w_reg_n730 ), .ZN(_w_reg_N427 ));
AND2_X2 _w_reg_U151  ( .A1(w_d[425]), .A2(_w_reg_n730 ), .ZN(_w_reg_N428 ));
AND2_X2 _w_reg_U150  ( .A1(w_d[426]), .A2(_w_reg_n730 ), .ZN(_w_reg_N429 ));
AND2_X2 _w_reg_U149  ( .A1(w_d[40]), .A2(_w_reg_n730 ), .ZN(_w_reg_N43 ) );
AND2_X2 _w_reg_U148  ( .A1(w_d[427]), .A2(_w_reg_n730 ), .ZN(_w_reg_N430 ));
AND2_X2 _w_reg_U147  ( .A1(w_d[428]), .A2(_w_reg_n730 ), .ZN(_w_reg_N431 ));
AND2_X2 _w_reg_U146  ( .A1(w_d[429]), .A2(_w_reg_n730 ), .ZN(_w_reg_N432 ));
AND2_X2 _w_reg_U145  ( .A1(w_d[430]), .A2(_w_reg_n720 ), .ZN(_w_reg_N433 ));
AND2_X2 _w_reg_U144  ( .A1(w_d[431]), .A2(_w_reg_n720 ), .ZN(_w_reg_N434 ));
AND2_X2 _w_reg_U143  ( .A1(w_d[432]), .A2(_w_reg_n720 ), .ZN(_w_reg_N435 ));
AND2_X2 _w_reg_U142  ( .A1(w_d[433]), .A2(_w_reg_n720 ), .ZN(_w_reg_N436 ));
AND2_X2 _w_reg_U141  ( .A1(w_d[434]), .A2(_w_reg_n720 ), .ZN(_w_reg_N437 ));
AND2_X2 _w_reg_U140  ( .A1(w_d[435]), .A2(_w_reg_n720 ), .ZN(_w_reg_N438 ));
AND2_X2 _w_reg_U139  ( .A1(w_d[436]), .A2(_w_reg_n720 ), .ZN(_w_reg_N439 ));
AND2_X2 _w_reg_U138  ( .A1(w_d[41]), .A2(_w_reg_n720 ), .ZN(_w_reg_N44 ) );
AND2_X2 _w_reg_U137  ( .A1(w_d[437]), .A2(_w_reg_n720 ), .ZN(_w_reg_N440 ));
AND2_X2 _w_reg_U136  ( .A1(w_d[438]), .A2(_w_reg_n720 ), .ZN(_w_reg_N441 ));
AND2_X2 _w_reg_U135  ( .A1(w_d[439]), .A2(_w_reg_n720 ), .ZN(_w_reg_N442 ));
AND2_X2 _w_reg_U134  ( .A1(w_d[440]), .A2(_w_reg_n710 ), .ZN(_w_reg_N443 ));
AND2_X2 _w_reg_U133  ( .A1(w_d[441]), .A2(_w_reg_n710 ), .ZN(_w_reg_N444 ));
AND2_X2 _w_reg_U132  ( .A1(w_d[442]), .A2(_w_reg_n710 ), .ZN(_w_reg_N445 ));
AND2_X2 _w_reg_U131  ( .A1(w_d[443]), .A2(_w_reg_n710 ), .ZN(_w_reg_N446 ));
AND2_X2 _w_reg_U130  ( .A1(w_d[444]), .A2(_w_reg_n710 ), .ZN(_w_reg_N447 ));
AND2_X2 _w_reg_U129  ( .A1(w_d[445]), .A2(_w_reg_n710 ), .ZN(_w_reg_N448 ));
AND2_X2 _w_reg_U128  ( .A1(w_d[446]), .A2(_w_reg_n710 ), .ZN(_w_reg_N449 ));
AND2_X2 _w_reg_U127  ( .A1(w_d[42]), .A2(_w_reg_n710 ), .ZN(_w_reg_N45 ) );
AND2_X2 _w_reg_U126  ( .A1(w_d[447]), .A2(_w_reg_n710 ), .ZN(_w_reg_N450 ));
AND2_X2 _w_reg_U125  ( .A1(w_d[448]), .A2(_w_reg_n710 ), .ZN(_w_reg_N451 ));
AND2_X2 _w_reg_U124  ( .A1(w_d[449]), .A2(_w_reg_n710 ), .ZN(_w_reg_N452 ));
AND2_X2 _w_reg_U123  ( .A1(w_d[450]), .A2(_w_reg_n700 ), .ZN(_w_reg_N453 ));
AND2_X2 _w_reg_U122  ( .A1(w_d[451]), .A2(_w_reg_n700 ), .ZN(_w_reg_N454 ));
AND2_X2 _w_reg_U121  ( .A1(w_d[452]), .A2(_w_reg_n700 ), .ZN(_w_reg_N455 ));
AND2_X2 _w_reg_U120  ( .A1(w_d[453]), .A2(_w_reg_n700 ), .ZN(_w_reg_N456 ));
AND2_X2 _w_reg_U119  ( .A1(w_d[454]), .A2(_w_reg_n700 ), .ZN(_w_reg_N457 ));
AND2_X2 _w_reg_U118  ( .A1(w_d[455]), .A2(_w_reg_n700 ), .ZN(_w_reg_N458 ));
AND2_X2 _w_reg_U117  ( .A1(w_d[456]), .A2(_w_reg_n700 ), .ZN(_w_reg_N459 ));
AND2_X2 _w_reg_U116  ( .A1(w_d[43]), .A2(_w_reg_n700 ), .ZN(_w_reg_N46 ) );
AND2_X2 _w_reg_U115  ( .A1(w_d[457]), .A2(_w_reg_n700 ), .ZN(_w_reg_N460 ));
AND2_X2 _w_reg_U114  ( .A1(w_d[458]), .A2(_w_reg_n700 ), .ZN(_w_reg_N461 ));
AND2_X2 _w_reg_U113  ( .A1(w_d[459]), .A2(_w_reg_n700 ), .ZN(_w_reg_N462 ));
AND2_X2 _w_reg_U112  ( .A1(w_d[460]), .A2(_w_reg_n690 ), .ZN(_w_reg_N463 ));
AND2_X2 _w_reg_U111  ( .A1(w_d[461]), .A2(_w_reg_n690 ), .ZN(_w_reg_N464 ));
AND2_X2 _w_reg_U110  ( .A1(w_d[462]), .A2(_w_reg_n690 ), .ZN(_w_reg_N465 ));
AND2_X2 _w_reg_U109  ( .A1(w_d[463]), .A2(_w_reg_n690 ), .ZN(_w_reg_N466 ));
AND2_X2 _w_reg_U108  ( .A1(w_d[464]), .A2(_w_reg_n690 ), .ZN(_w_reg_N467 ));
AND2_X2 _w_reg_U107  ( .A1(w_d[465]), .A2(_w_reg_n690 ), .ZN(_w_reg_N468 ));
AND2_X2 _w_reg_U106  ( .A1(w_d[466]), .A2(_w_reg_n690 ), .ZN(_w_reg_N469 ));
AND2_X2 _w_reg_U105  ( .A1(w_d[44]), .A2(_w_reg_n690 ), .ZN(_w_reg_N47 ) );
AND2_X2 _w_reg_U104  ( .A1(w_d[467]), .A2(_w_reg_n690 ), .ZN(_w_reg_N470 ));
AND2_X2 _w_reg_U103  ( .A1(w_d[468]), .A2(_w_reg_n690 ), .ZN(_w_reg_N471 ));
AND2_X2 _w_reg_U102  ( .A1(w_d[469]), .A2(_w_reg_n690 ), .ZN(_w_reg_N472 ));
AND2_X2 _w_reg_U101  ( .A1(w_d[470]), .A2(_w_reg_n680 ), .ZN(_w_reg_N473 ));
AND2_X2 _w_reg_U100  ( .A1(w_d[471]), .A2(_w_reg_n680 ), .ZN(_w_reg_N474 ));
AND2_X2 _w_reg_U99  ( .A1(w_d[472]), .A2(_w_reg_n680 ), .ZN(_w_reg_N475 ) );
AND2_X2 _w_reg_U98  ( .A1(w_d[473]), .A2(_w_reg_n680 ), .ZN(_w_reg_N476 ) );
AND2_X2 _w_reg_U97  ( .A1(w_d[474]), .A2(_w_reg_n680 ), .ZN(_w_reg_N477 ) );
AND2_X2 _w_reg_U96  ( .A1(w_d[475]), .A2(_w_reg_n680 ), .ZN(_w_reg_N478 ) );
AND2_X2 _w_reg_U95  ( .A1(w_d[476]), .A2(_w_reg_n680 ), .ZN(_w_reg_N479 ) );
AND2_X2 _w_reg_U94  ( .A1(w_d[45]), .A2(_w_reg_n680 ), .ZN(_w_reg_N48 ) );
AND2_X2 _w_reg_U93  ( .A1(w_d[477]), .A2(_w_reg_n680 ), .ZN(_w_reg_N480 ) );
AND2_X2 _w_reg_U92  ( .A1(w_d[478]), .A2(_w_reg_n680 ), .ZN(_w_reg_N481 ) );
AND2_X2 _w_reg_U91  ( .A1(w_d[479]), .A2(_w_reg_n680 ), .ZN(_w_reg_N482 ) );
AND2_X2 _w_reg_U83  ( .A1(w_d[46]), .A2(_w_reg_n670 ), .ZN(_w_reg_N49 ) );
AND2_X2 _w_reg_U71  ( .A1(w_d[47]), .A2(_w_reg_n670 ), .ZN(_w_reg_N50 ) );
AND2_X2 _w_reg_U69  ( .A1(w_d[498]), .A2(_w_reg_n670 ), .ZN(_w_reg_N501 ) );
AND2_X2 _w_reg_U68  ( .A1(w_d[499]), .A2(_w_reg_n670 ), .ZN(_w_reg_N502 ) );
AND2_X2 _w_reg_U67  ( .A1(w_d[500]), .A2(_w_reg_n670 ), .ZN(_w_reg_N503 ) );
AND2_X2 _w_reg_U66  ( .A1(w_d[501]), .A2(_w_reg_n670 ), .ZN(_w_reg_N504 ) );
AND2_X2 _w_reg_U65  ( .A1(w_d[502]), .A2(_w_reg_n670 ), .ZN(_w_reg_N505 ) );
AND2_X2 _w_reg_U64  ( .A1(w_d[503]), .A2(_w_reg_n670 ), .ZN(_w_reg_N506 ) );
AND2_X2 _w_reg_U63  ( .A1(w_d[504]), .A2(_w_reg_n670 ), .ZN(_w_reg_N507 ) );
AND2_X2 _w_reg_U62  ( .A1(w_d[505]), .A2(_w_reg_n670 ), .ZN(_w_reg_N508 ) );
AND2_X2 _w_reg_U61  ( .A1(w_d[506]), .A2(_w_reg_n660 ), .ZN(_w_reg_N509 ) );
AND2_X2 _w_reg_U60  ( .A1(w_d[48]), .A2(_w_reg_n660 ), .ZN(_w_reg_N51 ) );
AND2_X2 _w_reg_U59  ( .A1(w_d[507]), .A2(_w_reg_n660 ), .ZN(_w_reg_N510 ) );
AND2_X2 _w_reg_U58  ( .A1(w_d[508]), .A2(_w_reg_n660 ), .ZN(_w_reg_N511 ) );
AND2_X2 _w_reg_U57  ( .A1(w_d[509]), .A2(_w_reg_n660 ), .ZN(_w_reg_N512 ) );
AND2_X2 _w_reg_U56  ( .A1(w_d[510]), .A2(_w_reg_n660 ), .ZN(_w_reg_N513 ) );
AND2_X2 _w_reg_U55  ( .A1(w_d[511]), .A2(_w_reg_n660 ), .ZN(_w_reg_N514 ) );
AND2_X2 _w_reg_U54  ( .A1(w_d[49]), .A2(_w_reg_n660 ), .ZN(_w_reg_N52 ) );
AND2_X2 _w_reg_U53  ( .A1(w_d[50]), .A2(_w_reg_n660 ), .ZN(_w_reg_N53 ) );
AND2_X2 _w_reg_U52  ( .A1(w_d[51]), .A2(_w_reg_n660 ), .ZN(_w_reg_N54 ) );
AND2_X2 _w_reg_U51  ( .A1(w_d[52]), .A2(_w_reg_n660 ), .ZN(_w_reg_N55 ) );
AND2_X2 _w_reg_U50  ( .A1(w_d[53]), .A2(_w_reg_n650 ), .ZN(_w_reg_N56 ) );
AND2_X2 _w_reg_U49  ( .A1(w_d[54]), .A2(_w_reg_n650 ), .ZN(_w_reg_N57 ) );
AND2_X2 _w_reg_U48  ( .A1(w_d[55]), .A2(_w_reg_n650 ), .ZN(_w_reg_N58 ) );
AND2_X2 _w_reg_U47  ( .A1(w_d[56]), .A2(_w_reg_n650 ), .ZN(_w_reg_N59 ) );
AND2_X2 _w_reg_U45  ( .A1(w_d[57]), .A2(_w_reg_n650 ), .ZN(_w_reg_N60 ) );
AND2_X2 _w_reg_U44  ( .A1(w_d[58]), .A2(_w_reg_n650 ), .ZN(_w_reg_N61 ) );
AND2_X2 _w_reg_U43  ( .A1(w_d[59]), .A2(_w_reg_n650 ), .ZN(_w_reg_N62 ) );
AND2_X2 _w_reg_U42  ( .A1(w_d[60]), .A2(_w_reg_n650 ), .ZN(_w_reg_N63 ) );
AND2_X2 _w_reg_U41  ( .A1(w_d[61]), .A2(_w_reg_n650 ), .ZN(_w_reg_N64 ) );
AND2_X2 _w_reg_U40  ( .A1(w_d[62]), .A2(_w_reg_n650 ), .ZN(_w_reg_N65 ) );
AND2_X2 _w_reg_U39  ( .A1(w_d[63]), .A2(_w_reg_n640 ), .ZN(_w_reg_N66 ) );
AND2_X2 _w_reg_U38  ( .A1(w_d[64]), .A2(_w_reg_n640 ), .ZN(_w_reg_N67 ) );
AND2_X2 _w_reg_U37  ( .A1(w_d[65]), .A2(_w_reg_n640 ), .ZN(_w_reg_N68 ) );
AND2_X2 _w_reg_U36  ( .A1(w_d[66]), .A2(_w_reg_n640 ), .ZN(_w_reg_N69 ) );
AND2_X2 _w_reg_U34  ( .A1(w_d[67]), .A2(_w_reg_n640 ), .ZN(_w_reg_N70 ) );
AND2_X2 _w_reg_U33  ( .A1(w_d[68]), .A2(_w_reg_n640 ), .ZN(_w_reg_N71 ) );
AND2_X2 _w_reg_U32  ( .A1(w_d[69]), .A2(_w_reg_n640 ), .ZN(_w_reg_N72 ) );
AND2_X2 _w_reg_U31  ( .A1(w_d[70]), .A2(_w_reg_n640 ), .ZN(_w_reg_N73 ) );
AND2_X2 _w_reg_U30  ( .A1(w_d[71]), .A2(_w_reg_n640 ), .ZN(_w_reg_N74 ) );
AND2_X2 _w_reg_U29  ( .A1(w_d[72]), .A2(_w_reg_n640 ), .ZN(_w_reg_N75 ) );
AND2_X2 _w_reg_U28  ( .A1(w_d[73]), .A2(_w_reg_n630 ), .ZN(_w_reg_N76 ) );
AND2_X2 _w_reg_U27  ( .A1(w_d[74]), .A2(_w_reg_n630 ), .ZN(_w_reg_N77 ) );
AND2_X2 _w_reg_U26  ( .A1(w_d[75]), .A2(_w_reg_n630 ), .ZN(_w_reg_N78 ) );
AND2_X2 _w_reg_U25  ( .A1(w_d[76]), .A2(_w_reg_n630 ), .ZN(_w_reg_N79 ) );
AND2_X2 _w_reg_U23  ( .A1(w_d[77]), .A2(_w_reg_n630 ), .ZN(_w_reg_N80 ) );
AND2_X2 _w_reg_U22  ( .A1(w_d[78]), .A2(_w_reg_n630 ), .ZN(_w_reg_N81 ) );
AND2_X2 _w_reg_U21  ( .A1(w_d[79]), .A2(_w_reg_n630 ), .ZN(_w_reg_N82 ) );
AND2_X2 _w_reg_U20  ( .A1(w_d[80]), .A2(_w_reg_n630 ), .ZN(_w_reg_N83 ) );
AND2_X2 _w_reg_U19  ( .A1(w_d[81]), .A2(_w_reg_n630 ), .ZN(_w_reg_N84 ) );
AND2_X2 _w_reg_U18  ( .A1(w_d[82]), .A2(_w_reg_n630 ), .ZN(_w_reg_N85 ) );
AND2_X2 _w_reg_U17  ( .A1(w_d[83]), .A2(_w_reg_n620 ), .ZN(_w_reg_N86 ) );
AND2_X2 _w_reg_U16  ( .A1(w_d[84]), .A2(_w_reg_n620 ), .ZN(_w_reg_N87 ) );
AND2_X2 _w_reg_U15  ( .A1(w_d[85]), .A2(_w_reg_n620 ), .ZN(_w_reg_N88 ) );
AND2_X2 _w_reg_U14  ( .A1(w_d[86]), .A2(_w_reg_n620 ), .ZN(_w_reg_N89 ) );
AND2_X2 _w_reg_U12  ( .A1(w_d[87]), .A2(_w_reg_n620 ), .ZN(_w_reg_N90 ) );
AND2_X2 _w_reg_U11  ( .A1(w_d[88]), .A2(_w_reg_n620 ), .ZN(_w_reg_N91 ) );
AND2_X2 _w_reg_U10  ( .A1(w_d[89]), .A2(_w_reg_n620 ), .ZN(_w_reg_N92 ) );
AND2_X2 _w_reg_U9  ( .A1(w_d[90]), .A2(_w_reg_n620 ), .ZN(_w_reg_N93 ) );
AND2_X2 _w_reg_U8  ( .A1(w_d[91]), .A2(_w_reg_n620 ), .ZN(_w_reg_N94 ) );
AND2_X2 _w_reg_U7  ( .A1(w_d[92]), .A2(_w_reg_n620 ), .ZN(_w_reg_N95 ) );
AND2_X2 _w_reg_U6  ( .A1(w_d[93]), .A2(_w_reg_n610 ), .ZN(_w_reg_N96 ) );
AND2_X2 _w_reg_U5  ( .A1(w_d[94]), .A2(_w_reg_n610 ), .ZN(_w_reg_N97 ) );
AND2_X2 _w_reg_U4  ( .A1(w_d[95]), .A2(_w_reg_n610 ), .ZN(_w_reg_N98 ) );
AND2_X2 _w_reg_U3  ( .A1(w_d[96]), .A2(_w_reg_n610 ), .ZN(_w_reg_N99 ) );
DFF_X2 _w_reg_q_reg_0_  ( .D(_w_reg_N3 ), .CK(clk), .Q(w_q[0]), .QN() );
DFF_X2 _w_reg_q_reg_1_  ( .D(_w_reg_N4 ), .CK(clk), .Q(w_q[1]), .QN() );
DFF_X2 _w_reg_q_reg_2_  ( .D(_w_reg_N5 ), .CK(clk), .Q(w_q[2]), .QN() );
DFF_X2 _w_reg_q_reg_3_  ( .D(_w_reg_N6 ), .CK(clk), .Q(w_q[3]), .QN() );
DFF_X2 _w_reg_q_reg_4_  ( .D(_w_reg_N7 ), .CK(clk), .Q(w_q[4]), .QN() );
DFF_X2 _w_reg_q_reg_5_  ( .D(_w_reg_N8 ), .CK(clk), .Q(w_q[5]), .QN() );
DFF_X2 _w_reg_q_reg_6_  ( .D(_w_reg_N9 ), .CK(clk), .Q(w_q[6]), .QN() );
DFF_X2 _w_reg_q_reg_7_  ( .D(_w_reg_N10 ), .CK(clk), .Q(w_q[7]), .QN() );
DFF_X2 _w_reg_q_reg_8_  ( .D(_w_reg_N11 ), .CK(clk), .Q(w_q[8]), .QN() );
DFF_X2 _w_reg_q_reg_9_  ( .D(_w_reg_N12 ), .CK(clk), .Q(w_q[9]), .QN() );
DFF_X2 _w_reg_q_reg_10_  ( .D(_w_reg_N13 ), .CK(clk), .Q(w_q[10]), .QN() );
DFF_X2 _w_reg_q_reg_11_  ( .D(_w_reg_N14 ), .CK(clk), .Q(w_q[11]), .QN() );
DFF_X2 _w_reg_q_reg_12_  ( .D(_w_reg_N15 ), .CK(clk), .Q(w_q[12]), .QN() );
DFF_X2 _w_reg_q_reg_13_  ( .D(_w_reg_N16 ), .CK(clk), .Q(w_q[13]), .QN() );
DFF_X2 _w_reg_q_reg_14_  ( .D(_w_reg_N17 ), .CK(clk), .Q(w_q[14]), .QN() );
DFF_X2 _w_reg_q_reg_15_  ( .D(_w_reg_N18 ), .CK(clk), .Q(w_q[15]), .QN() );
DFF_X2 _w_reg_q_reg_16_  ( .D(_w_reg_N19 ), .CK(clk), .Q(w_q[16]), .QN() );
DFF_X2 _w_reg_q_reg_17_  ( .D(_w_reg_N20 ), .CK(clk), .Q(w_q[17]), .QN() );
DFF_X2 _w_reg_q_reg_18_  ( .D(_w_reg_N21 ), .CK(clk), .Q(w_q[18]), .QN() );
DFF_X2 _w_reg_q_reg_19_  ( .D(_w_reg_N22 ), .CK(clk), .Q(w_q[19]), .QN() );
DFF_X2 _w_reg_q_reg_20_  ( .D(_w_reg_N23 ), .CK(clk), .Q(w_q[20]), .QN() );
DFF_X2 _w_reg_q_reg_21_  ( .D(_w_reg_N24 ), .CK(clk), .Q(w_q[21]), .QN() );
DFF_X2 _w_reg_q_reg_22_  ( .D(_w_reg_N25 ), .CK(clk), .Q(w_q[22]), .QN() );
DFF_X2 _w_reg_q_reg_23_  ( .D(_w_reg_N26 ), .CK(clk), .Q(w_q[23]), .QN() );
DFF_X2 _w_reg_q_reg_24_  ( .D(_w_reg_N27 ), .CK(clk), .Q(w_q[24]), .QN() );
DFF_X2 _w_reg_q_reg_25_  ( .D(_w_reg_N28 ), .CK(clk), .Q(w_q[25]), .QN() );
DFF_X2 _w_reg_q_reg_26_  ( .D(_w_reg_N29 ), .CK(clk), .Q(w_q[26]), .QN() );
DFF_X2 _w_reg_q_reg_27_  ( .D(_w_reg_N30 ), .CK(clk), .Q(w_q[27]), .QN() );
DFF_X2 _w_reg_q_reg_28_  ( .D(_w_reg_N31 ), .CK(clk), .Q(w_q[28]), .QN() );
DFF_X2 _w_reg_q_reg_29_  ( .D(_w_reg_N32 ), .CK(clk), .Q(w_q[29]), .QN() );
DFF_X2 _w_reg_q_reg_30_  ( .D(_w_reg_N33 ), .CK(clk), .Q(w_q[30]), .QN() );
DFF_X2 _w_reg_q_reg_31_  ( .D(_w_reg_N34 ), .CK(clk), .Q(w_q[31]), .QN() );
DFF_X2 _w_reg_q_reg_32_  ( .D(_w_reg_N35 ), .CK(clk), .Q(w_q[32]), .QN() );
DFF_X2 _w_reg_q_reg_33_  ( .D(_w_reg_N36 ), .CK(clk), .Q(w_q[33]), .QN() );
DFF_X2 _w_reg_q_reg_34_  ( .D(_w_reg_N37 ), .CK(clk), .Q(w_q[34]), .QN() );
DFF_X2 _w_reg_q_reg_35_  ( .D(_w_reg_N38 ), .CK(clk), .Q(w_q[35]), .QN() );
DFF_X2 _w_reg_q_reg_36_  ( .D(_w_reg_N39 ), .CK(clk), .Q(w_q[36]), .QN() );
DFF_X2 _w_reg_q_reg_37_  ( .D(_w_reg_N40 ), .CK(clk), .Q(w_q[37]), .QN() );
DFF_X2 _w_reg_q_reg_38_  ( .D(_w_reg_N41 ), .CK(clk), .Q(w_q[38]), .QN() );
DFF_X2 _w_reg_q_reg_39_  ( .D(_w_reg_N42 ), .CK(clk), .Q(w_q[39]), .QN() );
DFF_X2 _w_reg_q_reg_40_  ( .D(_w_reg_N43 ), .CK(clk), .Q(w_q[40]), .QN() );
DFF_X2 _w_reg_q_reg_41_  ( .D(_w_reg_N44 ), .CK(clk), .Q(w_q[41]), .QN() );
DFF_X2 _w_reg_q_reg_42_  ( .D(_w_reg_N45 ), .CK(clk), .Q(w_q[42]), .QN() );
DFF_X2 _w_reg_q_reg_43_  ( .D(_w_reg_N46 ), .CK(clk), .Q(w_q[43]), .QN() );
DFF_X2 _w_reg_q_reg_44_  ( .D(_w_reg_N47 ), .CK(clk), .Q(w_q[44]), .QN() );
DFF_X2 _w_reg_q_reg_45_  ( .D(_w_reg_N48 ), .CK(clk), .Q(w_q[45]), .QN() );
DFF_X2 _w_reg_q_reg_46_  ( .D(_w_reg_N49 ), .CK(clk), .Q(w_q[46]), .QN() );
DFF_X2 _w_reg_q_reg_47_  ( .D(_w_reg_N50 ), .CK(clk), .Q(w_q[47]), .QN() );
DFF_X2 _w_reg_q_reg_48_  ( .D(_w_reg_N51 ), .CK(clk), .Q(w_q[48]), .QN() );
DFF_X2 _w_reg_q_reg_49_  ( .D(_w_reg_N52 ), .CK(clk), .Q(w_q[49]), .QN() );
DFF_X2 _w_reg_q_reg_50_  ( .D(_w_reg_N53 ), .CK(clk), .Q(w_q[50]), .QN() );
DFF_X2 _w_reg_q_reg_51_  ( .D(_w_reg_N54 ), .CK(clk), .Q(w_q[51]), .QN() );
DFF_X2 _w_reg_q_reg_52_  ( .D(_w_reg_N55 ), .CK(clk), .Q(w_q[52]), .QN() );
DFF_X2 _w_reg_q_reg_53_  ( .D(_w_reg_N56 ), .CK(clk), .Q(w_q[53]), .QN() );
DFF_X2 _w_reg_q_reg_54_  ( .D(_w_reg_N57 ), .CK(clk), .Q(w_q[54]), .QN() );
DFF_X2 _w_reg_q_reg_55_  ( .D(_w_reg_N58 ), .CK(clk), .Q(w_q[55]), .QN() );
DFF_X2 _w_reg_q_reg_56_  ( .D(_w_reg_N59 ), .CK(clk), .Q(w_q[56]), .QN() );
DFF_X2 _w_reg_q_reg_57_  ( .D(_w_reg_N60 ), .CK(clk), .Q(w_q[57]), .QN() );
DFF_X2 _w_reg_q_reg_58_  ( .D(_w_reg_N61 ), .CK(clk), .Q(w_q[58]), .QN() );
DFF_X2 _w_reg_q_reg_59_  ( .D(_w_reg_N62 ), .CK(clk), .Q(w_q[59]), .QN() );
DFF_X2 _w_reg_q_reg_60_  ( .D(_w_reg_N63 ), .CK(clk), .Q(w_q[60]), .QN() );
DFF_X2 _w_reg_q_reg_61_  ( .D(_w_reg_N64 ), .CK(clk), .Q(w_q[61]), .QN() );
DFF_X2 _w_reg_q_reg_62_  ( .D(_w_reg_N65 ), .CK(clk), .Q(w_q[62]), .QN() );
DFF_X2 _w_reg_q_reg_63_  ( .D(_w_reg_N66 ), .CK(clk), .Q(w_q[63]), .QN() );
DFF_X2 _w_reg_q_reg_64_  ( .D(_w_reg_N67 ), .CK(clk), .Q(w_q[64]), .QN() );
DFF_X2 _w_reg_q_reg_65_  ( .D(_w_reg_N68 ), .CK(clk), .Q(w_q[65]), .QN() );
DFF_X2 _w_reg_q_reg_66_  ( .D(_w_reg_N69 ), .CK(clk), .Q(w_q[66]), .QN() );
DFF_X2 _w_reg_q_reg_67_  ( .D(_w_reg_N70 ), .CK(clk), .Q(w_q[67]), .QN() );
DFF_X2 _w_reg_q_reg_68_  ( .D(_w_reg_N71 ), .CK(clk), .Q(w_q[68]), .QN() );
DFF_X2 _w_reg_q_reg_69_  ( .D(_w_reg_N72 ), .CK(clk), .Q(w_q[69]), .QN() );
DFF_X2 _w_reg_q_reg_70_  ( .D(_w_reg_N73 ), .CK(clk), .Q(w_q[70]), .QN() );
DFF_X2 _w_reg_q_reg_71_  ( .D(_w_reg_N74 ), .CK(clk), .Q(w_q[71]), .QN() );
DFF_X2 _w_reg_q_reg_72_  ( .D(_w_reg_N75 ), .CK(clk), .Q(w_q[72]), .QN() );
DFF_X2 _w_reg_q_reg_73_  ( .D(_w_reg_N76 ), .CK(clk), .Q(w_q[73]), .QN() );
DFF_X2 _w_reg_q_reg_74_  ( .D(_w_reg_N77 ), .CK(clk), .Q(w_q[74]), .QN() );
DFF_X2 _w_reg_q_reg_75_  ( .D(_w_reg_N78 ), .CK(clk), .Q(w_q[75]), .QN() );
DFF_X2 _w_reg_q_reg_76_  ( .D(_w_reg_N79 ), .CK(clk), .Q(w_q[76]), .QN() );
DFF_X2 _w_reg_q_reg_77_  ( .D(_w_reg_N80 ), .CK(clk), .Q(w_q[77]), .QN() );
DFF_X2 _w_reg_q_reg_78_  ( .D(_w_reg_N81 ), .CK(clk), .Q(w_q[78]), .QN() );
DFF_X2 _w_reg_q_reg_79_  ( .D(_w_reg_N82 ), .CK(clk), .Q(w_q[79]), .QN() );
DFF_X2 _w_reg_q_reg_80_  ( .D(_w_reg_N83 ), .CK(clk), .Q(w_q[80]), .QN() );
DFF_X2 _w_reg_q_reg_81_  ( .D(_w_reg_N84 ), .CK(clk), .Q(w_q[81]), .QN() );
DFF_X2 _w_reg_q_reg_82_  ( .D(_w_reg_N85 ), .CK(clk), .Q(w_q[82]), .QN() );
DFF_X2 _w_reg_q_reg_83_  ( .D(_w_reg_N86 ), .CK(clk), .Q(w_q[83]), .QN() );
DFF_X2 _w_reg_q_reg_84_  ( .D(_w_reg_N87 ), .CK(clk), .Q(w_q[84]), .QN() );
DFF_X2 _w_reg_q_reg_85_  ( .D(_w_reg_N88 ), .CK(clk), .Q(w_q[85]), .QN() );
DFF_X2 _w_reg_q_reg_86_  ( .D(_w_reg_N89 ), .CK(clk), .Q(w_q[86]), .QN() );
DFF_X2 _w_reg_q_reg_87_  ( .D(_w_reg_N90 ), .CK(clk), .Q(w_q[87]), .QN() );
DFF_X2 _w_reg_q_reg_88_  ( .D(_w_reg_N91 ), .CK(clk), .Q(w_q[88]), .QN() );
DFF_X2 _w_reg_q_reg_89_  ( .D(_w_reg_N92 ), .CK(clk), .Q(w_q[89]), .QN() );
DFF_X2 _w_reg_q_reg_90_  ( .D(_w_reg_N93 ), .CK(clk), .Q(w_q[90]), .QN() );
DFF_X2 _w_reg_q_reg_91_  ( .D(_w_reg_N94 ), .CK(clk), .Q(w_q[91]), .QN() );
DFF_X2 _w_reg_q_reg_92_  ( .D(_w_reg_N95 ), .CK(clk), .Q(w_q[92]), .QN() );
DFF_X2 _w_reg_q_reg_93_  ( .D(_w_reg_N96 ), .CK(clk), .Q(w_q[93]), .QN() );
DFF_X2 _w_reg_q_reg_94_  ( .D(_w_reg_N97 ), .CK(clk), .Q(w_q[94]), .QN() );
DFF_X2 _w_reg_q_reg_95_  ( .D(_w_reg_N98 ), .CK(clk), .Q(w_q[95]), .QN() );
DFF_X2 _w_reg_q_reg_96_  ( .D(_w_reg_N99 ), .CK(clk), .Q(w_q[96]), .QN() );
DFF_X2 _w_reg_q_reg_97_  ( .D(_w_reg_N100 ), .CK(clk), .Q(w_q[97]), .QN() );
DFF_X2 _w_reg_q_reg_98_  ( .D(_w_reg_N101 ), .CK(clk), .Q(w_q[98]), .QN() );
DFF_X2 _w_reg_q_reg_99_  ( .D(_w_reg_N102 ), .CK(clk), .Q(w_q[99]), .QN() );
DFF_X2 _w_reg_q_reg_100_  ( .D(_w_reg_N103 ), .CK(clk), .Q(w_q[100]), .QN());
DFF_X2 _w_reg_q_reg_101_  ( .D(_w_reg_N104 ), .CK(clk), .Q(w_q[101]), .QN());
DFF_X2 _w_reg_q_reg_102_  ( .D(_w_reg_N105 ), .CK(clk), .Q(w_q[102]), .QN());
DFF_X2 _w_reg_q_reg_103_  ( .D(_w_reg_N106 ), .CK(clk), .Q(w_q[103]), .QN());
DFF_X2 _w_reg_q_reg_104_  ( .D(_w_reg_N107 ), .CK(clk), .Q(w_q[104]), .QN());
DFF_X2 _w_reg_q_reg_105_  ( .D(_w_reg_N108 ), .CK(clk), .Q(w_q[105]), .QN());
DFF_X2 _w_reg_q_reg_106_  ( .D(_w_reg_N109 ), .CK(clk), .Q(w_q[106]), .QN());
DFF_X2 _w_reg_q_reg_107_  ( .D(_w_reg_N110 ), .CK(clk), .Q(w_q[107]), .QN());
DFF_X2 _w_reg_q_reg_108_  ( .D(_w_reg_N111 ), .CK(clk), .Q(w_q[108]), .QN());
DFF_X2 _w_reg_q_reg_109_  ( .D(_w_reg_N112 ), .CK(clk), .Q(w_q[109]), .QN());
DFF_X2 _w_reg_q_reg_110_  ( .D(_w_reg_N113 ), .CK(clk), .Q(w_q[110]), .QN());
DFF_X2 _w_reg_q_reg_111_  ( .D(_w_reg_N114 ), .CK(clk), .Q(w_q[111]), .QN());
DFF_X2 _w_reg_q_reg_112_  ( .D(_w_reg_N115 ), .CK(clk), .Q(w_q[112]), .QN());
DFF_X2 _w_reg_q_reg_113_  ( .D(_w_reg_N116 ), .CK(clk), .Q(w_q[113]), .QN());
DFF_X2 _w_reg_q_reg_114_  ( .D(_w_reg_N117 ), .CK(clk), .Q(w_q[114]), .QN());
DFF_X2 _w_reg_q_reg_115_  ( .D(_w_reg_N118 ), .CK(clk), .Q(w_q[115]), .QN());
DFF_X2 _w_reg_q_reg_116_  ( .D(_w_reg_N119 ), .CK(clk), .Q(w_q[116]), .QN());
DFF_X2 _w_reg_q_reg_117_  ( .D(_w_reg_N120 ), .CK(clk), .Q(w_q[117]), .QN());
DFF_X2 _w_reg_q_reg_118_  ( .D(_w_reg_N121 ), .CK(clk), .Q(w_q[118]), .QN());
DFF_X2 _w_reg_q_reg_119_  ( .D(_w_reg_N122 ), .CK(clk), .Q(w_q[119]), .QN());
DFF_X2 _w_reg_q_reg_120_  ( .D(_w_reg_N123 ), .CK(clk), .Q(w_q[120]), .QN());
DFF_X2 _w_reg_q_reg_121_  ( .D(_w_reg_N124 ), .CK(clk), .Q(w_q[121]), .QN());
DFF_X2 _w_reg_q_reg_122_  ( .D(_w_reg_N125 ), .CK(clk), .Q(w_q[122]), .QN());
DFF_X2 _w_reg_q_reg_123_  ( .D(_w_reg_N126 ), .CK(clk), .Q(w_q[123]), .QN());
DFF_X2 _w_reg_q_reg_124_  ( .D(_w_reg_N127 ), .CK(clk), .Q(w_q[124]), .QN());
DFF_X2 _w_reg_q_reg_125_  ( .D(_w_reg_N128 ), .CK(clk), .Q(w_q[125]), .QN());
DFF_X2 _w_reg_q_reg_126_  ( .D(_w_reg_N129 ), .CK(clk), .Q(w_q[126]), .QN());
DFF_X2 _w_reg_q_reg_127_  ( .D(_w_reg_N130 ), .CK(clk), .Q(w_q[127]), .QN());
DFF_X2 _w_reg_q_reg_128_  ( .D(_w_reg_N131 ), .CK(clk), .Q(w_q[128]), .QN());
DFF_X2 _w_reg_q_reg_129_  ( .D(_w_reg_N132 ), .CK(clk), .Q(w_q[129]), .QN());
DFF_X2 _w_reg_q_reg_130_  ( .D(_w_reg_N133 ), .CK(clk), .Q(w_q[130]), .QN());
DFF_X2 _w_reg_q_reg_131_  ( .D(_w_reg_N134 ), .CK(clk), .Q(w_q[131]), .QN());
DFF_X2 _w_reg_q_reg_132_  ( .D(_w_reg_N135 ), .CK(clk), .Q(w_q[132]), .QN());
DFF_X2 _w_reg_q_reg_133_  ( .D(_w_reg_N136 ), .CK(clk), .Q(w_q[133]), .QN());
DFF_X2 _w_reg_q_reg_134_  ( .D(_w_reg_N137 ), .CK(clk), .Q(w_q[134]), .QN());
DFF_X2 _w_reg_q_reg_135_  ( .D(_w_reg_N138 ), .CK(clk), .Q(w_q[135]), .QN());
DFF_X2 _w_reg_q_reg_136_  ( .D(_w_reg_N139 ), .CK(clk), .Q(w_q[136]), .QN());
DFF_X2 _w_reg_q_reg_137_  ( .D(_w_reg_N140 ), .CK(clk), .Q(w_q[137]), .QN());
DFF_X2 _w_reg_q_reg_138_  ( .D(_w_reg_N141 ), .CK(clk), .Q(w_q[138]), .QN());
DFF_X2 _w_reg_q_reg_139_  ( .D(_w_reg_N142 ), .CK(clk), .Q(w_q[139]), .QN());
DFF_X2 _w_reg_q_reg_140_  ( .D(_w_reg_N143 ), .CK(clk), .Q(w_q[140]), .QN());
DFF_X2 _w_reg_q_reg_141_  ( .D(_w_reg_N144 ), .CK(clk), .Q(w_q[141]), .QN());
DFF_X2 _w_reg_q_reg_142_  ( .D(_w_reg_N145 ), .CK(clk), .Q(w_q[142]), .QN());
DFF_X2 _w_reg_q_reg_143_  ( .D(_w_reg_N146 ), .CK(clk), .Q(w_q[143]), .QN());
DFF_X2 _w_reg_q_reg_144_  ( .D(_w_reg_N147 ), .CK(clk), .Q(w_q[144]), .QN());
DFF_X2 _w_reg_q_reg_145_  ( .D(_w_reg_N148 ), .CK(clk), .Q(w_q[145]), .QN());
DFF_X2 _w_reg_q_reg_146_  ( .D(_w_reg_N149 ), .CK(clk), .Q(w_q[146]), .QN());
DFF_X2 _w_reg_q_reg_147_  ( .D(_w_reg_N150 ), .CK(clk), .Q(w_q[147]), .QN());
DFF_X2 _w_reg_q_reg_148_  ( .D(_w_reg_N151 ), .CK(clk), .Q(w_q[148]), .QN());
DFF_X2 _w_reg_q_reg_149_  ( .D(_w_reg_N152 ), .CK(clk), .Q(w_q[149]), .QN());
DFF_X2 _w_reg_q_reg_150_  ( .D(_w_reg_N153 ), .CK(clk), .Q(w_q[150]), .QN());
DFF_X2 _w_reg_q_reg_151_  ( .D(_w_reg_N154 ), .CK(clk), .Q(w_q[151]), .QN());
DFF_X2 _w_reg_q_reg_152_  ( .D(_w_reg_N155 ), .CK(clk), .Q(w_q[152]), .QN());
DFF_X2 _w_reg_q_reg_153_  ( .D(_w_reg_N156 ), .CK(clk), .Q(w_q[153]), .QN());
DFF_X2 _w_reg_q_reg_154_  ( .D(_w_reg_N157 ), .CK(clk), .Q(w_q[154]), .QN());
DFF_X2 _w_reg_q_reg_155_  ( .D(_w_reg_N158 ), .CK(clk), .Q(w_q[155]), .QN());
DFF_X2 _w_reg_q_reg_156_  ( .D(_w_reg_N159 ), .CK(clk), .Q(w_q[156]), .QN());
DFF_X2 _w_reg_q_reg_157_  ( .D(_w_reg_N160 ), .CK(clk), .Q(w_q[157]), .QN());
DFF_X2 _w_reg_q_reg_158_  ( .D(_w_reg_N161 ), .CK(clk), .Q(w_q[158]), .QN());
DFF_X2 _w_reg_q_reg_159_  ( .D(_w_reg_N162 ), .CK(clk), .Q(w_q[159]), .QN());
DFF_X2 _w_reg_q_reg_160_  ( .D(_w_reg_N163 ), .CK(clk), .Q(w_q[160]), .QN());
DFF_X2 _w_reg_q_reg_161_  ( .D(_w_reg_N164 ), .CK(clk), .Q(w_q[161]), .QN());
DFF_X2 _w_reg_q_reg_162_  ( .D(_w_reg_N165 ), .CK(clk), .Q(w_q[162]), .QN());
DFF_X2 _w_reg_q_reg_163_  ( .D(_w_reg_N166 ), .CK(clk), .Q(w_q[163]), .QN());
DFF_X2 _w_reg_q_reg_164_  ( .D(_w_reg_N167 ), .CK(clk), .Q(w_q[164]), .QN());
DFF_X2 _w_reg_q_reg_165_  ( .D(_w_reg_N168 ), .CK(clk), .Q(w_q[165]), .QN());
DFF_X2 _w_reg_q_reg_166_  ( .D(_w_reg_N169 ), .CK(clk), .Q(w_q[166]), .QN());
DFF_X2 _w_reg_q_reg_167_  ( .D(_w_reg_N170 ), .CK(clk), .Q(w_q[167]), .QN());
DFF_X2 _w_reg_q_reg_168_  ( .D(_w_reg_N171 ), .CK(clk), .Q(w_q[168]), .QN());
DFF_X2 _w_reg_q_reg_169_  ( .D(_w_reg_N172 ), .CK(clk), .Q(w_q[169]), .QN());
DFF_X2 _w_reg_q_reg_170_  ( .D(_w_reg_N173 ), .CK(clk), .Q(w_q[170]), .QN());
DFF_X2 _w_reg_q_reg_171_  ( .D(_w_reg_N174 ), .CK(clk), .Q(w_q[171]), .QN());
DFF_X2 _w_reg_q_reg_172_  ( .D(_w_reg_N175 ), .CK(clk), .Q(w_q[172]), .QN());
DFF_X2 _w_reg_q_reg_173_  ( .D(_w_reg_N176 ), .CK(clk), .Q(w_q[173]), .QN());
DFF_X2 _w_reg_q_reg_174_  ( .D(_w_reg_N177 ), .CK(clk), .Q(w_q[174]), .QN());
DFF_X2 _w_reg_q_reg_175_  ( .D(_w_reg_N178 ), .CK(clk), .Q(w_q[175]), .QN());
DFF_X2 _w_reg_q_reg_176_  ( .D(_w_reg_N179 ), .CK(clk), .Q(w_q[176]), .QN());
DFF_X2 _w_reg_q_reg_177_  ( .D(_w_reg_N180 ), .CK(clk), .Q(w_q[177]), .QN());
DFF_X2 _w_reg_q_reg_178_  ( .D(_w_reg_N181 ), .CK(clk), .Q(w_q[178]), .QN());
DFF_X2 _w_reg_q_reg_179_  ( .D(_w_reg_N182 ), .CK(clk), .Q(w_q[179]), .QN());
DFF_X2 _w_reg_q_reg_180_  ( .D(_w_reg_N183 ), .CK(clk), .Q(w_q[180]), .QN());
DFF_X2 _w_reg_q_reg_181_  ( .D(_w_reg_N184 ), .CK(clk), .Q(w_q[181]), .QN());
DFF_X2 _w_reg_q_reg_182_  ( .D(_w_reg_N185 ), .CK(clk), .Q(w_q[182]), .QN());
DFF_X2 _w_reg_q_reg_183_  ( .D(_w_reg_N186 ), .CK(clk), .Q(w_q[183]), .QN());
DFF_X2 _w_reg_q_reg_184_  ( .D(_w_reg_N187 ), .CK(clk), .Q(w_q[184]), .QN());
DFF_X2 _w_reg_q_reg_185_  ( .D(_w_reg_N188 ), .CK(clk), .Q(w_q[185]), .QN());
DFF_X2 _w_reg_q_reg_186_  ( .D(_w_reg_N189 ), .CK(clk), .Q(w_q[186]), .QN());
DFF_X2 _w_reg_q_reg_187_  ( .D(_w_reg_N190 ), .CK(clk), .Q(w_q[187]), .QN());
DFF_X2 _w_reg_q_reg_188_  ( .D(_w_reg_N191 ), .CK(clk), .Q(w_q[188]), .QN());
DFF_X2 _w_reg_q_reg_189_  ( .D(_w_reg_N192 ), .CK(clk), .Q(w_q[189]), .QN());
DFF_X2 _w_reg_q_reg_190_  ( .D(_w_reg_N193 ), .CK(clk), .Q(w_q[190]), .QN());
DFF_X2 _w_reg_q_reg_191_  ( .D(_w_reg_N194 ), .CK(clk), .Q(w_q[191]), .QN());
DFF_X2 _w_reg_q_reg_192_  ( .D(_w_reg_N195 ), .CK(clk), .Q(w_q[192]), .QN());
DFF_X2 _w_reg_q_reg_193_  ( .D(_w_reg_N196 ), .CK(clk), .Q(w_q[193]), .QN());
DFF_X2 _w_reg_q_reg_194_  ( .D(_w_reg_N197 ), .CK(clk), .Q(w_q[194]), .QN());
DFF_X2 _w_reg_q_reg_195_  ( .D(_w_reg_N198 ), .CK(clk), .Q(w_q[195]), .QN());
DFF_X2 _w_reg_q_reg_196_  ( .D(_w_reg_N199 ), .CK(clk), .Q(w_q[196]), .QN());
DFF_X2 _w_reg_q_reg_197_  ( .D(_w_reg_N200 ), .CK(clk), .Q(w_q[197]), .QN());
DFF_X2 _w_reg_q_reg_198_  ( .D(_w_reg_N201 ), .CK(clk), .Q(w_q[198]), .QN());
DFF_X2 _w_reg_q_reg_199_  ( .D(_w_reg_N202 ), .CK(clk), .Q(w_q[199]), .QN());
DFF_X2 _w_reg_q_reg_200_  ( .D(_w_reg_N203 ), .CK(clk), .Q(w_q[200]), .QN());
DFF_X2 _w_reg_q_reg_201_  ( .D(_w_reg_N204 ), .CK(clk), .Q(w_q[201]), .QN());
DFF_X2 _w_reg_q_reg_202_  ( .D(_w_reg_N205 ), .CK(clk), .Q(w_q[202]), .QN());
DFF_X2 _w_reg_q_reg_203_  ( .D(_w_reg_N206 ), .CK(clk), .Q(w_q[203]), .QN());
DFF_X2 _w_reg_q_reg_204_  ( .D(_w_reg_N207 ), .CK(clk), .Q(w_q[204]), .QN());
DFF_X2 _w_reg_q_reg_205_  ( .D(_w_reg_N208 ), .CK(clk), .Q(w_q[205]), .QN());
DFF_X2 _w_reg_q_reg_206_  ( .D(_w_reg_N209 ), .CK(clk), .Q(w_q[206]), .QN());
DFF_X2 _w_reg_q_reg_207_  ( .D(_w_reg_N210 ), .CK(clk), .Q(w_q[207]), .QN());
DFF_X2 _w_reg_q_reg_208_  ( .D(_w_reg_N211 ), .CK(clk), .Q(w_q[208]), .QN());
DFF_X2 _w_reg_q_reg_209_  ( .D(_w_reg_N212 ), .CK(clk), .Q(w_q[209]), .QN());
DFF_X2 _w_reg_q_reg_210_  ( .D(_w_reg_N213 ), .CK(clk), .Q(w_q[210]), .QN());
DFF_X2 _w_reg_q_reg_211_  ( .D(_w_reg_N214 ), .CK(clk), .Q(w_q[211]), .QN());
DFF_X2 _w_reg_q_reg_212_  ( .D(_w_reg_N215 ), .CK(clk), .Q(w_q[212]), .QN());
DFF_X2 _w_reg_q_reg_213_  ( .D(_w_reg_N216 ), .CK(clk), .Q(w_q[213]), .QN());
DFF_X2 _w_reg_q_reg_214_  ( .D(_w_reg_N217 ), .CK(clk), .Q(w_q[214]), .QN());
DFF_X2 _w_reg_q_reg_215_  ( .D(_w_reg_N218 ), .CK(clk), .Q(w_q[215]), .QN());
DFF_X2 _w_reg_q_reg_216_  ( .D(_w_reg_N219 ), .CK(clk), .Q(w_q[216]), .QN());
DFF_X2 _w_reg_q_reg_217_  ( .D(_w_reg_N220 ), .CK(clk), .Q(w_q[217]), .QN());
DFF_X2 _w_reg_q_reg_218_  ( .D(_w_reg_N221 ), .CK(clk), .Q(w_q[218]), .QN());
DFF_X2 _w_reg_q_reg_219_  ( .D(_w_reg_N222 ), .CK(clk), .Q(w_q[219]), .QN());
DFF_X2 _w_reg_q_reg_220_  ( .D(_w_reg_N223 ), .CK(clk), .Q(w_q[220]), .QN());
DFF_X2 _w_reg_q_reg_221_  ( .D(_w_reg_N224 ), .CK(clk), .Q(w_q[221]), .QN());
DFF_X2 _w_reg_q_reg_222_  ( .D(_w_reg_N225 ), .CK(clk), .Q(w_q[222]), .QN());
DFF_X2 _w_reg_q_reg_223_  ( .D(_w_reg_N226 ), .CK(clk), .Q(w_q[223]), .QN());
DFF_X2 _w_reg_q_reg_224_  ( .D(_w_reg_N227 ), .CK(clk), .Q(w_q[224]), .QN());
DFF_X2 _w_reg_q_reg_225_  ( .D(_w_reg_N228 ), .CK(clk), .Q(w_q[225]), .QN());
DFF_X2 _w_reg_q_reg_226_  ( .D(_w_reg_N229 ), .CK(clk), .Q(w_q[226]), .QN());
DFF_X2 _w_reg_q_reg_227_  ( .D(_w_reg_N230 ), .CK(clk), .Q(w_q[227]), .QN());
DFF_X2 _w_reg_q_reg_228_  ( .D(_w_reg_N231 ), .CK(clk), .Q(w_q[228]), .QN());
DFF_X2 _w_reg_q_reg_229_  ( .D(_w_reg_N232 ), .CK(clk), .Q(w_q[229]), .QN());
DFF_X2 _w_reg_q_reg_230_  ( .D(_w_reg_N233 ), .CK(clk), .Q(w_q[230]), .QN());
DFF_X2 _w_reg_q_reg_231_  ( .D(_w_reg_N234 ), .CK(clk), .Q(w_q[231]), .QN());
DFF_X2 _w_reg_q_reg_232_  ( .D(_w_reg_N235 ), .CK(clk), .Q(w_q[232]), .QN());
DFF_X2 _w_reg_q_reg_233_  ( .D(_w_reg_N236 ), .CK(clk), .Q(w_q[233]), .QN());
DFF_X2 _w_reg_q_reg_234_  ( .D(_w_reg_N237 ), .CK(clk), .Q(w_q[234]), .QN());
DFF_X2 _w_reg_q_reg_235_  ( .D(_w_reg_N238 ), .CK(clk), .Q(w_q[235]), .QN());
DFF_X2 _w_reg_q_reg_236_  ( .D(_w_reg_N239 ), .CK(clk), .Q(w_q[236]), .QN());
DFF_X2 _w_reg_q_reg_237_  ( .D(_w_reg_N240 ), .CK(clk), .Q(w_q[237]), .QN());
DFF_X2 _w_reg_q_reg_238_  ( .D(_w_reg_N241 ), .CK(clk), .Q(w_q[238]), .QN());
DFF_X2 _w_reg_q_reg_239_  ( .D(_w_reg_N242 ), .CK(clk), .Q(w_q[239]), .QN());
DFF_X2 _w_reg_q_reg_240_  ( .D(_w_reg_N243 ), .CK(clk), .Q(w_q[240]), .QN());
DFF_X2 _w_reg_q_reg_241_  ( .D(_w_reg_N244 ), .CK(clk), .Q(w_q[241]), .QN());
DFF_X2 _w_reg_q_reg_242_  ( .D(_w_reg_N245 ), .CK(clk), .Q(w_q[242]), .QN());
DFF_X2 _w_reg_q_reg_243_  ( .D(_w_reg_N246 ), .CK(clk), .Q(w_q[243]), .QN());
DFF_X2 _w_reg_q_reg_244_  ( .D(_w_reg_N247 ), .CK(clk), .Q(w_q[244]), .QN());
DFF_X2 _w_reg_q_reg_245_  ( .D(_w_reg_N248 ), .CK(clk), .Q(w_q[245]), .QN());
DFF_X2 _w_reg_q_reg_246_  ( .D(_w_reg_N249 ), .CK(clk), .Q(w_q[246]), .QN());
DFF_X2 _w_reg_q_reg_247_  ( .D(_w_reg_N250 ), .CK(clk), .Q(w_q[247]), .QN());
DFF_X2 _w_reg_q_reg_248_  ( .D(_w_reg_N251 ), .CK(clk), .Q(w_q[248]), .QN());
DFF_X2 _w_reg_q_reg_249_  ( .D(_w_reg_N252 ), .CK(clk), .Q(w_q[249]), .QN());
DFF_X2 _w_reg_q_reg_250_  ( .D(_w_reg_N253 ), .CK(clk), .Q(w_q[250]), .QN());
DFF_X2 _w_reg_q_reg_251_  ( .D(_w_reg_N254 ), .CK(clk), .Q(w_q[251]), .QN());
DFF_X2 _w_reg_q_reg_252_  ( .D(_w_reg_N255 ), .CK(clk), .Q(w_q[252]), .QN());
DFF_X2 _w_reg_q_reg_253_  ( .D(_w_reg_N256 ), .CK(clk), .Q(w_q[253]), .QN());
DFF_X2 _w_reg_q_reg_254_  ( .D(_w_reg_N257 ), .CK(clk), .Q(w_q[254]), .QN());
DFF_X2 _w_reg_q_reg_255_  ( .D(_w_reg_N258 ), .CK(clk), .Q(w_q[255]), .QN());
DFF_X2 _w_reg_q_reg_256_  ( .D(_w_reg_N259 ), .CK(clk), .Q(w_q[256]), .QN());
DFF_X2 _w_reg_q_reg_257_  ( .D(_w_reg_N260 ), .CK(clk), .Q(w_q[257]), .QN());
DFF_X2 _w_reg_q_reg_258_  ( .D(_w_reg_N261 ), .CK(clk), .Q(w_q[258]), .QN());
DFF_X2 _w_reg_q_reg_259_  ( .D(_w_reg_N262 ), .CK(clk), .Q(w_q[259]), .QN());
DFF_X2 _w_reg_q_reg_260_  ( .D(_w_reg_N263 ), .CK(clk), .Q(w_q[260]), .QN());
DFF_X2 _w_reg_q_reg_261_  ( .D(_w_reg_N264 ), .CK(clk), .Q(w_q[261]), .QN());
DFF_X2 _w_reg_q_reg_262_  ( .D(_w_reg_N265 ), .CK(clk), .Q(w_q[262]), .QN());
DFF_X2 _w_reg_q_reg_263_  ( .D(_w_reg_N266 ), .CK(clk), .Q(w_q[263]), .QN());
DFF_X2 _w_reg_q_reg_264_  ( .D(_w_reg_N267 ), .CK(clk), .Q(w_q[264]), .QN());
DFF_X2 _w_reg_q_reg_265_  ( .D(_w_reg_N268 ), .CK(clk), .Q(w_q[265]), .QN());
DFF_X2 _w_reg_q_reg_266_  ( .D(_w_reg_N269 ), .CK(clk), .Q(w_q[266]), .QN());
DFF_X2 _w_reg_q_reg_267_  ( .D(_w_reg_N270 ), .CK(clk), .Q(w_q[267]), .QN());
DFF_X2 _w_reg_q_reg_268_  ( .D(_w_reg_N271 ), .CK(clk), .Q(w_q[268]), .QN());
DFF_X2 _w_reg_q_reg_269_  ( .D(_w_reg_N272 ), .CK(clk), .Q(w_q[269]), .QN());
DFF_X2 _w_reg_q_reg_270_  ( .D(_w_reg_N273 ), .CK(clk), .Q(w_q[270]), .QN());
DFF_X2 _w_reg_q_reg_271_  ( .D(_w_reg_N274 ), .CK(clk), .Q(w_q[271]), .QN());
DFF_X2 _w_reg_q_reg_272_  ( .D(_w_reg_N275 ), .CK(clk), .Q(w_q[272]), .QN());
DFF_X2 _w_reg_q_reg_273_  ( .D(_w_reg_N276 ), .CK(clk), .Q(w_q[273]), .QN());
DFF_X2 _w_reg_q_reg_274_  ( .D(_w_reg_N277 ), .CK(clk), .Q(w_q[274]), .QN());
DFF_X2 _w_reg_q_reg_275_  ( .D(_w_reg_N278 ), .CK(clk), .Q(w_q[275]), .QN());
DFF_X2 _w_reg_q_reg_276_  ( .D(_w_reg_N279 ), .CK(clk), .Q(w_q[276]), .QN());
DFF_X2 _w_reg_q_reg_277_  ( .D(_w_reg_N280 ), .CK(clk), .Q(w_q[277]), .QN());
DFF_X2 _w_reg_q_reg_278_  ( .D(_w_reg_N281 ), .CK(clk), .Q(w_q[278]), .QN());
DFF_X2 _w_reg_q_reg_279_  ( .D(_w_reg_N282 ), .CK(clk), .Q(w_q[279]), .QN());
DFF_X2 _w_reg_q_reg_280_  ( .D(_w_reg_N283 ), .CK(clk), .Q(w_q[280]), .QN());
DFF_X2 _w_reg_q_reg_281_  ( .D(_w_reg_N284 ), .CK(clk), .Q(w_q[281]), .QN());
DFF_X2 _w_reg_q_reg_282_  ( .D(_w_reg_N285 ), .CK(clk), .Q(w_q[282]), .QN());
DFF_X2 _w_reg_q_reg_283_  ( .D(_w_reg_N286 ), .CK(clk), .Q(w_q[283]), .QN());
DFF_X2 _w_reg_q_reg_284_  ( .D(_w_reg_N287 ), .CK(clk), .Q(w_q[284]), .QN());
DFF_X2 _w_reg_q_reg_285_  ( .D(_w_reg_N288 ), .CK(clk), .Q(w_q[285]), .QN());
DFF_X2 _w_reg_q_reg_286_  ( .D(_w_reg_N289 ), .CK(clk), .Q(w_q[286]), .QN());
DFF_X2 _w_reg_q_reg_287_  ( .D(_w_reg_N290 ), .CK(clk), .Q(w_q[287]), .QN());
DFF_X2 _w_reg_q_reg_288_  ( .D(_w_reg_N291 ), .CK(clk), .Q(w_q[288]), .QN());
DFF_X2 _w_reg_q_reg_289_  ( .D(_w_reg_N292 ), .CK(clk), .Q(w_q[289]), .QN());
DFF_X2 _w_reg_q_reg_290_  ( .D(_w_reg_N293 ), .CK(clk), .Q(w_q[290]), .QN());
DFF_X2 _w_reg_q_reg_291_  ( .D(_w_reg_N294 ), .CK(clk), .Q(w_q[291]), .QN());
DFF_X2 _w_reg_q_reg_292_  ( .D(_w_reg_N295 ), .CK(clk), .Q(w_q[292]), .QN());
DFF_X2 _w_reg_q_reg_293_  ( .D(_w_reg_N296 ), .CK(clk), .Q(w_q[293]), .QN());
DFF_X2 _w_reg_q_reg_294_  ( .D(_w_reg_N297 ), .CK(clk), .Q(w_q[294]), .QN());
DFF_X2 _w_reg_q_reg_295_  ( .D(_w_reg_N298 ), .CK(clk), .Q(w_q[295]), .QN());
DFF_X2 _w_reg_q_reg_296_  ( .D(_w_reg_N299 ), .CK(clk), .Q(w_q[296]), .QN());
DFF_X2 _w_reg_q_reg_297_  ( .D(_w_reg_N300 ), .CK(clk), .Q(w_q[297]), .QN());
DFF_X2 _w_reg_q_reg_298_  ( .D(_w_reg_N301 ), .CK(clk), .Q(w_q[298]), .QN());
DFF_X2 _w_reg_q_reg_299_  ( .D(_w_reg_N302 ), .CK(clk), .Q(w_q[299]), .QN());
DFF_X2 _w_reg_q_reg_300_  ( .D(_w_reg_N303 ), .CK(clk), .Q(w_q[300]), .QN());
DFF_X2 _w_reg_q_reg_301_  ( .D(_w_reg_N304 ), .CK(clk), .Q(w_q[301]), .QN());
DFF_X2 _w_reg_q_reg_302_  ( .D(_w_reg_N305 ), .CK(clk), .Q(w_q[302]), .QN());
DFF_X2 _w_reg_q_reg_303_  ( .D(_w_reg_N306 ), .CK(clk), .Q(w_q[303]), .QN());
DFF_X2 _w_reg_q_reg_304_  ( .D(_w_reg_N307 ), .CK(clk), .Q(w_q[304]), .QN());
DFF_X2 _w_reg_q_reg_305_  ( .D(_w_reg_N308 ), .CK(clk), .Q(w_q[305]), .QN());
DFF_X2 _w_reg_q_reg_306_  ( .D(_w_reg_N309 ), .CK(clk), .Q(w_q[306]), .QN());
DFF_X2 _w_reg_q_reg_307_  ( .D(_w_reg_N310 ), .CK(clk), .Q(w_q[307]), .QN());
DFF_X2 _w_reg_q_reg_308_  ( .D(_w_reg_N311 ), .CK(clk), .Q(w_q[308]), .QN());
DFF_X2 _w_reg_q_reg_309_  ( .D(_w_reg_N312 ), .CK(clk), .Q(w_q[309]), .QN());
DFF_X2 _w_reg_q_reg_310_  ( .D(_w_reg_N313 ), .CK(clk), .Q(w_q[310]), .QN());
DFF_X2 _w_reg_q_reg_311_  ( .D(_w_reg_N314 ), .CK(clk), .Q(w_q[311]), .QN());
DFF_X2 _w_reg_q_reg_312_  ( .D(_w_reg_N315 ), .CK(clk), .Q(w_q[312]), .QN());
DFF_X2 _w_reg_q_reg_313_  ( .D(_w_reg_N316 ), .CK(clk), .Q(w_q[313]), .QN());
DFF_X2 _w_reg_q_reg_314_  ( .D(_w_reg_N317 ), .CK(clk), .Q(w_q[314]), .QN());
DFF_X2 _w_reg_q_reg_315_  ( .D(_w_reg_N318 ), .CK(clk), .Q(w_q[315]), .QN());
DFF_X2 _w_reg_q_reg_316_  ( .D(_w_reg_N319 ), .CK(clk), .Q(w_q[316]), .QN());
DFF_X2 _w_reg_q_reg_317_  ( .D(_w_reg_N320 ), .CK(clk), .Q(w_q[317]), .QN());
DFF_X2 _w_reg_q_reg_318_  ( .D(_w_reg_N321 ), .CK(clk), .Q(w_q[318]), .QN());
DFF_X2 _w_reg_q_reg_319_  ( .D(_w_reg_N322 ), .CK(clk), .Q(w_q[319]), .QN());
DFF_X2 _w_reg_q_reg_320_  ( .D(_w_reg_N323 ), .CK(clk), .Q(w_q[320]), .QN());
DFF_X2 _w_reg_q_reg_321_  ( .D(_w_reg_N324 ), .CK(clk), .Q(w_q[321]), .QN());
DFF_X2 _w_reg_q_reg_322_  ( .D(_w_reg_N325 ), .CK(clk), .Q(w_q[322]), .QN());
DFF_X2 _w_reg_q_reg_323_  ( .D(_w_reg_N326 ), .CK(clk), .Q(w_q[323]), .QN());
DFF_X2 _w_reg_q_reg_324_  ( .D(_w_reg_N327 ), .CK(clk), .Q(w_q[324]), .QN());
DFF_X2 _w_reg_q_reg_325_  ( .D(_w_reg_N328 ), .CK(clk), .Q(w_q[325]), .QN());
DFF_X2 _w_reg_q_reg_326_  ( .D(_w_reg_N329 ), .CK(clk), .Q(w_q[326]), .QN());
DFF_X2 _w_reg_q_reg_327_  ( .D(_w_reg_N330 ), .CK(clk), .Q(w_q[327]), .QN());
DFF_X2 _w_reg_q_reg_328_  ( .D(_w_reg_N331 ), .CK(clk), .Q(w_q[328]), .QN());
DFF_X2 _w_reg_q_reg_329_  ( .D(_w_reg_N332 ), .CK(clk), .Q(w_q[329]), .QN());
DFF_X2 _w_reg_q_reg_330_  ( .D(_w_reg_N333 ), .CK(clk), .Q(w_q[330]), .QN());
DFF_X2 _w_reg_q_reg_331_  ( .D(_w_reg_N334 ), .CK(clk), .Q(w_q[331]), .QN());
DFF_X2 _w_reg_q_reg_332_  ( .D(_w_reg_N335 ), .CK(clk), .Q(w_q[332]), .QN());
DFF_X2 _w_reg_q_reg_333_  ( .D(_w_reg_N336 ), .CK(clk), .Q(w_q[333]), .QN());
DFF_X2 _w_reg_q_reg_334_  ( .D(_w_reg_N337 ), .CK(clk), .Q(w_q[334]), .QN());
DFF_X2 _w_reg_q_reg_335_  ( .D(_w_reg_N338 ), .CK(clk), .Q(w_q[335]), .QN());
DFF_X2 _w_reg_q_reg_336_  ( .D(_w_reg_N339 ), .CK(clk), .Q(w_q[336]), .QN());
DFF_X2 _w_reg_q_reg_337_  ( .D(_w_reg_N340 ), .CK(clk), .Q(w_q[337]), .QN());
DFF_X2 _w_reg_q_reg_338_  ( .D(_w_reg_N341 ), .CK(clk), .Q(w_q[338]), .QN());
DFF_X2 _w_reg_q_reg_339_  ( .D(_w_reg_N342 ), .CK(clk), .Q(w_q[339]), .QN());
DFF_X2 _w_reg_q_reg_340_  ( .D(_w_reg_N343 ), .CK(clk), .Q(w_q[340]), .QN());
DFF_X2 _w_reg_q_reg_341_  ( .D(_w_reg_N344 ), .CK(clk), .Q(w_q[341]), .QN());
DFF_X2 _w_reg_q_reg_342_  ( .D(_w_reg_N345 ), .CK(clk), .Q(w_q[342]), .QN());
DFF_X2 _w_reg_q_reg_343_  ( .D(_w_reg_N346 ), .CK(clk), .Q(w_q[343]), .QN());
DFF_X2 _w_reg_q_reg_344_  ( .D(_w_reg_N347 ), .CK(clk), .Q(w_q[344]), .QN());
DFF_X2 _w_reg_q_reg_345_  ( .D(_w_reg_N348 ), .CK(clk), .Q(w_q[345]), .QN());
DFF_X2 _w_reg_q_reg_346_  ( .D(_w_reg_N349 ), .CK(clk), .Q(w_q[346]), .QN());
DFF_X2 _w_reg_q_reg_347_  ( .D(_w_reg_N350 ), .CK(clk), .Q(w_q[347]), .QN());
DFF_X2 _w_reg_q_reg_348_  ( .D(_w_reg_N351 ), .CK(clk), .Q(w_q[348]), .QN());
DFF_X2 _w_reg_q_reg_349_  ( .D(_w_reg_N352 ), .CK(clk), .Q(w_q[349]), .QN());
DFF_X2 _w_reg_q_reg_350_  ( .D(_w_reg_N353 ), .CK(clk), .Q(w_q[350]), .QN());
DFF_X2 _w_reg_q_reg_351_  ( .D(_w_reg_N354 ), .CK(clk), .Q(w_q[351]), .QN());
DFF_X2 _w_reg_q_reg_352_  ( .D(_w_reg_N355 ), .CK(clk), .Q(w_q[352]), .QN());
DFF_X2 _w_reg_q_reg_353_  ( .D(_w_reg_N356 ), .CK(clk), .Q(w_q[353]), .QN());
DFF_X2 _w_reg_q_reg_354_  ( .D(_w_reg_N357 ), .CK(clk), .Q(w_q[354]), .QN());
DFF_X2 _w_reg_q_reg_355_  ( .D(_w_reg_N358 ), .CK(clk), .Q(w_q[355]), .QN());
DFF_X2 _w_reg_q_reg_356_  ( .D(_w_reg_N359 ), .CK(clk), .Q(w_q[356]), .QN());
DFF_X2 _w_reg_q_reg_357_  ( .D(_w_reg_N360 ), .CK(clk), .Q(w_q[357]), .QN());
DFF_X2 _w_reg_q_reg_358_  ( .D(_w_reg_N361 ), .CK(clk), .Q(w_q[358]), .QN());
DFF_X2 _w_reg_q_reg_359_  ( .D(_w_reg_N362 ), .CK(clk), .Q(w_q[359]), .QN());
DFF_X2 _w_reg_q_reg_360_  ( .D(_w_reg_N363 ), .CK(clk), .Q(w_q[360]), .QN());
DFF_X2 _w_reg_q_reg_361_  ( .D(_w_reg_N364 ), .CK(clk), .Q(w_q[361]), .QN());
DFF_X2 _w_reg_q_reg_362_  ( .D(_w_reg_N365 ), .CK(clk), .Q(w_q[362]), .QN());
DFF_X2 _w_reg_q_reg_363_  ( .D(_w_reg_N366 ), .CK(clk), .Q(w_q[363]), .QN());
DFF_X2 _w_reg_q_reg_364_  ( .D(_w_reg_N367 ), .CK(clk), .Q(w_q[364]), .QN());
DFF_X2 _w_reg_q_reg_365_  ( .D(_w_reg_N368 ), .CK(clk), .Q(w_q[365]), .QN());
DFF_X2 _w_reg_q_reg_366_  ( .D(_w_reg_N369 ), .CK(clk), .Q(w_q[366]), .QN());
DFF_X2 _w_reg_q_reg_367_  ( .D(_w_reg_N370 ), .CK(clk), .Q(w_q[367]), .QN());
DFF_X2 _w_reg_q_reg_368_  ( .D(_w_reg_N371 ), .CK(clk), .Q(w_q[368]), .QN());
DFF_X2 _w_reg_q_reg_369_  ( .D(_w_reg_N372 ), .CK(clk), .Q(w_q[369]), .QN());
DFF_X2 _w_reg_q_reg_370_  ( .D(_w_reg_N373 ), .CK(clk), .Q(w_q[370]), .QN());
DFF_X2 _w_reg_q_reg_371_  ( .D(_w_reg_N374 ), .CK(clk), .Q(w_q[371]), .QN());
DFF_X2 _w_reg_q_reg_372_  ( .D(_w_reg_N375 ), .CK(clk), .Q(w_q[372]), .QN());
DFF_X2 _w_reg_q_reg_373_  ( .D(_w_reg_N376 ), .CK(clk), .Q(w_q[373]), .QN());
DFF_X2 _w_reg_q_reg_374_  ( .D(_w_reg_N377 ), .CK(clk), .Q(w_q[374]), .QN());
DFF_X2 _w_reg_q_reg_375_  ( .D(_w_reg_N378 ), .CK(clk), .Q(w_q[375]), .QN());
DFF_X2 _w_reg_q_reg_376_  ( .D(_w_reg_N379 ), .CK(clk), .Q(w_q[376]), .QN());
DFF_X2 _w_reg_q_reg_377_  ( .D(_w_reg_N380 ), .CK(clk), .Q(w_q[377]), .QN());
DFF_X2 _w_reg_q_reg_378_  ( .D(_w_reg_N381 ), .CK(clk), .Q(w_q[378]), .QN());
DFF_X2 _w_reg_q_reg_379_  ( .D(_w_reg_N382 ), .CK(clk), .Q(w_q[379]), .QN());
DFF_X2 _w_reg_q_reg_380_  ( .D(_w_reg_N383 ), .CK(clk), .Q(w_q[380]), .QN());
DFF_X2 _w_reg_q_reg_381_  ( .D(_w_reg_N384 ), .CK(clk), .Q(w_q[381]), .QN());
DFF_X2 _w_reg_q_reg_382_  ( .D(_w_reg_N385 ), .CK(clk), .Q(w_q[382]), .QN());
DFF_X2 _w_reg_q_reg_383_  ( .D(_w_reg_N386 ), .CK(clk), .Q(w_q[383]), .QN());
DFF_X2 _w_reg_q_reg_384_  ( .D(_w_reg_N387 ), .CK(clk), .Q(w_q[384]), .QN());
DFF_X2 _w_reg_q_reg_385_  ( .D(_w_reg_N388 ), .CK(clk), .Q(w_q[385]), .QN());
DFF_X2 _w_reg_q_reg_386_  ( .D(_w_reg_N389 ), .CK(clk), .Q(w_q[386]), .QN());
DFF_X2 _w_reg_q_reg_387_  ( .D(_w_reg_N390 ), .CK(clk), .Q(w_q[387]), .QN());
DFF_X2 _w_reg_q_reg_388_  ( .D(_w_reg_N391 ), .CK(clk), .Q(w_q[388]), .QN());
DFF_X2 _w_reg_q_reg_389_  ( .D(_w_reg_N392 ), .CK(clk), .Q(w_q[389]), .QN());
DFF_X2 _w_reg_q_reg_390_  ( .D(_w_reg_N393 ), .CK(clk), .Q(w_q[390]), .QN());
DFF_X2 _w_reg_q_reg_391_  ( .D(_w_reg_N394 ), .CK(clk), .Q(w_q[391]), .QN());
DFF_X2 _w_reg_q_reg_392_  ( .D(_w_reg_N395 ), .CK(clk), .Q(w_q[392]), .QN());
DFF_X2 _w_reg_q_reg_393_  ( .D(_w_reg_N396 ), .CK(clk), .Q(w_q[393]), .QN());
DFF_X2 _w_reg_q_reg_394_  ( .D(_w_reg_N397 ), .CK(clk), .Q(w_q[394]), .QN());
DFF_X2 _w_reg_q_reg_395_  ( .D(_w_reg_N398 ), .CK(clk), .Q(w_q[395]), .QN());
DFF_X2 _w_reg_q_reg_396_  ( .D(_w_reg_N399 ), .CK(clk), .Q(w_q[396]), .QN());
DFF_X2 _w_reg_q_reg_397_  ( .D(_w_reg_N400 ), .CK(clk), .Q(w_q[397]), .QN());
DFF_X2 _w_reg_q_reg_398_  ( .D(_w_reg_N401 ), .CK(clk), .Q(w_q[398]), .QN());
DFF_X2 _w_reg_q_reg_399_  ( .D(_w_reg_N402 ), .CK(clk), .Q(w_q[399]), .QN());
DFF_X2 _w_reg_q_reg_400_  ( .D(_w_reg_N403 ), .CK(clk), .Q(w_q[400]), .QN());
DFF_X2 _w_reg_q_reg_401_  ( .D(_w_reg_N404 ), .CK(clk), .Q(w_q[401]), .QN());
DFF_X2 _w_reg_q_reg_402_  ( .D(_w_reg_N405 ), .CK(clk), .Q(w_q[402]), .QN());
DFF_X2 _w_reg_q_reg_403_  ( .D(_w_reg_N406 ), .CK(clk), .Q(w_q[403]), .QN());
DFF_X2 _w_reg_q_reg_404_  ( .D(_w_reg_N407 ), .CK(clk), .Q(w_q[404]), .QN());
DFF_X2 _w_reg_q_reg_405_  ( .D(_w_reg_N408 ), .CK(clk), .Q(w_q[405]), .QN());
DFF_X2 _w_reg_q_reg_406_  ( .D(_w_reg_N409 ), .CK(clk), .Q(w_q[406]), .QN());
DFF_X2 _w_reg_q_reg_407_  ( .D(_w_reg_N410 ), .CK(clk), .Q(w_q[407]), .QN());
DFF_X2 _w_reg_q_reg_408_  ( .D(_w_reg_N411 ), .CK(clk), .Q(w_q[408]), .QN());
DFF_X2 _w_reg_q_reg_409_  ( .D(_w_reg_N412 ), .CK(clk), .Q(w_q[409]), .QN());
DFF_X2 _w_reg_q_reg_410_  ( .D(_w_reg_N413 ), .CK(clk), .Q(w_q[410]), .QN());
DFF_X2 _w_reg_q_reg_411_  ( .D(_w_reg_N414 ), .CK(clk), .Q(w_q[411]), .QN());
DFF_X2 _w_reg_q_reg_412_  ( .D(_w_reg_N415 ), .CK(clk), .Q(w_q[412]), .QN());
DFF_X2 _w_reg_q_reg_413_  ( .D(_w_reg_N416 ), .CK(clk), .Q(w_q[413]), .QN());
DFF_X2 _w_reg_q_reg_414_  ( .D(_w_reg_N417 ), .CK(clk), .Q(w_q[414]), .QN());
DFF_X2 _w_reg_q_reg_415_  ( .D(_w_reg_N418 ), .CK(clk), .Q(w_q[415]), .QN());
DFF_X2 _w_reg_q_reg_416_  ( .D(_w_reg_N419 ), .CK(clk), .Q(w_q[416]), .QN());
DFF_X2 _w_reg_q_reg_417_  ( .D(_w_reg_N420 ), .CK(clk), .Q(w_q[417]), .QN());
DFF_X2 _w_reg_q_reg_418_  ( .D(_w_reg_N421 ), .CK(clk), .Q(w_q[418]), .QN());
DFF_X2 _w_reg_q_reg_419_  ( .D(_w_reg_N422 ), .CK(clk), .Q(w_q[419]), .QN());
DFF_X2 _w_reg_q_reg_420_  ( .D(_w_reg_N423 ), .CK(clk), .Q(w_q[420]), .QN());
DFF_X2 _w_reg_q_reg_421_  ( .D(_w_reg_N424 ), .CK(clk), .Q(w_q[421]), .QN());
DFF_X2 _w_reg_q_reg_422_  ( .D(_w_reg_N425 ), .CK(clk), .Q(w_q[422]), .QN());
DFF_X2 _w_reg_q_reg_423_  ( .D(_w_reg_N426 ), .CK(clk), .Q(w_q[423]), .QN());
DFF_X2 _w_reg_q_reg_424_  ( .D(_w_reg_N427 ), .CK(clk), .Q(w_q[424]), .QN());
DFF_X2 _w_reg_q_reg_425_  ( .D(_w_reg_N428 ), .CK(clk), .Q(w_q[425]), .QN());
DFF_X2 _w_reg_q_reg_426_  ( .D(_w_reg_N429 ), .CK(clk), .Q(w_q[426]), .QN());
DFF_X2 _w_reg_q_reg_427_  ( .D(_w_reg_N430 ), .CK(clk), .Q(w_q[427]), .QN());
DFF_X2 _w_reg_q_reg_428_  ( .D(_w_reg_N431 ), .CK(clk), .Q(w_q[428]), .QN());
DFF_X2 _w_reg_q_reg_429_  ( .D(_w_reg_N432 ), .CK(clk), .Q(w_q[429]), .QN());
DFF_X2 _w_reg_q_reg_430_  ( .D(_w_reg_N433 ), .CK(clk), .Q(w_q[430]), .QN());
DFF_X2 _w_reg_q_reg_431_  ( .D(_w_reg_N434 ), .CK(clk), .Q(w_q[431]), .QN());
DFF_X2 _w_reg_q_reg_432_  ( .D(_w_reg_N435 ), .CK(clk), .Q(w_q[432]), .QN());
DFF_X2 _w_reg_q_reg_433_  ( .D(_w_reg_N436 ), .CK(clk), .Q(w_q[433]), .QN());
DFF_X2 _w_reg_q_reg_434_  ( .D(_w_reg_N437 ), .CK(clk), .Q(w_q[434]), .QN());
DFF_X2 _w_reg_q_reg_435_  ( .D(_w_reg_N438 ), .CK(clk), .Q(w_q[435]), .QN());
DFF_X2 _w_reg_q_reg_436_  ( .D(_w_reg_N439 ), .CK(clk), .Q(w_q[436]), .QN());
DFF_X2 _w_reg_q_reg_437_  ( .D(_w_reg_N440 ), .CK(clk), .Q(w_q[437]), .QN());
DFF_X2 _w_reg_q_reg_438_  ( .D(_w_reg_N441 ), .CK(clk), .Q(w_q[438]), .QN());
DFF_X2 _w_reg_q_reg_439_  ( .D(_w_reg_N442 ), .CK(clk), .Q(w_q[439]), .QN());
DFF_X2 _w_reg_q_reg_440_  ( .D(_w_reg_N443 ), .CK(clk), .Q(w_q[440]), .QN());
DFF_X2 _w_reg_q_reg_441_  ( .D(_w_reg_N444 ), .CK(clk), .Q(w_q[441]), .QN());
DFF_X2 _w_reg_q_reg_442_  ( .D(_w_reg_N445 ), .CK(clk), .Q(w_q[442]), .QN());
DFF_X2 _w_reg_q_reg_443_  ( .D(_w_reg_N446 ), .CK(clk), .Q(w_q[443]), .QN());
DFF_X2 _w_reg_q_reg_444_  ( .D(_w_reg_N447 ), .CK(clk), .Q(w_q[444]), .QN());
DFF_X2 _w_reg_q_reg_445_  ( .D(_w_reg_N448 ), .CK(clk), .Q(w_q[445]), .QN());
DFF_X2 _w_reg_q_reg_446_  ( .D(_w_reg_N449 ), .CK(clk), .Q(w_q[446]), .QN());
DFF_X2 _w_reg_q_reg_447_  ( .D(_w_reg_N450 ), .CK(clk), .Q(w_q[447]), .QN());
DFF_X2 _w_reg_q_reg_448_  ( .D(_w_reg_N451 ), .CK(clk), .Q(w_q[448]), .QN());
DFF_X2 _w_reg_q_reg_449_  ( .D(_w_reg_N452 ), .CK(clk), .Q(w_q[449]), .QN());
DFF_X2 _w_reg_q_reg_450_  ( .D(_w_reg_N453 ), .CK(clk), .Q(w_q[450]), .QN());
DFF_X2 _w_reg_q_reg_451_  ( .D(_w_reg_N454 ), .CK(clk), .Q(w_q[451]), .QN());
DFF_X2 _w_reg_q_reg_452_  ( .D(_w_reg_N455 ), .CK(clk), .Q(w_q[452]), .QN());
DFF_X2 _w_reg_q_reg_453_  ( .D(_w_reg_N456 ), .CK(clk), .Q(w_q[453]), .QN());
DFF_X2 _w_reg_q_reg_454_  ( .D(_w_reg_N457 ), .CK(clk), .Q(w_q[454]), .QN());
DFF_X2 _w_reg_q_reg_455_  ( .D(_w_reg_N458 ), .CK(clk), .Q(w_q[455]), .QN());
DFF_X2 _w_reg_q_reg_456_  ( .D(_w_reg_N459 ), .CK(clk), .Q(w_q[456]), .QN());
DFF_X2 _w_reg_q_reg_457_  ( .D(_w_reg_N460 ), .CK(clk), .Q(w_q[457]), .QN());
DFF_X2 _w_reg_q_reg_458_  ( .D(_w_reg_N461 ), .CK(clk), .Q(w_q[458]), .QN());
DFF_X2 _w_reg_q_reg_459_  ( .D(_w_reg_N462 ), .CK(clk), .Q(w_q[459]), .QN());
DFF_X2 _w_reg_q_reg_460_  ( .D(_w_reg_N463 ), .CK(clk), .Q(w_q[460]), .QN());
DFF_X2 _w_reg_q_reg_461_  ( .D(_w_reg_N464 ), .CK(clk), .Q(w_q[461]), .QN());
DFF_X2 _w_reg_q_reg_462_  ( .D(_w_reg_N465 ), .CK(clk), .Q(w_q[462]), .QN());
DFF_X2 _w_reg_q_reg_463_  ( .D(_w_reg_N466 ), .CK(clk), .Q(w_q[463]), .QN());
DFF_X2 _w_reg_q_reg_464_  ( .D(_w_reg_N467 ), .CK(clk), .Q(w_q[464]), .QN());
DFF_X2 _w_reg_q_reg_465_  ( .D(_w_reg_N468 ), .CK(clk), .Q(w_q[465]), .QN());
DFF_X2 _w_reg_q_reg_466_  ( .D(_w_reg_N469 ), .CK(clk), .Q(w_q[466]), .QN());
DFF_X2 _w_reg_q_reg_467_  ( .D(_w_reg_N470 ), .CK(clk), .Q(w_q[467]), .QN());
DFF_X2 _w_reg_q_reg_468_  ( .D(_w_reg_N471 ), .CK(clk), .Q(w_q[468]), .QN());
DFF_X2 _w_reg_q_reg_469_  ( .D(_w_reg_N472 ), .CK(clk), .Q(w_q[469]), .QN());
DFF_X2 _w_reg_q_reg_470_  ( .D(_w_reg_N473 ), .CK(clk), .Q(w_q[470]), .QN());
DFF_X2 _w_reg_q_reg_471_  ( .D(_w_reg_N474 ), .CK(clk), .Q(w_q[471]), .QN());
DFF_X2 _w_reg_q_reg_472_  ( .D(_w_reg_N475 ), .CK(clk), .Q(w_q[472]), .QN());
DFF_X2 _w_reg_q_reg_473_  ( .D(_w_reg_N476 ), .CK(clk), .Q(w_q[473]), .QN());
DFF_X2 _w_reg_q_reg_474_  ( .D(_w_reg_N477 ), .CK(clk), .Q(w_q[474]), .QN());
DFF_X2 _w_reg_q_reg_475_  ( .D(_w_reg_N478 ), .CK(clk), .Q(w_q[475]), .QN());
DFF_X2 _w_reg_q_reg_476_  ( .D(_w_reg_N479 ), .CK(clk), .Q(w_q[476]), .QN());
DFF_X2 _w_reg_q_reg_477_  ( .D(_w_reg_N480 ), .CK(clk), .Q(w_q[477]), .QN());
DFF_X2 _w_reg_q_reg_478_  ( .D(_w_reg_N481 ), .CK(clk), .Q(w_q[478]), .QN());
DFF_X2 _w_reg_q_reg_479_  ( .D(_w_reg_N482 ), .CK(clk), .Q(w_q[479]), .QN());
DFF_X2 _w_reg_q_reg_480_  ( .D(_w_reg_N483 ), .CK(clk), .Q(w[0]), .QN() );
DFF_X2 _w_reg_q_reg_481_  ( .D(_w_reg_N484 ), .CK(clk), .Q(w[1]), .QN() );
DFF_X2 _w_reg_q_reg_482_  ( .D(_w_reg_N485 ), .CK(clk), .Q(w[2]), .QN() );
DFF_X2 _w_reg_q_reg_483_  ( .D(_w_reg_N486 ), .CK(clk), .Q(w[3]), .QN() );
DFF_X2 _w_reg_q_reg_484_  ( .D(_w_reg_N487 ), .CK(clk), .Q(w[4]), .QN() );
DFF_X2 _w_reg_q_reg_485_  ( .D(_w_reg_N488 ), .CK(clk), .Q(w[5]), .QN() );
DFF_X2 _w_reg_q_reg_486_  ( .D(_w_reg_N489 ), .CK(clk), .Q(w[6]), .QN() );
DFF_X2 _w_reg_q_reg_487_  ( .D(_w_reg_N490 ), .CK(clk), .Q(w[7]), .QN() );
DFF_X2 _w_reg_q_reg_488_  ( .D(_w_reg_N491 ), .CK(clk), .Q(w[8]), .QN() );
DFF_X2 _w_reg_q_reg_489_  ( .D(_w_reg_N492 ), .CK(clk), .Q(w[9]), .QN() );
DFF_X2 _w_reg_q_reg_490_  ( .D(_w_reg_N493 ), .CK(clk), .Q(w[10]), .QN() );
DFF_X2 _w_reg_q_reg_491_  ( .D(_w_reg_N494 ), .CK(clk), .Q(w[11]), .QN() );
DFF_X2 _w_reg_q_reg_492_  ( .D(_w_reg_N495 ), .CK(clk), .Q(w[12]), .QN() );
DFF_X2 _w_reg_q_reg_493_  ( .D(_w_reg_N496 ), .CK(clk), .Q(w[13]), .QN() );
DFF_X2 _w_reg_q_reg_494_  ( .D(_w_reg_N497 ), .CK(clk), .Q(w[14]), .QN() );
DFF_X2 _w_reg_q_reg_495_  ( .D(_w_reg_N498 ), .CK(clk), .Q(w[15]), .QN() );
DFF_X2 _w_reg_q_reg_496_  ( .D(_w_reg_N499 ), .CK(clk), .Q(w[16]), .QN() );
DFF_X2 _w_reg_q_reg_497_  ( .D(_w_reg_N500 ), .CK(clk), .Q(w[17]), .QN() );
DFF_X2 _w_reg_q_reg_498_  ( .D(_w_reg_N501 ), .CK(clk), .Q(w[18]), .QN() );
DFF_X2 _w_reg_q_reg_499_  ( .D(_w_reg_N502 ), .CK(clk), .Q(w[19]), .QN() );
DFF_X2 _w_reg_q_reg_500_  ( .D(_w_reg_N503 ), .CK(clk), .Q(w[20]), .QN() );
DFF_X2 _w_reg_q_reg_501_  ( .D(_w_reg_N504 ), .CK(clk), .Q(w[21]), .QN() );
DFF_X2 _w_reg_q_reg_502_  ( .D(_w_reg_N505 ), .CK(clk), .Q(w[22]), .QN() );
DFF_X2 _w_reg_q_reg_503_  ( .D(_w_reg_N506 ), .CK(clk), .Q(w[23]), .QN() );
DFF_X2 _w_reg_q_reg_504_  ( .D(_w_reg_N507 ), .CK(clk), .Q(w[24]), .QN() );
DFF_X2 _w_reg_q_reg_505_  ( .D(_w_reg_N508 ), .CK(clk), .Q(w[25]), .QN() );
DFF_X2 _w_reg_q_reg_506_  ( .D(_w_reg_N509 ), .CK(clk), .Q(w[26]), .QN() );
DFF_X2 _w_reg_q_reg_507_  ( .D(_w_reg_N510 ), .CK(clk), .Q(w[27]), .QN() );
DFF_X2 _w_reg_q_reg_508_  ( .D(_w_reg_N511 ), .CK(clk), .Q(w[28]), .QN() );
DFF_X2 _w_reg_q_reg_509_  ( .D(_w_reg_N512 ), .CK(clk), .Q(w[29]), .QN() );
DFF_X2 _w_reg_q_reg_510_  ( .D(_w_reg_N513 ), .CK(clk), .Q(w[30]), .QN() );
DFF_X2 _w_reg_q_reg_511_  ( .D(_w_reg_N514 ), .CK(clk), .Q(w[31]), .QN() );
AND2_X2 _cv_reg_U179  ( .A1(cv_d[137]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N140 ) );
AND2_X2 _cv_reg_U178  ( .A1(cv_d[136]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N139 ) );
AND2_X2 _cv_reg_U177  ( .A1(cv_d[135]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N138 ) );
AND2_X2 _cv_reg_U176  ( .A1(cv_d[134]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N137 ) );
AND2_X2 _cv_reg_U175  ( .A1(cv_d[133]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N136 ) );
AND2_X2 _cv_reg_U174  ( .A1(cv_d[132]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N135 ) );
AND2_X2 _cv_reg_U173  ( .A1(cv_d[131]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N134 ) );
AND2_X2 _cv_reg_U172  ( .A1(cv_d[130]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N133 ) );
AND2_X2 _cv_reg_U171  ( .A1(cv_d[129]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N132 ) );
AND2_X2 _cv_reg_U170  ( .A1(cv_d[128]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N131 ) );
AND2_X2 _cv_reg_U169  ( .A1(cv_d[111]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N114 ) );
AND2_X2 _cv_reg_U168  ( .A1(cv_d[110]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N113 ) );
AND2_X2 _cv_reg_U167  ( .A1(cv_d[109]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N112 ) );
AND2_X2 _cv_reg_U166  ( .A1(cv_d[108]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N111 ) );
AND2_X2 _cv_reg_U165  ( .A1(cv_d[107]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N110 ) );
AND2_X2 _cv_reg_U164  ( .A1(cv_d[106]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N109 ) );
AND2_X2 _cv_reg_U163  ( .A1(cv_d[105]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N108 ) );
AND2_X2 _cv_reg_U162  ( .A1(cv_d[104]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N107 ) );
AND2_X2 _cv_reg_U161  ( .A1(cv_d[103]), .A2(_cv_reg_n220 ), .ZN(_cv_reg_N106 ) );
AND2_X2 _cv_reg_U160  ( .A1(cv_d[102]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N105 ) );
AND2_X2 _cv_reg_U159  ( .A1(cv_d[101]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N104 ) );
AND2_X2 _cv_reg_U158  ( .A1(cv_d[100]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N103 ) );
AND2_X2 _cv_reg_U157  ( .A1(cv_d[99]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N102 ) );
AND2_X2 _cv_reg_U156  ( .A1(cv_d[98]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N101 ) );
AND2_X2 _cv_reg_U155  ( .A1(cv_d[97]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N100 ) );
AND2_X2 _cv_reg_U154  ( .A1(cv_d[96]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N99 ));
AND2_X2 _cv_reg_U153  ( .A1(cv_d[79]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N82 ));
AND2_X2 _cv_reg_U152  ( .A1(cv_d[78]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N81 ));
AND2_X2 _cv_reg_U151  ( .A1(cv_d[77]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N80 ));
AND2_X2 _cv_reg_U150  ( .A1(cv_d[76]), .A2(_cv_reg_n210 ), .ZN(_cv_reg_N79 ));
AND2_X2 _cv_reg_U149  ( .A1(cv_d[75]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N78 ));
AND2_X2 _cv_reg_U148  ( .A1(cv_d[74]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N77 ));
AND2_X2 _cv_reg_U147  ( .A1(cv_d[73]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N76 ));
AND2_X2 _cv_reg_U146  ( .A1(cv_d[72]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N75 ));
AND2_X2 _cv_reg_U140  ( .A1(cv_d[71]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N74 ));
AND2_X2 _cv_reg_U129  ( .A1(cv_d[70]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N73 ));
AND2_X2 _cv_reg_U127  ( .A1(cv_d[69]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N72 ));
AND2_X2 _cv_reg_U126  ( .A1(cv_d[68]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N71 ));
AND2_X2 _cv_reg_U125  ( .A1(cv_d[67]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N70 ));
AND2_X2 _cv_reg_U124  ( .A1(cv_d[66]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N69 ));
AND2_X2 _cv_reg_U123  ( .A1(cv_d[65]), .A2(_cv_reg_n200 ), .ZN(_cv_reg_N68 ));
AND2_X2 _cv_reg_U122  ( .A1(cv_d[64]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N67 ));
AND2_X2 _cv_reg_U121  ( .A1(cv_d[47]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N50 ));
AND2_X2 _cv_reg_U120  ( .A1(cv_d[46]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N49 ));
AND2_X2 _cv_reg_U119  ( .A1(cv_d[45]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N48 ));
AND2_X2 _cv_reg_U118  ( .A1(cv_d[44]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N47 ));
AND2_X2 _cv_reg_U117  ( .A1(cv_d[43]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N46 ));
AND2_X2 _cv_reg_U116  ( .A1(cv_d[42]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N45 ));
AND2_X2 _cv_reg_U115  ( .A1(cv_d[41]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N44 ));
AND2_X2 _cv_reg_U114  ( .A1(cv_d[40]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N43 ));
AND2_X2 _cv_reg_U113  ( .A1(cv_d[39]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N42 ));
AND2_X2 _cv_reg_U112  ( .A1(cv_d[38]), .A2(_cv_reg_n190 ), .ZN(_cv_reg_N41 ));
AND2_X2 _cv_reg_U111  ( .A1(cv_d[37]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N40 ));
AND2_X2 _cv_reg_U110  ( .A1(cv_d[36]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N39 ));
AND2_X2 _cv_reg_U109  ( .A1(cv_d[35]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N38 ));
AND2_X2 _cv_reg_U108  ( .A1(cv_d[34]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N37 ));
AND2_X2 _cv_reg_U107  ( .A1(cv_d[33]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N36 ));
AND2_X2 _cv_reg_U106  ( .A1(cv_d[32]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N35 ));
AND2_X2 _cv_reg_U105  ( .A1(cv_d[15]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N18 ));
AND2_X2 _cv_reg_U102  ( .A1(cv_d[14]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N17 ));
AND2_X2 _cv_reg_U101  ( .A1(cv_d[13]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N16 ));
AND2_X2 _cv_reg_U97  ( .A1(cv_d[12]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N15 ));
AND2_X2 _cv_reg_U96  ( .A1(cv_d[11]), .A2(_cv_reg_n180 ), .ZN(_cv_reg_N14 ));
AND2_X2 _cv_reg_U95  ( .A1(cv_d[10]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N13 ));
AND2_X2 _cv_reg_U92  ( .A1(cv_d[9]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N12 ));
AND2_X2 _cv_reg_U91  ( .A1(cv_d[8]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N11 ));
AND2_X2 _cv_reg_U79  ( .A1(cv_d[7]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N10 ));
AND2_X2 _cv_reg_U73  ( .A1(cv_d[6]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N9 ) );
AND2_X2 _cv_reg_U72  ( .A1(cv_d[5]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N8 ) );
AND2_X2 _cv_reg_U71  ( .A1(cv_d[4]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N7 ) );
AND2_X2 _cv_reg_U70  ( .A1(cv_d[3]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N6 ) );
AND2_X2 _cv_reg_U69  ( .A1(cv_d[2]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N5 ) );
AND2_X2 _cv_reg_U68  ( .A1(cv_d[1]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N4 ) );
AND2_X2 _cv_reg_U67  ( .A1(cv_d[0]), .A2(_cv_reg_n170 ), .ZN(_cv_reg_N3 ) );
INV_X4 _cv_reg_U66  ( .A(n7117), .ZN(_cv_reg_n330 ) );
INV_X4 _cv_reg_U65  ( .A(_cv_reg_n330 ), .ZN(_cv_reg_n320 ) );
INV_X4 _cv_reg_U64  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n310 ) );
INV_X4 _cv_reg_U63  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n220 ) );
INV_X4 _cv_reg_U62  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n210 ) );
INV_X4 _cv_reg_U61  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n200 ) );
INV_X4 _cv_reg_U60  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n190 ) );
INV_X4 _cv_reg_U59  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n180 ) );
INV_X4 _cv_reg_U58  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n170 ) );
INV_X4 _cv_reg_U57  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n280 ) );
INV_X4 _cv_reg_U56  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n290 ) );
INV_X4 _cv_reg_U46  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n300 ) );
INV_X4 _cv_reg_U38  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n240 ) );
INV_X4 _cv_reg_U37  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n230 ) );
INV_X4 _cv_reg_U36  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n250 ) );
INV_X4 _cv_reg_U35  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n260 ) );
INV_X4 _cv_reg_U34  ( .A(_cv_reg_n320 ), .ZN(_cv_reg_n270 ) );
AND2_X1 _cv_reg_U33  ( .A1(cv_d[157]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N160 ) );
AND2_X1 _cv_reg_U32  ( .A1(cv_d[156]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N159 ) );
AND2_X1 _cv_reg_U31  ( .A1(cv_d[152]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N155 ) );
AND2_X1 _cv_reg_U30  ( .A1(cv_d[151]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N154 ) );
AND2_X1 _cv_reg_U29  ( .A1(cv_d[148]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N151 ) );
AND2_X1 _cv_reg_U28  ( .A1(cv_d[147]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N150 ) );
AND2_X1 _cv_reg_U27  ( .A1(cv_d[146]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N149 ) );
AND2_X1 _cv_reg_U26  ( .A1(cv_d[145]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N148 ) );
AND2_X1 _cv_reg_U25  ( .A1(cv_d[144]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N147 ) );
AND2_X1 _cv_reg_U24  ( .A1(cv_d[143]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N146 ) );
AND2_X1 _cv_reg_U23  ( .A1(cv_d[142]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N145 ) );
AND2_X1 _cv_reg_U22  ( .A1(cv_d[141]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N144 ) );
AND2_X1 _cv_reg_U21  ( .A1(cv_d[140]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N143 ) );
AND2_X1 _cv_reg_U13  ( .A1(cv_d[139]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N142 ) );
AND2_X1 _cv_reg_U3  ( .A1(cv_d[138]), .A2(_cv_reg_n230 ), .ZN(_cv_reg_N141 ));
AND2_X2 _cv_reg_U145  ( .A1(cv_d[112]), .A2(_cv_reg_n310 ), .ZN(_cv_reg_N115 ) );
AND2_X2 _cv_reg_U144  ( .A1(cv_d[113]), .A2(_cv_reg_n310 ), .ZN(_cv_reg_N116 ) );
AND2_X2 _cv_reg_U143  ( .A1(cv_d[114]), .A2(_cv_reg_n310 ), .ZN(_cv_reg_N117 ) );
AND2_X2 _cv_reg_U142  ( .A1(cv_d[115]), .A2(_cv_reg_n310 ), .ZN(_cv_reg_N118 ) );
AND2_X2 _cv_reg_U141  ( .A1(cv_d[116]), .A2(_cv_reg_n310 ), .ZN(_cv_reg_N119 ) );
AND2_X2 _cv_reg_U139  ( .A1(cv_d[117]), .A2(_cv_reg_n310 ), .ZN(_cv_reg_N120 ) );
AND2_X2 _cv_reg_U138  ( .A1(cv_d[118]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N121 ) );
AND2_X2 _cv_reg_U137  ( .A1(cv_d[119]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N122 ) );
AND2_X2 _cv_reg_U136  ( .A1(cv_d[120]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N123 ) );
AND2_X2 _cv_reg_U135  ( .A1(cv_d[121]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N124 ) );
AND2_X2 _cv_reg_U134  ( .A1(cv_d[122]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N125 ) );
AND2_X2 _cv_reg_U133  ( .A1(cv_d[123]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N126 ) );
AND2_X2 _cv_reg_U132  ( .A1(cv_d[124]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N127 ) );
AND2_X2 _cv_reg_U131  ( .A1(cv_d[125]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N128 ) );
AND2_X2 _cv_reg_U130  ( .A1(cv_d[126]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N129 ) );
AND2_X2 _cv_reg_U128  ( .A1(cv_d[127]), .A2(_cv_reg_n300 ), .ZN(_cv_reg_N130 ) );
AND2_X2 _cv_reg_U104  ( .A1(cv_d[149]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N152 ) );
AND2_X2 _cv_reg_U103  ( .A1(cv_d[150]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N153 ) );
AND2_X2 _cv_reg_U100  ( .A1(cv_d[153]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N156 ) );
AND2_X2 _cv_reg_U99  ( .A1(cv_d[154]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N157 ) );
AND2_X2 _cv_reg_U98  ( .A1(cv_d[155]), .A2(_cv_reg_n290 ), .ZN(_cv_reg_N158 ) );
AND2_X2 _cv_reg_U94  ( .A1(cv_d[158]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N161 ) );
AND2_X2 _cv_reg_U93  ( .A1(cv_d[159]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N162 ) );
AND2_X2 _cv_reg_U90  ( .A1(cv_d[16]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N19 ));
AND2_X2 _cv_reg_U89  ( .A1(cv_d[17]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N20 ));
AND2_X2 _cv_reg_U88  ( .A1(cv_d[18]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N21 ));
AND2_X2 _cv_reg_U87  ( .A1(cv_d[19]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N22 ));
AND2_X2 _cv_reg_U86  ( .A1(cv_d[20]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N23 ));
AND2_X2 _cv_reg_U85  ( .A1(cv_d[21]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N24 ));
AND2_X2 _cv_reg_U84  ( .A1(cv_d[22]), .A2(_cv_reg_n280 ), .ZN(_cv_reg_N25 ));
AND2_X2 _cv_reg_U83  ( .A1(cv_d[23]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N26 ));
AND2_X2 _cv_reg_U82  ( .A1(cv_d[24]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N27 ));
AND2_X2 _cv_reg_U81  ( .A1(cv_d[25]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N28 ));
AND2_X2 _cv_reg_U80  ( .A1(cv_d[26]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N29 ));
AND2_X2 _cv_reg_U78  ( .A1(cv_d[27]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N30 ));
AND2_X2 _cv_reg_U77  ( .A1(cv_d[28]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N31 ));
AND2_X2 _cv_reg_U76  ( .A1(cv_d[29]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N32 ));
AND2_X2 _cv_reg_U75  ( .A1(cv_d[30]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N33 ));
AND2_X2 _cv_reg_U74  ( .A1(cv_d[31]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N34 ));
AND2_X2 _cv_reg_U55  ( .A1(cv_d[48]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N51 ));
AND2_X2 _cv_reg_U54  ( .A1(cv_d[49]), .A2(_cv_reg_n270 ), .ZN(_cv_reg_N52 ));
AND2_X2 _cv_reg_U53  ( .A1(cv_d[50]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N53 ));
AND2_X2 _cv_reg_U52  ( .A1(cv_d[51]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N54 ));
AND2_X2 _cv_reg_U51  ( .A1(cv_d[52]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N55 ));
AND2_X2 _cv_reg_U50  ( .A1(cv_d[53]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N56 ));
AND2_X2 _cv_reg_U49  ( .A1(cv_d[54]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N57 ));
AND2_X2 _cv_reg_U48  ( .A1(cv_d[55]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N58 ));
AND2_X2 _cv_reg_U47  ( .A1(cv_d[56]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N59 ));
AND2_X2 _cv_reg_U45  ( .A1(cv_d[57]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N60 ));
AND2_X2 _cv_reg_U44  ( .A1(cv_d[58]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N61 ));
AND2_X2 _cv_reg_U43  ( .A1(cv_d[59]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N62 ));
AND2_X2 _cv_reg_U42  ( .A1(cv_d[60]), .A2(_cv_reg_n260 ), .ZN(_cv_reg_N63 ));
AND2_X2 _cv_reg_U41  ( .A1(cv_d[61]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N64 ));
AND2_X2 _cv_reg_U40  ( .A1(cv_d[62]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N65 ));
AND2_X2 _cv_reg_U39  ( .A1(cv_d[63]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N66 ));
AND2_X2 _cv_reg_U20  ( .A1(cv_d[80]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N83 ));
AND2_X2 _cv_reg_U19  ( .A1(cv_d[81]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N84 ));
AND2_X2 _cv_reg_U18  ( .A1(cv_d[82]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N85 ));
AND2_X2 _cv_reg_U17  ( .A1(cv_d[83]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N86 ));
AND2_X2 _cv_reg_U16  ( .A1(cv_d[84]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N87 ));
AND2_X2 _cv_reg_U15  ( .A1(cv_d[85]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N88 ));
AND2_X2 _cv_reg_U14  ( .A1(cv_d[86]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N89 ));
AND2_X2 _cv_reg_U12  ( .A1(cv_d[87]), .A2(_cv_reg_n250 ), .ZN(_cv_reg_N90 ));
AND2_X2 _cv_reg_U11  ( .A1(cv_d[88]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N91 ));
AND2_X2 _cv_reg_U10  ( .A1(cv_d[89]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N92 ));
AND2_X2 _cv_reg_U9  ( .A1(cv_d[90]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N93 ));
AND2_X2 _cv_reg_U8  ( .A1(cv_d[91]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N94 ));
AND2_X2 _cv_reg_U7  ( .A1(cv_d[92]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N95 ));
AND2_X2 _cv_reg_U6  ( .A1(cv_d[93]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N96 ));
AND2_X2 _cv_reg_U5  ( .A1(cv_d[94]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N97 ));
AND2_X2 _cv_reg_U4  ( .A1(cv_d[95]), .A2(_cv_reg_n240 ), .ZN(_cv_reg_N98 ));
DFF_X2 _cv_reg_q_reg_0_  ( .D(_cv_reg_N3 ), .CK(clk), .Q(cv_q[0]), .QN() );
DFF_X2 _cv_reg_q_reg_1_  ( .D(_cv_reg_N4 ), .CK(clk), .Q(cv_q[1]), .QN() );
DFF_X2 _cv_reg_q_reg_2_  ( .D(_cv_reg_N5 ), .CK(clk), .Q(cv_q[2]), .QN() );
DFF_X2 _cv_reg_q_reg_3_  ( .D(_cv_reg_N6 ), .CK(clk), .Q(cv_q[3]), .QN() );
DFF_X2 _cv_reg_q_reg_4_  ( .D(_cv_reg_N7 ), .CK(clk), .Q(cv_q[4]), .QN() );
DFF_X2 _cv_reg_q_reg_5_  ( .D(_cv_reg_N8 ), .CK(clk), .Q(cv_q[5]), .QN() );
DFF_X2 _cv_reg_q_reg_6_  ( .D(_cv_reg_N9 ), .CK(clk), .Q(cv_q[6]), .QN() );
DFF_X2 _cv_reg_q_reg_7_  ( .D(_cv_reg_N10 ), .CK(clk), .Q(cv_q[7]), .QN() );
DFF_X2 _cv_reg_q_reg_8_  ( .D(_cv_reg_N11 ), .CK(clk), .Q(cv_q[8]), .QN() );
DFF_X2 _cv_reg_q_reg_9_  ( .D(_cv_reg_N12 ), .CK(clk), .Q(cv_q[9]), .QN() );
DFF_X2 _cv_reg_q_reg_10_  ( .D(_cv_reg_N13 ), .CK(clk), .Q(cv_q[10]), .QN());
DFF_X2 _cv_reg_q_reg_11_  ( .D(_cv_reg_N14 ), .CK(clk), .Q(cv_q[11]), .QN());
DFF_X2 _cv_reg_q_reg_12_  ( .D(_cv_reg_N15 ), .CK(clk), .Q(cv_q[12]), .QN());
DFF_X2 _cv_reg_q_reg_13_  ( .D(_cv_reg_N16 ), .CK(clk), .Q(cv_q[13]), .QN());
DFF_X2 _cv_reg_q_reg_14_  ( .D(_cv_reg_N17 ), .CK(clk), .Q(cv_q[14]), .QN());
DFF_X2 _cv_reg_q_reg_15_  ( .D(_cv_reg_N18 ), .CK(clk), .Q(cv_q[15]), .QN());
DFF_X2 _cv_reg_q_reg_16_  ( .D(_cv_reg_N19 ), .CK(clk), .Q(cv_q[16]), .QN());
DFF_X2 _cv_reg_q_reg_17_  ( .D(_cv_reg_N20 ), .CK(clk), .Q(cv_q[17]), .QN());
DFF_X2 _cv_reg_q_reg_18_  ( .D(_cv_reg_N21 ), .CK(clk), .Q(cv_q[18]), .QN());
DFF_X2 _cv_reg_q_reg_19_  ( .D(_cv_reg_N22 ), .CK(clk), .Q(cv_q[19]), .QN());
DFF_X2 _cv_reg_q_reg_20_  ( .D(_cv_reg_N23 ), .CK(clk), .Q(cv_q[20]), .QN());
DFF_X2 _cv_reg_q_reg_21_  ( .D(_cv_reg_N24 ), .CK(clk), .Q(cv_q[21]), .QN());
DFF_X2 _cv_reg_q_reg_22_  ( .D(_cv_reg_N25 ), .CK(clk), .Q(cv_q[22]), .QN());
DFF_X2 _cv_reg_q_reg_23_  ( .D(_cv_reg_N26 ), .CK(clk), .Q(cv_q[23]), .QN());
DFF_X2 _cv_reg_q_reg_24_  ( .D(_cv_reg_N27 ), .CK(clk), .Q(cv_q[24]), .QN());
DFF_X2 _cv_reg_q_reg_25_  ( .D(_cv_reg_N28 ), .CK(clk), .Q(cv_q[25]), .QN());
DFF_X2 _cv_reg_q_reg_26_  ( .D(_cv_reg_N29 ), .CK(clk), .Q(cv_q[26]), .QN());
DFF_X2 _cv_reg_q_reg_27_  ( .D(_cv_reg_N30 ), .CK(clk), .Q(cv_q[27]), .QN());
DFF_X2 _cv_reg_q_reg_28_  ( .D(_cv_reg_N31 ), .CK(clk), .Q(cv_q[28]), .QN());
DFF_X2 _cv_reg_q_reg_29_  ( .D(_cv_reg_N32 ), .CK(clk), .Q(cv_q[29]), .QN());
DFF_X2 _cv_reg_q_reg_30_  ( .D(_cv_reg_N33 ), .CK(clk), .Q(cv_q[30]), .QN());
DFF_X2 _cv_reg_q_reg_31_  ( .D(_cv_reg_N34 ), .CK(clk), .Q(cv_q[31]), .QN());
DFF_X2 _cv_reg_q_reg_32_  ( .D(_cv_reg_N35 ), .CK(clk), .Q(cv_q[32]), .QN());
DFF_X2 _cv_reg_q_reg_33_  ( .D(_cv_reg_N36 ), .CK(clk), .Q(cv_q[33]), .QN());
DFF_X2 _cv_reg_q_reg_34_  ( .D(_cv_reg_N37 ), .CK(clk), .Q(cv_q[34]), .QN());
DFF_X2 _cv_reg_q_reg_35_  ( .D(_cv_reg_N38 ), .CK(clk), .Q(cv_q[35]), .QN());
DFF_X2 _cv_reg_q_reg_36_  ( .D(_cv_reg_N39 ), .CK(clk), .Q(cv_q[36]), .QN());
DFF_X2 _cv_reg_q_reg_37_  ( .D(_cv_reg_N40 ), .CK(clk), .Q(cv_q[37]), .QN());
DFF_X2 _cv_reg_q_reg_38_  ( .D(_cv_reg_N41 ), .CK(clk), .Q(cv_q[38]), .QN());
DFF_X2 _cv_reg_q_reg_39_  ( .D(_cv_reg_N42 ), .CK(clk), .Q(cv_q[39]), .QN());
DFF_X2 _cv_reg_q_reg_40_  ( .D(_cv_reg_N43 ), .CK(clk), .Q(cv_q[40]), .QN());
DFF_X2 _cv_reg_q_reg_41_  ( .D(_cv_reg_N44 ), .CK(clk), .Q(cv_q[41]), .QN());
DFF_X2 _cv_reg_q_reg_42_  ( .D(_cv_reg_N45 ), .CK(clk), .Q(cv_q[42]), .QN());
DFF_X2 _cv_reg_q_reg_43_  ( .D(_cv_reg_N46 ), .CK(clk), .Q(cv_q[43]), .QN());
DFF_X2 _cv_reg_q_reg_44_  ( .D(_cv_reg_N47 ), .CK(clk), .Q(cv_q[44]), .QN());
DFF_X2 _cv_reg_q_reg_45_  ( .D(_cv_reg_N48 ), .CK(clk), .Q(cv_q[45]), .QN());
DFF_X2 _cv_reg_q_reg_46_  ( .D(_cv_reg_N49 ), .CK(clk), .Q(cv_q[46]), .QN());
DFF_X2 _cv_reg_q_reg_47_  ( .D(_cv_reg_N50 ), .CK(clk), .Q(cv_q[47]), .QN());
DFF_X2 _cv_reg_q_reg_48_  ( .D(_cv_reg_N51 ), .CK(clk), .Q(cv_q[48]), .QN());
DFF_X2 _cv_reg_q_reg_49_  ( .D(_cv_reg_N52 ), .CK(clk), .Q(cv_q[49]), .QN());
DFF_X2 _cv_reg_q_reg_50_  ( .D(_cv_reg_N53 ), .CK(clk), .Q(cv_q[50]), .QN());
DFF_X2 _cv_reg_q_reg_51_  ( .D(_cv_reg_N54 ), .CK(clk), .Q(cv_q[51]), .QN());
DFF_X2 _cv_reg_q_reg_52_  ( .D(_cv_reg_N55 ), .CK(clk), .Q(cv_q[52]), .QN());
DFF_X2 _cv_reg_q_reg_53_  ( .D(_cv_reg_N56 ), .CK(clk), .Q(cv_q[53]), .QN());
DFF_X2 _cv_reg_q_reg_54_  ( .D(_cv_reg_N57 ), .CK(clk), .Q(cv_q[54]), .QN());
DFF_X2 _cv_reg_q_reg_55_  ( .D(_cv_reg_N58 ), .CK(clk), .Q(cv_q[55]), .QN());
DFF_X2 _cv_reg_q_reg_56_  ( .D(_cv_reg_N59 ), .CK(clk), .Q(cv_q[56]), .QN());
DFF_X2 _cv_reg_q_reg_57_  ( .D(_cv_reg_N60 ), .CK(clk), .Q(cv_q[57]), .QN());
DFF_X2 _cv_reg_q_reg_58_  ( .D(_cv_reg_N61 ), .CK(clk), .Q(cv_q[58]), .QN());
DFF_X2 _cv_reg_q_reg_59_  ( .D(_cv_reg_N62 ), .CK(clk), .Q(cv_q[59]), .QN());
DFF_X2 _cv_reg_q_reg_60_  ( .D(_cv_reg_N63 ), .CK(clk), .Q(cv_q[60]), .QN());
DFF_X2 _cv_reg_q_reg_61_  ( .D(_cv_reg_N64 ), .CK(clk), .Q(cv_q[61]), .QN());
DFF_X2 _cv_reg_q_reg_62_  ( .D(_cv_reg_N65 ), .CK(clk), .Q(cv_q[62]), .QN());
DFF_X2 _cv_reg_q_reg_63_  ( .D(_cv_reg_N66 ), .CK(clk), .Q(cv_q[63]), .QN());
DFF_X2 _cv_reg_q_reg_64_  ( .D(_cv_reg_N67 ), .CK(clk), .Q(cv_q[64]), .QN());
DFF_X2 _cv_reg_q_reg_65_  ( .D(_cv_reg_N68 ), .CK(clk), .Q(cv_q[65]), .QN());
DFF_X2 _cv_reg_q_reg_66_  ( .D(_cv_reg_N69 ), .CK(clk), .Q(cv_q[66]), .QN());
DFF_X2 _cv_reg_q_reg_67_  ( .D(_cv_reg_N70 ), .CK(clk), .Q(cv_q[67]), .QN());
DFF_X2 _cv_reg_q_reg_68_  ( .D(_cv_reg_N71 ), .CK(clk), .Q(cv_q[68]), .QN());
DFF_X2 _cv_reg_q_reg_69_  ( .D(_cv_reg_N72 ), .CK(clk), .Q(cv_q[69]), .QN());
DFF_X2 _cv_reg_q_reg_70_  ( .D(_cv_reg_N73 ), .CK(clk), .Q(cv_q[70]), .QN());
DFF_X2 _cv_reg_q_reg_71_  ( .D(_cv_reg_N74 ), .CK(clk), .Q(cv_q[71]), .QN());
DFF_X2 _cv_reg_q_reg_72_  ( .D(_cv_reg_N75 ), .CK(clk), .Q(cv_q[72]), .QN());
DFF_X2 _cv_reg_q_reg_73_  ( .D(_cv_reg_N76 ), .CK(clk), .Q(cv_q[73]), .QN());
DFF_X2 _cv_reg_q_reg_74_  ( .D(_cv_reg_N77 ), .CK(clk), .Q(cv_q[74]), .QN());
DFF_X2 _cv_reg_q_reg_75_  ( .D(_cv_reg_N78 ), .CK(clk), .Q(cv_q[75]), .QN());
DFF_X2 _cv_reg_q_reg_76_  ( .D(_cv_reg_N79 ), .CK(clk), .Q(cv_q[76]), .QN());
DFF_X2 _cv_reg_q_reg_77_  ( .D(_cv_reg_N80 ), .CK(clk), .Q(cv_q[77]), .QN());
DFF_X2 _cv_reg_q_reg_78_  ( .D(_cv_reg_N81 ), .CK(clk), .Q(cv_q[78]), .QN());
DFF_X2 _cv_reg_q_reg_79_  ( .D(_cv_reg_N82 ), .CK(clk), .Q(cv_q[79]), .QN());
DFF_X2 _cv_reg_q_reg_80_  ( .D(_cv_reg_N83 ), .CK(clk), .Q(cv_q[80]), .QN());
DFF_X2 _cv_reg_q_reg_81_  ( .D(_cv_reg_N84 ), .CK(clk), .Q(cv_q[81]), .QN());
DFF_X2 _cv_reg_q_reg_82_  ( .D(_cv_reg_N85 ), .CK(clk), .Q(cv_q[82]), .QN());
DFF_X2 _cv_reg_q_reg_83_  ( .D(_cv_reg_N86 ), .CK(clk), .Q(cv_q[83]), .QN());
DFF_X2 _cv_reg_q_reg_84_  ( .D(_cv_reg_N87 ), .CK(clk), .Q(cv_q[84]), .QN());
DFF_X2 _cv_reg_q_reg_85_  ( .D(_cv_reg_N88 ), .CK(clk), .Q(cv_q[85]), .QN());
DFF_X2 _cv_reg_q_reg_86_  ( .D(_cv_reg_N89 ), .CK(clk), .Q(cv_q[86]), .QN());
DFF_X2 _cv_reg_q_reg_87_  ( .D(_cv_reg_N90 ), .CK(clk), .Q(cv_q[87]), .QN());
DFF_X2 _cv_reg_q_reg_88_  ( .D(_cv_reg_N91 ), .CK(clk), .Q(cv_q[88]), .QN());
DFF_X2 _cv_reg_q_reg_89_  ( .D(_cv_reg_N92 ), .CK(clk), .Q(cv_q[89]), .QN());
DFF_X2 _cv_reg_q_reg_90_  ( .D(_cv_reg_N93 ), .CK(clk), .Q(cv_q[90]), .QN());
DFF_X2 _cv_reg_q_reg_91_  ( .D(_cv_reg_N94 ), .CK(clk), .Q(cv_q[91]), .QN());
DFF_X2 _cv_reg_q_reg_92_  ( .D(_cv_reg_N95 ), .CK(clk), .Q(cv_q[92]), .QN());
DFF_X2 _cv_reg_q_reg_93_  ( .D(_cv_reg_N96 ), .CK(clk), .Q(cv_q[93]), .QN());
DFF_X2 _cv_reg_q_reg_94_  ( .D(_cv_reg_N97 ), .CK(clk), .Q(cv_q[94]), .QN());
DFF_X2 _cv_reg_q_reg_95_  ( .D(_cv_reg_N98 ), .CK(clk), .Q(cv_q[95]), .QN());
DFF_X2 _cv_reg_q_reg_96_  ( .D(_cv_reg_N99 ), .CK(clk), .Q(cv_q[96]), .QN());
DFF_X2 _cv_reg_q_reg_97_  ( .D(_cv_reg_N100 ), .CK(clk), .Q(cv_q[97]), .QN());
DFF_X2 _cv_reg_q_reg_98_  ( .D(_cv_reg_N101 ), .CK(clk), .Q(cv_q[98]), .QN());
DFF_X2 _cv_reg_q_reg_99_  ( .D(_cv_reg_N102 ), .CK(clk), .Q(cv_q[99]), .QN());
DFF_X2 _cv_reg_q_reg_100_  ( .D(_cv_reg_N103 ), .CK(clk), .Q(cv_q[100]),.QN() );
DFF_X2 _cv_reg_q_reg_101_  ( .D(_cv_reg_N104 ), .CK(clk), .Q(cv_q[101]),.QN() );
DFF_X2 _cv_reg_q_reg_102_  ( .D(_cv_reg_N105 ), .CK(clk), .Q(cv_q[102]),.QN() );
DFF_X2 _cv_reg_q_reg_103_  ( .D(_cv_reg_N106 ), .CK(clk), .Q(cv_q[103]),.QN() );
DFF_X2 _cv_reg_q_reg_104_  ( .D(_cv_reg_N107 ), .CK(clk), .Q(cv_q[104]),.QN() );
DFF_X2 _cv_reg_q_reg_105_  ( .D(_cv_reg_N108 ), .CK(clk), .Q(cv_q[105]),.QN() );
DFF_X2 _cv_reg_q_reg_106_  ( .D(_cv_reg_N109 ), .CK(clk), .Q(cv_q[106]),.QN() );
DFF_X2 _cv_reg_q_reg_107_  ( .D(_cv_reg_N110 ), .CK(clk), .Q(cv_q[107]),.QN() );
DFF_X2 _cv_reg_q_reg_108_  ( .D(_cv_reg_N111 ), .CK(clk), .Q(cv_q[108]),.QN() );
DFF_X2 _cv_reg_q_reg_109_  ( .D(_cv_reg_N112 ), .CK(clk), .Q(cv_q[109]),.QN() );
DFF_X2 _cv_reg_q_reg_110_  ( .D(_cv_reg_N113 ), .CK(clk), .Q(cv_q[110]),.QN() );
DFF_X2 _cv_reg_q_reg_111_  ( .D(_cv_reg_N114 ), .CK(clk), .Q(cv_q[111]),.QN() );
DFF_X2 _cv_reg_q_reg_112_  ( .D(_cv_reg_N115 ), .CK(clk), .Q(cv_q[112]),.QN() );
DFF_X2 _cv_reg_q_reg_113_  ( .D(_cv_reg_N116 ), .CK(clk), .Q(cv_q[113]),.QN() );
DFF_X2 _cv_reg_q_reg_114_  ( .D(_cv_reg_N117 ), .CK(clk), .Q(cv_q[114]),.QN() );
DFF_X2 _cv_reg_q_reg_115_  ( .D(_cv_reg_N118 ), .CK(clk), .Q(cv_q[115]),.QN() );
DFF_X2 _cv_reg_q_reg_116_  ( .D(_cv_reg_N119 ), .CK(clk), .Q(cv_q[116]),.QN() );
DFF_X2 _cv_reg_q_reg_117_  ( .D(_cv_reg_N120 ), .CK(clk), .Q(cv_q[117]),.QN() );
DFF_X2 _cv_reg_q_reg_118_  ( .D(_cv_reg_N121 ), .CK(clk), .Q(cv_q[118]),.QN() );
DFF_X2 _cv_reg_q_reg_119_  ( .D(_cv_reg_N122 ), .CK(clk), .Q(cv_q[119]),.QN() );
DFF_X2 _cv_reg_q_reg_120_  ( .D(_cv_reg_N123 ), .CK(clk), .Q(cv_q[120]),.QN() );
DFF_X2 _cv_reg_q_reg_121_  ( .D(_cv_reg_N124 ), .CK(clk), .Q(cv_q[121]),.QN() );
DFF_X2 _cv_reg_q_reg_122_  ( .D(_cv_reg_N125 ), .CK(clk), .Q(cv_q[122]),.QN() );
DFF_X2 _cv_reg_q_reg_123_  ( .D(_cv_reg_N126 ), .CK(clk), .Q(cv_q[123]),.QN() );
DFF_X2 _cv_reg_q_reg_124_  ( .D(_cv_reg_N127 ), .CK(clk), .Q(cv_q[124]),.QN() );
DFF_X2 _cv_reg_q_reg_125_  ( .D(_cv_reg_N128 ), .CK(clk), .Q(cv_q[125]),.QN() );
DFF_X2 _cv_reg_q_reg_126_  ( .D(_cv_reg_N129 ), .CK(clk), .Q(cv_q[126]),.QN() );
DFF_X2 _cv_reg_q_reg_127_  ( .D(_cv_reg_N130 ), .CK(clk), .Q(cv_q[127]),.QN() );
DFF_X2 _cv_reg_q_reg_128_  ( .D(_cv_reg_N131 ), .CK(clk), .Q(cv_q[128]),.QN() );
DFF_X2 _cv_reg_q_reg_129_  ( .D(_cv_reg_N132 ), .CK(clk), .Q(cv_q[129]),.QN() );
DFF_X2 _cv_reg_q_reg_130_  ( .D(_cv_reg_N133 ), .CK(clk), .Q(cv_q[130]),.QN() );
DFF_X2 _cv_reg_q_reg_131_  ( .D(_cv_reg_N134 ), .CK(clk), .Q(cv_q[131]),.QN() );
DFF_X2 _cv_reg_q_reg_132_  ( .D(_cv_reg_N135 ), .CK(clk), .Q(cv_q[132]),.QN() );
DFF_X2 _cv_reg_q_reg_133_  ( .D(_cv_reg_N136 ), .CK(clk), .Q(cv_q[133]),.QN() );
DFF_X2 _cv_reg_q_reg_134_  ( .D(_cv_reg_N137 ), .CK(clk), .Q(cv_q[134]),.QN() );
DFF_X2 _cv_reg_q_reg_135_  ( .D(_cv_reg_N138 ), .CK(clk), .Q(cv_q[135]),.QN() );
DFF_X2 _cv_reg_q_reg_136_  ( .D(_cv_reg_N139 ), .CK(clk), .Q(cv_q[136]),.QN() );
DFF_X2 _cv_reg_q_reg_137_  ( .D(_cv_reg_N140 ), .CK(clk), .Q(cv_q[137]),.QN() );
DFF_X2 _cv_reg_q_reg_138_  ( .D(_cv_reg_N141 ), .CK(clk), .Q(cv_q[138]),.QN() );
DFF_X2 _cv_reg_q_reg_139_  ( .D(_cv_reg_N142 ), .CK(clk), .Q(cv_q[139]),.QN() );
DFF_X2 _cv_reg_q_reg_140_  ( .D(_cv_reg_N143 ), .CK(clk), .Q(cv_q[140]),.QN() );
DFF_X2 _cv_reg_q_reg_141_  ( .D(_cv_reg_N144 ), .CK(clk), .Q(cv_q[141]),.QN() );
DFF_X2 _cv_reg_q_reg_142_  ( .D(_cv_reg_N145 ), .CK(clk), .Q(cv_q[142]),.QN() );
DFF_X2 _cv_reg_q_reg_143_  ( .D(_cv_reg_N146 ), .CK(clk), .Q(cv_q[143]),.QN() );
DFF_X2 _cv_reg_q_reg_144_  ( .D(_cv_reg_N147 ), .CK(clk), .Q(cv_q[144]),.QN() );
DFF_X2 _cv_reg_q_reg_145_  ( .D(_cv_reg_N148 ), .CK(clk), .Q(cv_q[145]),.QN() );
DFF_X2 _cv_reg_q_reg_146_  ( .D(_cv_reg_N149 ), .CK(clk), .Q(cv_q[146]),.QN() );
DFF_X2 _cv_reg_q_reg_147_  ( .D(_cv_reg_N150 ), .CK(clk), .Q(cv_q[147]),.QN() );
DFF_X2 _cv_reg_q_reg_148_  ( .D(_cv_reg_N151 ), .CK(clk), .Q(cv_q[148]),.QN() );
DFF_X2 _cv_reg_q_reg_149_  ( .D(_cv_reg_N152 ), .CK(clk), .Q(cv_q[149]),.QN() );
DFF_X2 _cv_reg_q_reg_150_  ( .D(_cv_reg_N153 ), .CK(clk), .Q(cv_q[150]),.QN() );
DFF_X2 _cv_reg_q_reg_151_  ( .D(_cv_reg_N154 ), .CK(clk), .Q(cv_q[151]),.QN() );
DFF_X2 _cv_reg_q_reg_152_  ( .D(_cv_reg_N155 ), .CK(clk), .Q(cv_q[152]),.QN() );
DFF_X2 _cv_reg_q_reg_153_  ( .D(_cv_reg_N156 ), .CK(clk), .Q(cv_q[153]),.QN() );
DFF_X2 _cv_reg_q_reg_154_  ( .D(_cv_reg_N157 ), .CK(clk), .Q(cv_q[154]),.QN() );
DFF_X2 _cv_reg_q_reg_155_  ( .D(_cv_reg_N158 ), .CK(clk), .Q(cv_q[155]),.QN() );
DFF_X2 _cv_reg_q_reg_156_  ( .D(_cv_reg_N159 ), .CK(clk), .Q(cv_q[156]),.QN() );
DFF_X2 _cv_reg_q_reg_157_  ( .D(_cv_reg_N160 ), .CK(clk), .Q(cv_q[157]),.QN() );
DFF_X2 _cv_reg_q_reg_158_  ( .D(_cv_reg_N161 ), .CK(clk), .Q(cv_q[158]),.QN() );
DFF_X2 _cv_reg_q_reg_159_  ( .D(_cv_reg_N162 ), .CK(clk), .Q(cv_q[159]),.QN() );
AND2_X2 _rnd_reg_U178  ( .A1(rnd_d[159]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N162 ) );
AND2_X2 _rnd_reg_U177  ( .A1(rnd_d[158]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N161 ) );
AND2_X2 _rnd_reg_U176  ( .A1(rnd_d[157]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N160 ) );
AND2_X2 _rnd_reg_U175  ( .A1(rnd_d[156]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N159 ) );
AND2_X2 _rnd_reg_U174  ( .A1(rnd_d[154]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N157 ) );
AND2_X2 _rnd_reg_U173  ( .A1(rnd_d[153]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N156 ) );
AND2_X2 _rnd_reg_U172  ( .A1(rnd_d[152]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N155 ) );
AND2_X2 _rnd_reg_U171  ( .A1(rnd_d[151]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N154 ) );
AND2_X2 _rnd_reg_U170  ( .A1(rnd_d[149]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N152 ) );
AND2_X2 _rnd_reg_U169  ( .A1(rnd_d[148]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N151 ) );
AND2_X2 _rnd_reg_U168  ( .A1(rnd_d[147]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N150 ) );
AND2_X2 _rnd_reg_U167  ( .A1(rnd_d[146]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N149 ) );
AND2_X2 _rnd_reg_U166  ( .A1(rnd_d[145]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N148 ) );
AND2_X2 _rnd_reg_U165  ( .A1(rnd_d[144]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N147 ) );
AND2_X2 _rnd_reg_U164  ( .A1(rnd_d[143]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N146 ) );
AND2_X2 _rnd_reg_U163  ( .A1(rnd_d[142]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N145 ) );
AND2_X2 _rnd_reg_U162  ( .A1(rnd_d[141]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N144 ) );
AND2_X2 _rnd_reg_U161  ( .A1(rnd_d[140]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N143 ) );
AND2_X2 _rnd_reg_U160  ( .A1(rnd_d[139]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N142 ) );
AND2_X2 _rnd_reg_U159  ( .A1(rnd_d[138]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N141 ) );
AND2_X2 _rnd_reg_U158  ( .A1(rnd_d[137]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N140 ) );
AND2_X2 _rnd_reg_U157  ( .A1(rnd_d[136]), .A2(_rnd_reg_n250 ), .ZN(_rnd_reg_N139 ) );
AND2_X2 _rnd_reg_U156  ( .A1(rnd_d[135]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N138 ) );
AND2_X2 _rnd_reg_U155  ( .A1(rnd_d[134]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N137 ) );
AND2_X2 _rnd_reg_U154  ( .A1(rnd_d[133]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N136 ) );
AND2_X2 _rnd_reg_U153  ( .A1(rnd_d[132]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N135 ) );
AND2_X2 _rnd_reg_U152  ( .A1(rnd_d[131]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N134 ) );
AND2_X2 _rnd_reg_U151  ( .A1(rnd_d[130]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N133 ) );
AND2_X2 _rnd_reg_U150  ( .A1(rnd_d[129]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N132 ) );
AND2_X2 _rnd_reg_U149  ( .A1(rnd_d[128]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N131 ) );
AND2_X2 _rnd_reg_U148  ( .A1(rnd_d[116]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N119 ) );
AND2_X2 _rnd_reg_U147  ( .A1(rnd_d[115]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N118 ) );
AND2_X2 _rnd_reg_U146  ( .A1(rnd_d[114]), .A2(_rnd_reg_n240 ), .ZN(_rnd_reg_N117 ) );
AND2_X2 _rnd_reg_U145  ( .A1(rnd_d[113]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N116 ) );
AND2_X2 _rnd_reg_U144  ( .A1(rnd_d[112]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N115 ) );
AND2_X2 _rnd_reg_U143  ( .A1(rnd_d[111]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N114 ) );
AND2_X2 _rnd_reg_U142  ( .A1(rnd_d[110]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N113 ) );
AND2_X2 _rnd_reg_U141  ( .A1(rnd_d[109]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N112 ) );
AND2_X2 _rnd_reg_U140  ( .A1(rnd_d[108]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N111 ) );
AND2_X2 _rnd_reg_U129  ( .A1(rnd_d[107]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N110 ) );
AND2_X2 _rnd_reg_U127  ( .A1(rnd_d[106]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N109 ) );
AND2_X2 _rnd_reg_U126  ( .A1(rnd_d[105]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N108 ) );
AND2_X2 _rnd_reg_U125  ( .A1(rnd_d[104]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N107 ) );
AND2_X2 _rnd_reg_U124  ( .A1(rnd_d[103]), .A2(_rnd_reg_n230 ), .ZN(_rnd_reg_N106 ) );
AND2_X2 _rnd_reg_U123  ( .A1(rnd_d[102]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N105 ) );
AND2_X2 _rnd_reg_U122  ( .A1(rnd_d[101]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N104 ) );
AND2_X2 _rnd_reg_U121  ( .A1(rnd_d[100]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N103 ) );
AND2_X2 _rnd_reg_U120  ( .A1(rnd_d[99]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N102 ) );
AND2_X2 _rnd_reg_U119  ( .A1(rnd_d[98]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N101 ) );
AND2_X2 _rnd_reg_U118  ( .A1(rnd_d[97]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N100 ) );
AND2_X2 _rnd_reg_U117  ( .A1(rnd_d[96]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N99 ) );
AND2_X2 _rnd_reg_U116  ( .A1(rnd_d[83]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N86 ) );
AND2_X2 _rnd_reg_U115  ( .A1(rnd_d[82]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N85 ) );
AND2_X2 _rnd_reg_U114  ( .A1(rnd_d[81]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N84 ) );
AND2_X2 _rnd_reg_U113  ( .A1(rnd_d[80]), .A2(_rnd_reg_n220 ), .ZN(_rnd_reg_N83 ) );
AND2_X2 _rnd_reg_U112  ( .A1(rnd_d[79]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N82 ) );
AND2_X2 _rnd_reg_U111  ( .A1(rnd_d[78]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N81 ) );
AND2_X2 _rnd_reg_U110  ( .A1(rnd_d[77]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N80 ) );
AND2_X2 _rnd_reg_U109  ( .A1(rnd_d[76]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N79 ) );
AND2_X2 _rnd_reg_U108  ( .A1(rnd_d[75]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N78 ) );
AND2_X2 _rnd_reg_U107  ( .A1(rnd_d[74]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N77 ) );
AND2_X2 _rnd_reg_U106  ( .A1(rnd_d[73]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N76 ) );
AND2_X2 _rnd_reg_U105  ( .A1(rnd_d[72]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N75 ) );
AND2_X2 _rnd_reg_U104  ( .A1(rnd_d[71]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N74 ) );
AND2_X2 _rnd_reg_U103  ( .A1(rnd_d[70]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N73 ) );
AND2_X2 _rnd_reg_U102  ( .A1(rnd_d[69]), .A2(_rnd_reg_n210 ), .ZN(_rnd_reg_N72 ) );
AND2_X2 _rnd_reg_U101  ( .A1(rnd_d[68]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N71 ) );
AND2_X2 _rnd_reg_U100  ( .A1(rnd_d[67]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N70 ) );
AND2_X2 _rnd_reg_U99  ( .A1(rnd_d[66]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N69 ) );
AND2_X2 _rnd_reg_U98  ( .A1(rnd_d[65]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N68 ) );
AND2_X2 _rnd_reg_U97  ( .A1(rnd_d[64]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N67 ) );
AND2_X2 _rnd_reg_U96  ( .A1(rnd_d[51]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N54 ) );
AND2_X2 _rnd_reg_U95  ( .A1(rnd_d[50]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N53 ) );
AND2_X2 _rnd_reg_U94  ( .A1(rnd_d[49]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N52 ) );
AND2_X2 _rnd_reg_U93  ( .A1(rnd_d[48]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N51 ) );
AND2_X2 _rnd_reg_U92  ( .A1(rnd_d[47]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N50 ) );
AND2_X2 _rnd_reg_U91  ( .A1(rnd_d[46]), .A2(_rnd_reg_n200 ), .ZN(_rnd_reg_N49 ) );
AND2_X2 _rnd_reg_U90  ( .A1(rnd_d[45]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N48 ) );
AND2_X2 _rnd_reg_U89  ( .A1(rnd_d[44]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N47 ) );
AND2_X2 _rnd_reg_U88  ( .A1(rnd_d[43]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N46 ) );
AND2_X2 _rnd_reg_U79  ( .A1(rnd_d[42]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N45 ) );
AND2_X2 _rnd_reg_U73  ( .A1(rnd_d[41]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N44 ) );
AND2_X2 _rnd_reg_U72  ( .A1(rnd_d[40]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N43 ) );
AND2_X2 _rnd_reg_U71  ( .A1(rnd_d[39]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N42 ) );
AND2_X2 _rnd_reg_U70  ( .A1(rnd_d[38]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N41 ) );
AND2_X2 _rnd_reg_U69  ( .A1(rnd_d[37]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N40 ) );
AND2_X2 _rnd_reg_U68  ( .A1(rnd_d[36]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N39 ) );
AND2_X2 _rnd_reg_U67  ( .A1(rnd_d[35]), .A2(_rnd_reg_n190 ), .ZN(_rnd_reg_N38 ) );
AND2_X2 _rnd_reg_U66  ( .A1(rnd_d[34]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N37 ) );
AND2_X2 _rnd_reg_U65  ( .A1(rnd_d[33]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N36 ) );
AND2_X2 _rnd_reg_U64  ( .A1(rnd_d[32]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N35 ) );
AND2_X2 _rnd_reg_U63  ( .A1(rnd_d[18]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N21 ) );
AND2_X2 _rnd_reg_U62  ( .A1(rnd_d[17]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N20 ) );
AND2_X2 _rnd_reg_U61  ( .A1(rnd_d[16]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N19 ) );
AND2_X2 _rnd_reg_U60  ( .A1(rnd_d[15]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N18 ) );
AND2_X2 _rnd_reg_U59  ( .A1(rnd_d[14]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N17 ) );
AND2_X2 _rnd_reg_U58  ( .A1(rnd_d[13]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N16 ) );
AND2_X2 _rnd_reg_U57  ( .A1(rnd_d[12]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N15 ) );
AND2_X2 _rnd_reg_U56  ( .A1(rnd_d[11]), .A2(_rnd_reg_n180 ), .ZN(_rnd_reg_N14 ) );
AND2_X2 _rnd_reg_U55  ( .A1(rnd_d[10]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N13 ) );
AND2_X2 _rnd_reg_U54  ( .A1(rnd_d[9]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N12 ) );
AND2_X2 _rnd_reg_U53  ( .A1(rnd_d[8]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N11 ) );
AND2_X2 _rnd_reg_U52  ( .A1(rnd_d[7]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N10 ) );
AND2_X2 _rnd_reg_U46  ( .A1(rnd_d[6]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N9 ) );
AND2_X2 _rnd_reg_U38  ( .A1(rnd_d[5]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N8 ) );
AND2_X2 _rnd_reg_U37  ( .A1(rnd_d[4]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N7 ) );
AND2_X2 _rnd_reg_U36  ( .A1(rnd_d[3]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N6 ) );
AND2_X2 _rnd_reg_U35  ( .A1(rnd_d[2]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N5 ) );
AND2_X2 _rnd_reg_U34  ( .A1(rnd_d[1]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N4 ) );
AND2_X2 _rnd_reg_U33  ( .A1(rnd_d[0]), .A2(_rnd_reg_n170 ), .ZN(_rnd_reg_N3 ) );
INV_X4 _rnd_reg_U32  ( .A(_rnd_reg_n190 ), .ZN(_rnd_reg_n320 ) );
INV_X4 _rnd_reg_U31  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n310 ) );
INV_X4 _rnd_reg_U30  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n220 ) );
INV_X4 _rnd_reg_U29  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n210 ) );
INV_X4 _rnd_reg_U28  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n200 ) );
INV_X4 _rnd_reg_U27  ( .A(n7117), .ZN(_rnd_reg_n190 ) );
INV_X4 _rnd_reg_U26  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n180 ) );
INV_X4 _rnd_reg_U25  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n170 ) );
INV_X4 _rnd_reg_U24  ( .A(n7117), .ZN(_rnd_reg_n260 ) );
INV_X4 _rnd_reg_U23  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n250 ) );
INV_X4 _rnd_reg_U22  ( .A(n7117), .ZN(_rnd_reg_n240 ) );
INV_X4 _rnd_reg_U21  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n300 ) );
INV_X4 _rnd_reg_U20  ( .A(n7117), .ZN(_rnd_reg_n230 ) );
INV_X4 _rnd_reg_U19  ( .A(n7117), .ZN(_rnd_reg_n270 ) );
INV_X4 _rnd_reg_U18  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n280 ) );
INV_X4 _rnd_reg_U17  ( .A(_rnd_reg_n320 ), .ZN(_rnd_reg_n290 ) );
AND2_X4 _rnd_reg_U13  ( .A1(rnd_d[155]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N158 ) );
AND2_X4 _rnd_reg_U3  ( .A1(rnd_d[150]), .A2(_rnd_reg_n260 ), .ZN(_rnd_reg_N153 ) );
DFF_X2 _rnd_reg_q_reg_156_  ( .D(_rnd_reg_N159 ), .CK(clk), .Q(rnd_q[156]),.QN() );
DFF_X2 _rnd_reg_q_reg_155_  ( .D(_rnd_reg_N158 ), .CK(clk), .Q(rnd_q[155]),.QN() );
DFF_X2 _rnd_reg_q_reg_158_  ( .D(_rnd_reg_N161 ), .CK(clk), .Q(rnd_q[158]),.QN() );
DFF_X2 _rnd_reg_q_reg_157_  ( .D(_rnd_reg_N160 ), .CK(clk), .Q(rnd_q[157]),.QN() );
DFF_X2 _rnd_reg_q_reg_159_  ( .D(_rnd_reg_N162 ), .CK(clk), .Q(rnd_q[159]),.QN() );
DFF_X2 _rnd_reg_q_reg_150_  ( .D(_rnd_reg_N153 ), .CK(clk), .Q(rnd_q[150]),.QN() );
DFF_X2 _rnd_reg_q_reg_154_  ( .D(_rnd_reg_N157 ), .CK(clk), .Q(rnd_q[154]),.QN() );
DFF_X2 _rnd_reg_q_reg_153_  ( .D(_rnd_reg_N156 ), .CK(clk), .Q(rnd_q[153]),.QN() );
DFF_X2 _rnd_reg_q_reg_151_  ( .D(_rnd_reg_N154 ), .CK(clk), .Q(rnd_q[151]),.QN() );
AND2_X2 _rnd_reg_U139  ( .A1(rnd_d[117]), .A2(_rnd_reg_n310 ), .ZN(_rnd_reg_N120 ) );
AND2_X2 _rnd_reg_U138  ( .A1(rnd_d[118]), .A2(_rnd_reg_n310 ), .ZN(_rnd_reg_N121 ) );
AND2_X2 _rnd_reg_U137  ( .A1(rnd_d[119]), .A2(_rnd_reg_n310 ), .ZN(_rnd_reg_N122 ) );
AND2_X2 _rnd_reg_U136  ( .A1(rnd_d[120]), .A2(_rnd_reg_n310 ), .ZN(_rnd_reg_N123 ) );
AND2_X2 _rnd_reg_U135  ( .A1(rnd_d[121]), .A2(_rnd_reg_n310 ), .ZN(_rnd_reg_N124 ) );
AND2_X2 _rnd_reg_U134  ( .A1(rnd_d[122]), .A2(_rnd_reg_n310 ), .ZN(_rnd_reg_N125 ) );
AND2_X2 _rnd_reg_U133  ( .A1(rnd_d[123]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N126 ) );
AND2_X2 _rnd_reg_U132  ( .A1(rnd_d[124]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N127 ) );
AND2_X2 _rnd_reg_U131  ( .A1(rnd_d[125]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N128 ) );
AND2_X2 _rnd_reg_U130  ( .A1(rnd_d[126]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N129 ) );
AND2_X2 _rnd_reg_U128  ( .A1(rnd_d[127]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N130 ) );
AND2_X2 _rnd_reg_U87  ( .A1(rnd_d[19]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N22 ) );
AND2_X2 _rnd_reg_U86  ( .A1(rnd_d[20]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N23 ) );
AND2_X2 _rnd_reg_U85  ( .A1(rnd_d[21]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N24 ) );
AND2_X2 _rnd_reg_U84  ( .A1(rnd_d[22]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N25 ) );
AND2_X2 _rnd_reg_U83  ( .A1(rnd_d[23]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N26 ) );
AND2_X2 _rnd_reg_U82  ( .A1(rnd_d[24]), .A2(_rnd_reg_n300 ), .ZN(_rnd_reg_N27 ) );
AND2_X2 _rnd_reg_U81  ( .A1(rnd_d[25]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N28 ) );
AND2_X2 _rnd_reg_U80  ( .A1(rnd_d[26]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N29 ) );
AND2_X2 _rnd_reg_U78  ( .A1(rnd_d[27]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N30 ) );
AND2_X2 _rnd_reg_U77  ( .A1(rnd_d[28]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N31 ) );
AND2_X2 _rnd_reg_U76  ( .A1(rnd_d[29]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N32 ) );
AND2_X2 _rnd_reg_U75  ( .A1(rnd_d[30]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N33 ) );
AND2_X2 _rnd_reg_U74  ( .A1(rnd_d[31]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N34 ) );
AND2_X2 _rnd_reg_U51  ( .A1(rnd_d[52]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N55 ) );
AND2_X2 _rnd_reg_U50  ( .A1(rnd_d[53]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N56 ) );
AND2_X2 _rnd_reg_U49  ( .A1(rnd_d[54]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N57 ) );
AND2_X2 _rnd_reg_U48  ( .A1(rnd_d[55]), .A2(_rnd_reg_n290 ), .ZN(_rnd_reg_N58 ) );
AND2_X2 _rnd_reg_U47  ( .A1(rnd_d[56]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N59 ) );
AND2_X2 _rnd_reg_U45  ( .A1(rnd_d[57]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N60 ) );
AND2_X2 _rnd_reg_U44  ( .A1(rnd_d[58]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N61 ) );
AND2_X2 _rnd_reg_U43  ( .A1(rnd_d[59]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N62 ) );
AND2_X2 _rnd_reg_U42  ( .A1(rnd_d[60]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N63 ) );
AND2_X2 _rnd_reg_U41  ( .A1(rnd_d[61]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N64 ) );
AND2_X2 _rnd_reg_U40  ( .A1(rnd_d[62]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N65 ) );
AND2_X2 _rnd_reg_U39  ( .A1(rnd_d[63]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N66 ) );
AND2_X2 _rnd_reg_U16  ( .A1(rnd_d[84]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N87 ) );
AND2_X2 _rnd_reg_U15  ( .A1(rnd_d[85]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N88 ) );
AND2_X2 _rnd_reg_U14  ( .A1(rnd_d[86]), .A2(_rnd_reg_n280 ), .ZN(_rnd_reg_N89 ) );
AND2_X2 _rnd_reg_U12  ( .A1(rnd_d[87]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N90 ) );
AND2_X2 _rnd_reg_U11  ( .A1(rnd_d[88]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N91 ) );
AND2_X2 _rnd_reg_U10  ( .A1(rnd_d[89]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N92 ) );
AND2_X2 _rnd_reg_U9  ( .A1(rnd_d[90]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N93 ) );
AND2_X2 _rnd_reg_U8  ( .A1(rnd_d[91]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N94 ) );
AND2_X2 _rnd_reg_U7  ( .A1(rnd_d[92]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N95 ) );
AND2_X2 _rnd_reg_U6  ( .A1(rnd_d[93]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N96 ) );
AND2_X2 _rnd_reg_U5  ( .A1(rnd_d[94]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N97 ) );
AND2_X2 _rnd_reg_U4  ( .A1(rnd_d[95]), .A2(_rnd_reg_n270 ), .ZN(_rnd_reg_N98 ) );
DFF_X2 _rnd_reg_q_reg_0_  ( .D(_rnd_reg_N3 ), .CK(clk), .Q(rnd_q[0]), .QN());
DFF_X2 _rnd_reg_q_reg_1_  ( .D(_rnd_reg_N4 ), .CK(clk), .Q(rnd_q[1]), .QN());
DFF_X2 _rnd_reg_q_reg_2_  ( .D(_rnd_reg_N5 ), .CK(clk), .Q(rnd_q[2]), .QN());
DFF_X2 _rnd_reg_q_reg_3_  ( .D(_rnd_reg_N6 ), .CK(clk), .Q(rnd_q[3]), .QN());
DFF_X2 _rnd_reg_q_reg_4_  ( .D(_rnd_reg_N7 ), .CK(clk), .Q(rnd_q[4]), .QN());
DFF_X2 _rnd_reg_q_reg_5_  ( .D(_rnd_reg_N8 ), .CK(clk), .Q(rnd_q[5]), .QN());
DFF_X2 _rnd_reg_q_reg_6_  ( .D(_rnd_reg_N9 ), .CK(clk), .Q(rnd_q[6]), .QN());
DFF_X2 _rnd_reg_q_reg_7_  ( .D(_rnd_reg_N10 ), .CK(clk), .Q(rnd_q[7]), .QN());
DFF_X2 _rnd_reg_q_reg_8_  ( .D(_rnd_reg_N11 ), .CK(clk), .Q(rnd_q[8]), .QN());
DFF_X2 _rnd_reg_q_reg_9_  ( .D(_rnd_reg_N12 ), .CK(clk), .Q(rnd_q[9]), .QN());
DFF_X2 _rnd_reg_q_reg_10_  ( .D(_rnd_reg_N13 ), .CK(clk), .Q(rnd_q[10]),.QN() );
DFF_X2 _rnd_reg_q_reg_11_  ( .D(_rnd_reg_N14 ), .CK(clk), .Q(rnd_q[11]),.QN() );
DFF_X2 _rnd_reg_q_reg_12_  ( .D(_rnd_reg_N15 ), .CK(clk), .Q(rnd_q[12]),.QN() );
DFF_X2 _rnd_reg_q_reg_13_  ( .D(_rnd_reg_N16 ), .CK(clk), .Q(rnd_q[13]),.QN() );
DFF_X2 _rnd_reg_q_reg_14_  ( .D(_rnd_reg_N17 ), .CK(clk), .Q(rnd_q[14]),.QN() );
DFF_X2 _rnd_reg_q_reg_15_  ( .D(_rnd_reg_N18 ), .CK(clk), .Q(rnd_q[15]),.QN() );
DFF_X2 _rnd_reg_q_reg_16_  ( .D(_rnd_reg_N19 ), .CK(clk), .Q(rnd_q[16]),.QN() );
DFF_X2 _rnd_reg_q_reg_17_  ( .D(_rnd_reg_N20 ), .CK(clk), .Q(rnd_q[17]),.QN() );
DFF_X2 _rnd_reg_q_reg_18_  ( .D(_rnd_reg_N21 ), .CK(clk), .Q(rnd_q[18]),.QN() );
DFF_X2 _rnd_reg_q_reg_19_  ( .D(_rnd_reg_N22 ), .CK(clk), .Q(rnd_q[19]),.QN() );
DFF_X2 _rnd_reg_q_reg_20_  ( .D(_rnd_reg_N23 ), .CK(clk), .Q(rnd_q[20]),.QN() );
DFF_X2 _rnd_reg_q_reg_21_  ( .D(_rnd_reg_N24 ), .CK(clk), .Q(rnd_q[21]),.QN() );
DFF_X2 _rnd_reg_q_reg_22_  ( .D(_rnd_reg_N25 ), .CK(clk), .Q(rnd_q[22]),.QN() );
DFF_X2 _rnd_reg_q_reg_23_  ( .D(_rnd_reg_N26 ), .CK(clk), .Q(rnd_q[23]),.QN() );
DFF_X2 _rnd_reg_q_reg_24_  ( .D(_rnd_reg_N27 ), .CK(clk), .Q(rnd_q[24]),.QN() );
DFF_X2 _rnd_reg_q_reg_25_  ( .D(_rnd_reg_N28 ), .CK(clk), .Q(rnd_q[25]),.QN() );
DFF_X2 _rnd_reg_q_reg_26_  ( .D(_rnd_reg_N29 ), .CK(clk), .Q(rnd_q[26]),.QN() );
DFF_X2 _rnd_reg_q_reg_27_  ( .D(_rnd_reg_N30 ), .CK(clk), .Q(rnd_q[27]),.QN() );
DFF_X2 _rnd_reg_q_reg_28_  ( .D(_rnd_reg_N31 ), .CK(clk), .Q(rnd_q[28]),.QN() );
DFF_X2 _rnd_reg_q_reg_29_  ( .D(_rnd_reg_N32 ), .CK(clk), .Q(rnd_q[29]),.QN() );
DFF_X2 _rnd_reg_q_reg_30_  ( .D(_rnd_reg_N33 ), .CK(clk), .Q(rnd_q[30]),.QN() );
DFF_X2 _rnd_reg_q_reg_31_  ( .D(_rnd_reg_N34 ), .CK(clk), .Q(rnd_q[31]),.QN() );
DFF_X2 _rnd_reg_q_reg_32_  ( .D(_rnd_reg_N35 ), .CK(clk), .Q(rnd_q[32]),.QN() );
DFF_X2 _rnd_reg_q_reg_33_  ( .D(_rnd_reg_N36 ), .CK(clk), .Q(rnd_q[33]),.QN() );
DFF_X2 _rnd_reg_q_reg_34_  ( .D(_rnd_reg_N37 ), .CK(clk), .Q(rnd_q[34]),.QN() );
DFF_X2 _rnd_reg_q_reg_35_  ( .D(_rnd_reg_N38 ), .CK(clk), .Q(rnd_q[35]),.QN() );
DFF_X2 _rnd_reg_q_reg_36_  ( .D(_rnd_reg_N39 ), .CK(clk), .Q(rnd_q[36]),.QN() );
DFF_X2 _rnd_reg_q_reg_37_  ( .D(_rnd_reg_N40 ), .CK(clk), .Q(rnd_q[37]),.QN() );
DFF_X2 _rnd_reg_q_reg_38_  ( .D(_rnd_reg_N41 ), .CK(clk), .Q(rnd_q[38]),.QN() );
DFF_X2 _rnd_reg_q_reg_39_  ( .D(_rnd_reg_N42 ), .CK(clk), .Q(rnd_q[39]),.QN() );
DFF_X2 _rnd_reg_q_reg_40_  ( .D(_rnd_reg_N43 ), .CK(clk), .Q(rnd_q[40]),.QN() );
DFF_X2 _rnd_reg_q_reg_41_  ( .D(_rnd_reg_N44 ), .CK(clk), .Q(rnd_q[41]),.QN() );
DFF_X2 _rnd_reg_q_reg_42_  ( .D(_rnd_reg_N45 ), .CK(clk), .Q(rnd_q[42]),.QN() );
DFF_X2 _rnd_reg_q_reg_43_  ( .D(_rnd_reg_N46 ), .CK(clk), .Q(rnd_q[43]),.QN() );
DFF_X2 _rnd_reg_q_reg_44_  ( .D(_rnd_reg_N47 ), .CK(clk), .Q(rnd_q[44]),.QN() );
DFF_X2 _rnd_reg_q_reg_45_  ( .D(_rnd_reg_N48 ), .CK(clk), .Q(rnd_q[45]),.QN() );
DFF_X2 _rnd_reg_q_reg_46_  ( .D(_rnd_reg_N49 ), .CK(clk), .Q(rnd_q[46]),.QN() );
DFF_X2 _rnd_reg_q_reg_47_  ( .D(_rnd_reg_N50 ), .CK(clk), .Q(rnd_q[47]),.QN() );
DFF_X2 _rnd_reg_q_reg_48_  ( .D(_rnd_reg_N51 ), .CK(clk), .Q(rnd_q[48]),.QN() );
DFF_X2 _rnd_reg_q_reg_49_  ( .D(_rnd_reg_N52 ), .CK(clk), .Q(rnd_q[49]),.QN() );
DFF_X2 _rnd_reg_q_reg_50_  ( .D(_rnd_reg_N53 ), .CK(clk), .Q(rnd_q[50]),.QN() );
DFF_X2 _rnd_reg_q_reg_51_  ( .D(_rnd_reg_N54 ), .CK(clk), .Q(rnd_q[51]),.QN() );
DFF_X2 _rnd_reg_q_reg_52_  ( .D(_rnd_reg_N55 ), .CK(clk), .Q(rnd_q[52]),.QN() );
DFF_X2 _rnd_reg_q_reg_53_  ( .D(_rnd_reg_N56 ), .CK(clk), .Q(rnd_q[53]),.QN() );
DFF_X2 _rnd_reg_q_reg_54_  ( .D(_rnd_reg_N57 ), .CK(clk), .Q(rnd_q[54]),.QN() );
DFF_X2 _rnd_reg_q_reg_55_  ( .D(_rnd_reg_N58 ), .CK(clk), .Q(rnd_q[55]),.QN() );
DFF_X2 _rnd_reg_q_reg_56_  ( .D(_rnd_reg_N59 ), .CK(clk), .Q(rnd_q[56]),.QN() );
DFF_X2 _rnd_reg_q_reg_57_  ( .D(_rnd_reg_N60 ), .CK(clk), .Q(rnd_q[57]),.QN() );
DFF_X2 _rnd_reg_q_reg_58_  ( .D(_rnd_reg_N61 ), .CK(clk), .Q(rnd_q[58]),.QN() );
DFF_X2 _rnd_reg_q_reg_59_  ( .D(_rnd_reg_N62 ), .CK(clk), .Q(rnd_q[59]),.QN() );
DFF_X2 _rnd_reg_q_reg_60_  ( .D(_rnd_reg_N63 ), .CK(clk), .Q(rnd_q[60]),.QN() );
DFF_X2 _rnd_reg_q_reg_61_  ( .D(_rnd_reg_N64 ), .CK(clk), .Q(rnd_q[61]),.QN() );
DFF_X2 _rnd_reg_q_reg_62_  ( .D(_rnd_reg_N65 ), .CK(clk), .Q(rnd_q[62]),.QN() );
DFF_X2 _rnd_reg_q_reg_63_  ( .D(_rnd_reg_N66 ), .CK(clk), .Q(rnd_q[63]),.QN() );
DFF_X2 _rnd_reg_q_reg_64_  ( .D(_rnd_reg_N67 ), .CK(clk), .Q(rnd_q[64]),.QN() );
DFF_X2 _rnd_reg_q_reg_65_  ( .D(_rnd_reg_N68 ), .CK(clk), .Q(rnd_q[65]),.QN() );
DFF_X2 _rnd_reg_q_reg_66_  ( .D(_rnd_reg_N69 ), .CK(clk), .Q(rnd_q[66]),.QN() );
DFF_X2 _rnd_reg_q_reg_67_  ( .D(_rnd_reg_N70 ), .CK(clk), .Q(rnd_q[67]),.QN() );
DFF_X2 _rnd_reg_q_reg_68_  ( .D(_rnd_reg_N71 ), .CK(clk), .Q(rnd_q[68]),.QN() );
DFF_X2 _rnd_reg_q_reg_69_  ( .D(_rnd_reg_N72 ), .CK(clk), .Q(rnd_q[69]),.QN() );
DFF_X2 _rnd_reg_q_reg_70_  ( .D(_rnd_reg_N73 ), .CK(clk), .Q(rnd_q[70]),.QN() );
DFF_X2 _rnd_reg_q_reg_71_  ( .D(_rnd_reg_N74 ), .CK(clk), .Q(rnd_q[71]),.QN() );
DFF_X2 _rnd_reg_q_reg_72_  ( .D(_rnd_reg_N75 ), .CK(clk), .Q(rnd_q[72]),.QN() );
DFF_X2 _rnd_reg_q_reg_73_  ( .D(_rnd_reg_N76 ), .CK(clk), .Q(rnd_q[73]),.QN() );
DFF_X2 _rnd_reg_q_reg_74_  ( .D(_rnd_reg_N77 ), .CK(clk), .Q(rnd_q[74]),.QN() );
DFF_X2 _rnd_reg_q_reg_75_  ( .D(_rnd_reg_N78 ), .CK(clk), .Q(rnd_q[75]),.QN() );
DFF_X2 _rnd_reg_q_reg_76_  ( .D(_rnd_reg_N79 ), .CK(clk), .Q(rnd_q[76]),.QN() );
DFF_X2 _rnd_reg_q_reg_77_  ( .D(_rnd_reg_N80 ), .CK(clk), .Q(rnd_q[77]),.QN() );
DFF_X2 _rnd_reg_q_reg_78_  ( .D(_rnd_reg_N81 ), .CK(clk), .Q(rnd_q[78]),.QN() );
DFF_X2 _rnd_reg_q_reg_79_  ( .D(_rnd_reg_N82 ), .CK(clk), .Q(rnd_q[79]),.QN() );
DFF_X2 _rnd_reg_q_reg_80_  ( .D(_rnd_reg_N83 ), .CK(clk), .Q(rnd_q[80]),.QN() );
DFF_X2 _rnd_reg_q_reg_81_  ( .D(_rnd_reg_N84 ), .CK(clk), .Q(rnd_q[81]),.QN() );
DFF_X2 _rnd_reg_q_reg_82_  ( .D(_rnd_reg_N85 ), .CK(clk), .Q(rnd_q[82]),.QN() );
DFF_X2 _rnd_reg_q_reg_83_  ( .D(_rnd_reg_N86 ), .CK(clk), .Q(rnd_q[83]),.QN() );
DFF_X2 _rnd_reg_q_reg_84_  ( .D(_rnd_reg_N87 ), .CK(clk), .Q(rnd_q[84]),.QN() );
DFF_X2 _rnd_reg_q_reg_85_  ( .D(_rnd_reg_N88 ), .CK(clk), .Q(rnd_q[85]),.QN() );
DFF_X2 _rnd_reg_q_reg_86_  ( .D(_rnd_reg_N89 ), .CK(clk), .Q(rnd_q[86]),.QN() );
DFF_X2 _rnd_reg_q_reg_87_  ( .D(_rnd_reg_N90 ), .CK(clk), .Q(rnd_q[87]),.QN() );
DFF_X2 _rnd_reg_q_reg_88_  ( .D(_rnd_reg_N91 ), .CK(clk), .Q(rnd_q[88]),.QN() );
DFF_X2 _rnd_reg_q_reg_89_  ( .D(_rnd_reg_N92 ), .CK(clk), .Q(rnd_q[89]),.QN() );
DFF_X2 _rnd_reg_q_reg_90_  ( .D(_rnd_reg_N93 ), .CK(clk), .Q(rnd_q[90]),.QN() );
DFF_X2 _rnd_reg_q_reg_91_  ( .D(_rnd_reg_N94 ), .CK(clk), .Q(rnd_q[91]),.QN() );
DFF_X2 _rnd_reg_q_reg_92_  ( .D(_rnd_reg_N95 ), .CK(clk), .Q(rnd_q[92]),.QN() );
DFF_X2 _rnd_reg_q_reg_93_  ( .D(_rnd_reg_N96 ), .CK(clk), .Q(rnd_q[93]),.QN() );
DFF_X2 _rnd_reg_q_reg_94_  ( .D(_rnd_reg_N97 ), .CK(clk), .Q(rnd_q[94]),.QN() );
DFF_X2 _rnd_reg_q_reg_95_  ( .D(_rnd_reg_N98 ), .CK(clk), .Q(rnd_q[95]),.QN() );
DFF_X2 _rnd_reg_q_reg_96_  ( .D(_rnd_reg_N99 ), .CK(clk), .Q(rnd_q[96]),.QN() );
DFF_X2 _rnd_reg_q_reg_97_  ( .D(_rnd_reg_N100 ), .CK(clk), .Q(rnd_q[97]),.QN() );
DFF_X2 _rnd_reg_q_reg_98_  ( .D(_rnd_reg_N101 ), .CK(clk), .Q(rnd_q[98]),.QN() );
DFF_X2 _rnd_reg_q_reg_99_  ( .D(_rnd_reg_N102 ), .CK(clk), .Q(rnd_q[99]),.QN() );
DFF_X2 _rnd_reg_q_reg_100_  ( .D(_rnd_reg_N103 ), .CK(clk), .Q(rnd_q[100]),.QN() );
DFF_X2 _rnd_reg_q_reg_101_  ( .D(_rnd_reg_N104 ), .CK(clk), .Q(rnd_q[101]),.QN() );
DFF_X2 _rnd_reg_q_reg_102_  ( .D(_rnd_reg_N105 ), .CK(clk), .Q(rnd_q[102]),.QN() );
DFF_X2 _rnd_reg_q_reg_103_  ( .D(_rnd_reg_N106 ), .CK(clk), .Q(rnd_q[103]),.QN() );
DFF_X2 _rnd_reg_q_reg_104_  ( .D(_rnd_reg_N107 ), .CK(clk), .Q(rnd_q[104]),.QN() );
DFF_X2 _rnd_reg_q_reg_105_  ( .D(_rnd_reg_N108 ), .CK(clk), .Q(rnd_q[105]),.QN() );
DFF_X2 _rnd_reg_q_reg_106_  ( .D(_rnd_reg_N109 ), .CK(clk), .Q(rnd_q[106]),.QN() );
DFF_X2 _rnd_reg_q_reg_107_  ( .D(_rnd_reg_N110 ), .CK(clk), .Q(rnd_q[107]),.QN() );
DFF_X2 _rnd_reg_q_reg_108_  ( .D(_rnd_reg_N111 ), .CK(clk), .Q(rnd_q[108]),.QN() );
DFF_X2 _rnd_reg_q_reg_109_  ( .D(_rnd_reg_N112 ), .CK(clk), .Q(rnd_q[109]),.QN() );
DFF_X2 _rnd_reg_q_reg_110_  ( .D(_rnd_reg_N113 ), .CK(clk), .Q(rnd_q[110]),.QN() );
DFF_X2 _rnd_reg_q_reg_111_  ( .D(_rnd_reg_N114 ), .CK(clk), .Q(rnd_q[111]),.QN() );
DFF_X2 _rnd_reg_q_reg_112_  ( .D(_rnd_reg_N115 ), .CK(clk), .Q(rnd_q[112]),.QN() );
DFF_X2 _rnd_reg_q_reg_113_  ( .D(_rnd_reg_N116 ), .CK(clk), .Q(rnd_q[113]),.QN() );
DFF_X2 _rnd_reg_q_reg_114_  ( .D(_rnd_reg_N117 ), .CK(clk), .Q(rnd_q[114]),.QN() );
DFF_X2 _rnd_reg_q_reg_115_  ( .D(_rnd_reg_N118 ), .CK(clk), .Q(rnd_q[115]),.QN() );
DFF_X2 _rnd_reg_q_reg_116_  ( .D(_rnd_reg_N119 ), .CK(clk), .Q(rnd_q[116]),.QN() );
DFF_X2 _rnd_reg_q_reg_117_  ( .D(_rnd_reg_N120 ), .CK(clk), .Q(rnd_q[117]),.QN() );
DFF_X2 _rnd_reg_q_reg_118_  ( .D(_rnd_reg_N121 ), .CK(clk), .Q(rnd_q[118]),.QN() );
DFF_X2 _rnd_reg_q_reg_119_  ( .D(_rnd_reg_N122 ), .CK(clk), .Q(rnd_q[119]),.QN() );
DFF_X2 _rnd_reg_q_reg_120_  ( .D(_rnd_reg_N123 ), .CK(clk), .Q(rnd_q[120]),.QN() );
DFF_X2 _rnd_reg_q_reg_121_  ( .D(_rnd_reg_N124 ), .CK(clk), .Q(rnd_q[121]),.QN() );
DFF_X2 _rnd_reg_q_reg_122_  ( .D(_rnd_reg_N125 ), .CK(clk), .Q(rnd_q[122]),.QN() );
DFF_X2 _rnd_reg_q_reg_123_  ( .D(_rnd_reg_N126 ), .CK(clk), .Q(rnd_q[123]),.QN() );
DFF_X2 _rnd_reg_q_reg_124_  ( .D(_rnd_reg_N127 ), .CK(clk), .Q(rnd_q[124]),.QN() );
DFF_X2 _rnd_reg_q_reg_125_  ( .D(_rnd_reg_N128 ), .CK(clk), .Q(rnd_q[125]),.QN() );
DFF_X2 _rnd_reg_q_reg_126_  ( .D(_rnd_reg_N129 ), .CK(clk), .Q(rnd_q[126]),.QN() );
DFF_X2 _rnd_reg_q_reg_127_  ( .D(_rnd_reg_N130 ), .CK(clk), .Q(rnd_q[127]),.QN() );
DFF_X2 _rnd_reg_q_reg_128_  ( .D(_rnd_reg_N131 ), .CK(clk), .Q(rnd_q[128]),.QN() );
DFF_X2 _rnd_reg_q_reg_129_  ( .D(_rnd_reg_N132 ), .CK(clk), .Q(rnd_q[129]),.QN() );
DFF_X2 _rnd_reg_q_reg_130_  ( .D(_rnd_reg_N133 ), .CK(clk), .Q(rnd_q[130]),.QN() );
DFF_X2 _rnd_reg_q_reg_131_  ( .D(_rnd_reg_N134 ), .CK(clk), .Q(rnd_q[131]),.QN() );
DFF_X2 _rnd_reg_q_reg_132_  ( .D(_rnd_reg_N135 ), .CK(clk), .Q(rnd_q[132]),.QN() );
DFF_X2 _rnd_reg_q_reg_133_  ( .D(_rnd_reg_N136 ), .CK(clk), .Q(rnd_q[133]),.QN() );
DFF_X2 _rnd_reg_q_reg_134_  ( .D(_rnd_reg_N137 ), .CK(clk), .Q(rnd_q[134]),.QN() );
DFF_X2 _rnd_reg_q_reg_135_  ( .D(_rnd_reg_N138 ), .CK(clk), .Q(rnd_q[135]),.QN() );
DFF_X2 _rnd_reg_q_reg_136_  ( .D(_rnd_reg_N139 ), .CK(clk), .Q(rnd_q[136]),.QN() );
DFF_X2 _rnd_reg_q_reg_137_  ( .D(_rnd_reg_N140 ), .CK(clk), .Q(rnd_q[137]),.QN() );
DFF_X2 _rnd_reg_q_reg_138_  ( .D(_rnd_reg_N141 ), .CK(clk), .Q(rnd_q[138]),.QN() );
DFF_X2 _rnd_reg_q_reg_139_  ( .D(_rnd_reg_N142 ), .CK(clk), .Q(rnd_q[139]),.QN() );
DFF_X2 _rnd_reg_q_reg_140_  ( .D(_rnd_reg_N143 ), .CK(clk), .Q(rnd_q[140]),.QN() );
DFF_X2 _rnd_reg_q_reg_141_  ( .D(_rnd_reg_N144 ), .CK(clk), .Q(rnd_q[141]),.QN() );
DFF_X2 _rnd_reg_q_reg_142_  ( .D(_rnd_reg_N145 ), .CK(clk), .Q(rnd_q[142]),.QN() );
DFF_X2 _rnd_reg_q_reg_143_  ( .D(_rnd_reg_N146 ), .CK(clk), .Q(rnd_q[143]),.QN() );
DFF_X2 _rnd_reg_q_reg_144_  ( .D(_rnd_reg_N147 ), .CK(clk), .Q(rnd_q[144]),.QN() );
DFF_X2 _rnd_reg_q_reg_145_  ( .D(_rnd_reg_N148 ), .CK(clk), .Q(rnd_q[145]),.QN() );
DFF_X2 _rnd_reg_q_reg_146_  ( .D(_rnd_reg_N149 ), .CK(clk), .Q(rnd_q[146]),.QN() );
DFF_X2 _rnd_reg_q_reg_147_  ( .D(_rnd_reg_N150 ), .CK(clk), .Q(rnd_q[147]),.QN() );
DFF_X2 _rnd_reg_q_reg_148_  ( .D(_rnd_reg_N151 ), .CK(clk), .Q(rnd_q[148]),.QN() );
DFF_X2 _rnd_reg_q_reg_149_  ( .D(_rnd_reg_N152 ), .CK(clk), .Q(rnd_q[149]),.QN() );
DFF_X2 _rnd_reg_q_reg_152_  ( .D(_rnd_reg_N155 ), .CK(clk), .Q(rnd_q[152]),.QN() );
AND2_X2 _cv_next_reg_U178  ( .A1(cv_next_d[159]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N162 ) );
AND2_X2 _cv_next_reg_U177  ( .A1(cv_next_d[158]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N161 ) );
AND2_X2 _cv_next_reg_U176  ( .A1(cv_next_d[157]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N160 ) );
AND2_X2 _cv_next_reg_U175  ( .A1(cv_next_d[156]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N159 ) );
AND2_X2 _cv_next_reg_U174  ( .A1(cv_next_d[155]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N158 ) );
AND2_X2 _cv_next_reg_U173  ( .A1(cv_next_d[154]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N157 ) );
AND2_X2 _cv_next_reg_U172  ( .A1(cv_next_d[153]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N156 ) );
AND2_X2 _cv_next_reg_U171  ( .A1(cv_next_d[152]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N155 ) );
AND2_X2 _cv_next_reg_U170  ( .A1(cv_next_d[151]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N154 ) );
AND2_X2 _cv_next_reg_U169  ( .A1(cv_next_d[150]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N153 ) );
AND2_X2 _cv_next_reg_U168  ( .A1(cv_next_d[149]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N152 ) );
AND2_X2 _cv_next_reg_U167  ( .A1(cv_next_d[148]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N151 ) );
AND2_X2 _cv_next_reg_U166  ( .A1(cv_next_d[147]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N150 ) );
AND2_X2 _cv_next_reg_U165  ( .A1(cv_next_d[146]), .A2(_cv_next_reg_n230 ),.ZN(_cv_next_reg_N149 ) );
AND2_X2 _cv_next_reg_U164  ( .A1(cv_next_d[145]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N148 ) );
AND2_X2 _cv_next_reg_U163  ( .A1(cv_next_d[144]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N147 ) );
AND2_X2 _cv_next_reg_U145  ( .A1(cv_next_d[127]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N130 ) );
AND2_X2 _cv_next_reg_U144  ( .A1(cv_next_d[126]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N129 ) );
AND2_X2 _cv_next_reg_U143  ( .A1(cv_next_d[125]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N128 ) );
AND2_X2 _cv_next_reg_U142  ( .A1(cv_next_d[124]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N127 ) );
AND2_X2 _cv_next_reg_U141  ( .A1(cv_next_d[123]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N126 ) );
AND2_X2 _cv_next_reg_U139  ( .A1(cv_next_d[122]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N125 ) );
AND2_X2 _cv_next_reg_U138  ( .A1(cv_next_d[121]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N124 ) );
AND2_X2 _cv_next_reg_U137  ( .A1(cv_next_d[120]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N123 ) );
AND2_X2 _cv_next_reg_U136  ( .A1(cv_next_d[119]), .A2(_cv_next_reg_n220 ),.ZN(_cv_next_reg_N122 ) );
AND2_X2 _cv_next_reg_U135  ( .A1(cv_next_d[118]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N121 ) );
AND2_X2 _cv_next_reg_U134  ( .A1(cv_next_d[117]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N120 ) );
AND2_X2 _cv_next_reg_U133  ( .A1(cv_next_d[116]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N119 ) );
AND2_X2 _cv_next_reg_U132  ( .A1(cv_next_d[115]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N118 ) );
AND2_X2 _cv_next_reg_U131  ( .A1(cv_next_d[114]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N117 ) );
AND2_X2 _cv_next_reg_U130  ( .A1(cv_next_d[113]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N116 ) );
AND2_X2 _cv_next_reg_U128  ( .A1(cv_next_d[112]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N115 ) );
AND2_X2 _cv_next_reg_U110  ( .A1(cv_next_d[95]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N98 ) );
AND2_X2 _cv_next_reg_U109  ( .A1(cv_next_d[94]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N97 ) );
AND2_X2 _cv_next_reg_U108  ( .A1(cv_next_d[93]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N96 ) );
AND2_X2 _cv_next_reg_U106  ( .A1(cv_next_d[92]), .A2(_cv_next_reg_n210 ),.ZN(_cv_next_reg_N95 ) );
AND2_X2 _cv_next_reg_U105  ( .A1(cv_next_d[91]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N94 ) );
AND2_X2 _cv_next_reg_U104  ( .A1(cv_next_d[90]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N93 ) );
AND2_X2 _cv_next_reg_U103  ( .A1(cv_next_d[89]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N92 ) );
AND2_X2 _cv_next_reg_U102  ( .A1(cv_next_d[88]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N91 ) );
AND2_X2 _cv_next_reg_U101  ( .A1(cv_next_d[87]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N90 ) );
AND2_X2 _cv_next_reg_U100  ( .A1(cv_next_d[86]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N89 ) );
AND2_X2 _cv_next_reg_U99  ( .A1(cv_next_d[85]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N88 ) );
AND2_X2 _cv_next_reg_U98  ( .A1(cv_next_d[84]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N87 ) );
AND2_X2 _cv_next_reg_U97  ( .A1(cv_next_d[83]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N86 ) );
AND2_X2 _cv_next_reg_U95  ( .A1(cv_next_d[82]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N85 ) );
AND2_X2 _cv_next_reg_U94  ( .A1(cv_next_d[81]), .A2(_cv_next_reg_n200 ),.ZN(_cv_next_reg_N84 ) );
AND2_X2 _cv_next_reg_U93  ( .A1(cv_next_d[80]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N83 ) );
AND2_X2 _cv_next_reg_U90  ( .A1(cv_next_d[63]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N66 ) );
AND2_X2 _cv_next_reg_U89  ( .A1(cv_next_d[62]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N65 ) );
AND2_X2 _cv_next_reg_U88  ( .A1(cv_next_d[61]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N64 ) );
AND2_X2 _cv_next_reg_U87  ( .A1(cv_next_d[60]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N63 ) );
AND2_X2 _cv_next_reg_U86  ( .A1(cv_next_d[59]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N62 ) );
AND2_X2 _cv_next_reg_U85  ( .A1(cv_next_d[58]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N61 ) );
AND2_X2 _cv_next_reg_U84  ( .A1(cv_next_d[57]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N60 ) );
AND2_X2 _cv_next_reg_U83  ( .A1(cv_next_d[56]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N59 ) );
AND2_X2 _cv_next_reg_U82  ( .A1(cv_next_d[55]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N58 ) );
AND2_X2 _cv_next_reg_U81  ( .A1(cv_next_d[54]), .A2(_cv_next_reg_n190 ),.ZN(_cv_next_reg_N57 ) );
AND2_X2 _cv_next_reg_U80  ( .A1(cv_next_d[53]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N56 ) );
AND2_X2 _cv_next_reg_U78  ( .A1(cv_next_d[52]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N55 ) );
AND2_X2 _cv_next_reg_U77  ( .A1(cv_next_d[51]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N54 ) );
AND2_X2 _cv_next_reg_U76  ( .A1(cv_next_d[50]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N53 ) );
AND2_X2 _cv_next_reg_U75  ( .A1(cv_next_d[49]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N52 ) );
AND2_X2 _cv_next_reg_U74  ( .A1(cv_next_d[48]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N51 ) );
AND2_X2 _cv_next_reg_U55  ( .A1(cv_next_d[31]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N34 ) );
AND2_X2 _cv_next_reg_U54  ( .A1(cv_next_d[30]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N33 ) );
AND2_X2 _cv_next_reg_U53  ( .A1(cv_next_d[29]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N32 ) );
AND2_X2 _cv_next_reg_U52  ( .A1(cv_next_d[28]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N31 ) );
AND2_X2 _cv_next_reg_U51  ( .A1(cv_next_d[27]), .A2(_cv_next_reg_n180 ),.ZN(_cv_next_reg_N30 ) );
AND2_X2 _cv_next_reg_U50  ( .A1(cv_next_d[26]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N29 ) );
AND2_X2 _cv_next_reg_U49  ( .A1(cv_next_d[25]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N28 ) );
AND2_X2 _cv_next_reg_U48  ( .A1(cv_next_d[24]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N27 ) );
AND2_X2 _cv_next_reg_U47  ( .A1(cv_next_d[23]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N26 ) );
AND2_X2 _cv_next_reg_U45  ( .A1(cv_next_d[22]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N25 ) );
AND2_X2 _cv_next_reg_U44  ( .A1(cv_next_d[21]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N24 ) );
AND2_X2 _cv_next_reg_U43  ( .A1(cv_next_d[20]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N23 ) );
AND2_X2 _cv_next_reg_U42  ( .A1(cv_next_d[19]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N22 ) );
AND2_X2 _cv_next_reg_U41  ( .A1(cv_next_d[18]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N21 ) );
AND2_X2 _cv_next_reg_U40  ( .A1(cv_next_d[17]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N20 ) );
AND2_X2 _cv_next_reg_U39  ( .A1(cv_next_d[16]), .A2(_cv_next_reg_n170 ),.ZN(_cv_next_reg_N19 ) );
INV_X4 _cv_next_reg_U20  ( .A(_cv_next_reg_n250 ), .ZN(_cv_next_reg_n320 ));
INV_X4 _cv_next_reg_U19  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n310 ));
INV_X4 _cv_next_reg_U18  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n220 ));
INV_X4 _cv_next_reg_U17  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n210 ));
INV_X4 _cv_next_reg_U16  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n200 ));
INV_X4 _cv_next_reg_U15  ( .A(n7117), .ZN(_cv_next_reg_n190 ) );
INV_X4 _cv_next_reg_U14  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n180 ));
INV_X4 _cv_next_reg_U12  ( .A(n7117), .ZN(_cv_next_reg_n170 ) );
INV_X4 _cv_next_reg_U11  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n240 ));
INV_X4 _cv_next_reg_U10  ( .A(n7117), .ZN(_cv_next_reg_n230 ) );
INV_X4 _cv_next_reg_U9  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n280 ) );
INV_X4 _cv_next_reg_U8  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n290 ) );
INV_X4 _cv_next_reg_U7  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n300 ) );
INV_X4 _cv_next_reg_U6  ( .A(n7117), .ZN(_cv_next_reg_n250 ) );
INV_X4 _cv_next_reg_U5  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n260 ) );
INV_X4 _cv_next_reg_U4  ( .A(_cv_next_reg_n320 ), .ZN(_cv_next_reg_n270 ) );
AND2_X2 _cv_next_reg_U162  ( .A1(cv_next_d[7]), .A2(_cv_next_reg_n310 ),.ZN(_cv_next_reg_N10 ) );
AND2_X2 _cv_next_reg_U161  ( .A1(cv_next_d[97]), .A2(_cv_next_reg_n310 ),.ZN(_cv_next_reg_N100 ) );
AND2_X2 _cv_next_reg_U160  ( .A1(cv_next_d[98]), .A2(_cv_next_reg_n310 ),.ZN(_cv_next_reg_N101 ) );
AND2_X2 _cv_next_reg_U159  ( .A1(cv_next_d[99]), .A2(_cv_next_reg_n310 ),.ZN(_cv_next_reg_N102 ) );
AND2_X2 _cv_next_reg_U158  ( .A1(cv_next_d[100]), .A2(_cv_next_reg_n310 ),.ZN(_cv_next_reg_N103 ) );
AND2_X2 _cv_next_reg_U157  ( .A1(cv_next_d[101]), .A2(_cv_next_reg_n310 ),.ZN(_cv_next_reg_N104 ) );
AND2_X2 _cv_next_reg_U156  ( .A1(cv_next_d[102]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N105 ) );
AND2_X2 _cv_next_reg_U155  ( .A1(cv_next_d[103]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N106 ) );
AND2_X2 _cv_next_reg_U154  ( .A1(cv_next_d[104]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N107 ) );
AND2_X2 _cv_next_reg_U153  ( .A1(cv_next_d[105]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N108 ) );
AND2_X2 _cv_next_reg_U152  ( .A1(cv_next_d[106]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N109 ) );
AND2_X2 _cv_next_reg_U151  ( .A1(cv_next_d[8]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N11 ) );
AND2_X2 _cv_next_reg_U150  ( .A1(cv_next_d[107]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N110 ) );
AND2_X2 _cv_next_reg_U149  ( .A1(cv_next_d[108]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N111 ) );
AND2_X2 _cv_next_reg_U148  ( .A1(cv_next_d[109]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N112 ) );
AND2_X2 _cv_next_reg_U147  ( .A1(cv_next_d[110]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N113 ) );
AND2_X2 _cv_next_reg_U146  ( .A1(cv_next_d[111]), .A2(_cv_next_reg_n300 ),.ZN(_cv_next_reg_N114 ) );
AND2_X2 _cv_next_reg_U140  ( .A1(cv_next_d[9]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N12 ) );
AND2_X2 _cv_next_reg_U129  ( .A1(cv_next_d[10]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N13 ) );
AND2_X2 _cv_next_reg_U127  ( .A1(cv_next_d[128]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N131 ) );
AND2_X2 _cv_next_reg_U126  ( .A1(cv_next_d[129]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N132 ) );
AND2_X2 _cv_next_reg_U125  ( .A1(cv_next_d[130]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N133 ) );
AND2_X2 _cv_next_reg_U124  ( .A1(cv_next_d[131]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N134 ) );
AND2_X2 _cv_next_reg_U123  ( .A1(cv_next_d[132]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N135 ) );
AND2_X2 _cv_next_reg_U122  ( .A1(cv_next_d[133]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N136 ) );
AND2_X2 _cv_next_reg_U121  ( .A1(cv_next_d[134]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N137 ) );
AND2_X2 _cv_next_reg_U120  ( .A1(cv_next_d[135]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N138 ) );
AND2_X2 _cv_next_reg_U119  ( .A1(cv_next_d[136]), .A2(_cv_next_reg_n290 ),.ZN(_cv_next_reg_N139 ) );
AND2_X2 _cv_next_reg_U118  ( .A1(cv_next_d[11]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N14 ) );
AND2_X2 _cv_next_reg_U117  ( .A1(cv_next_d[137]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N140 ) );
AND2_X2 _cv_next_reg_U116  ( .A1(cv_next_d[138]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N141 ) );
AND2_X2 _cv_next_reg_U115  ( .A1(cv_next_d[139]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N142 ) );
AND2_X2 _cv_next_reg_U114  ( .A1(cv_next_d[140]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N143 ) );
AND2_X2 _cv_next_reg_U113  ( .A1(cv_next_d[141]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N144 ) );
AND2_X2 _cv_next_reg_U112  ( .A1(cv_next_d[142]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N145 ) );
AND2_X2 _cv_next_reg_U111  ( .A1(cv_next_d[143]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N146 ) );
AND2_X2 _cv_next_reg_U107  ( .A1(cv_next_d[12]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N15 ) );
AND2_X2 _cv_next_reg_U96  ( .A1(cv_next_d[13]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N16 ) );
AND2_X2 _cv_next_reg_U92  ( .A1(cv_next_d[14]), .A2(_cv_next_reg_n280 ),.ZN(_cv_next_reg_N17 ) );
AND2_X2 _cv_next_reg_U91  ( .A1(cv_next_d[15]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N18 ) );
AND2_X2 _cv_next_reg_U79  ( .A1(cv_next_d[0]), .A2(_cv_next_reg_n270 ), .ZN(_cv_next_reg_N3 ) );
AND2_X2 _cv_next_reg_U73  ( .A1(cv_next_d[32]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N35 ) );
AND2_X2 _cv_next_reg_U72  ( .A1(cv_next_d[33]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N36 ) );
AND2_X2 _cv_next_reg_U71  ( .A1(cv_next_d[34]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N37 ) );
AND2_X2 _cv_next_reg_U70  ( .A1(cv_next_d[35]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N38 ) );
AND2_X2 _cv_next_reg_U69  ( .A1(cv_next_d[36]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N39 ) );
AND2_X2 _cv_next_reg_U68  ( .A1(cv_next_d[1]), .A2(_cv_next_reg_n270 ), .ZN(_cv_next_reg_N4 ) );
AND2_X2 _cv_next_reg_U67  ( .A1(cv_next_d[37]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N40 ) );
AND2_X2 _cv_next_reg_U66  ( .A1(cv_next_d[38]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N41 ) );
AND2_X2 _cv_next_reg_U65  ( .A1(cv_next_d[39]), .A2(_cv_next_reg_n270 ),.ZN(_cv_next_reg_N42 ) );
AND2_X2 _cv_next_reg_U64  ( .A1(cv_next_d[40]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N43 ) );
AND2_X2 _cv_next_reg_U63  ( .A1(cv_next_d[41]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N44 ) );
AND2_X2 _cv_next_reg_U62  ( .A1(cv_next_d[42]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N45 ) );
AND2_X2 _cv_next_reg_U61  ( .A1(cv_next_d[43]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N46 ) );
AND2_X2 _cv_next_reg_U60  ( .A1(cv_next_d[44]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N47 ) );
AND2_X2 _cv_next_reg_U59  ( .A1(cv_next_d[45]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N48 ) );
AND2_X2 _cv_next_reg_U58  ( .A1(cv_next_d[46]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N49 ) );
AND2_X2 _cv_next_reg_U57  ( .A1(cv_next_d[2]), .A2(_cv_next_reg_n260 ), .ZN(_cv_next_reg_N5 ) );
AND2_X2 _cv_next_reg_U56  ( .A1(cv_next_d[47]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N50 ) );
AND2_X2 _cv_next_reg_U46  ( .A1(cv_next_d[3]), .A2(_cv_next_reg_n260 ), .ZN(_cv_next_reg_N6 ) );
AND2_X2 _cv_next_reg_U38  ( .A1(cv_next_d[64]), .A2(_cv_next_reg_n260 ),.ZN(_cv_next_reg_N67 ) );
AND2_X2 _cv_next_reg_U37  ( .A1(cv_next_d[65]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N68 ) );
AND2_X2 _cv_next_reg_U36  ( .A1(cv_next_d[66]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N69 ) );
AND2_X2 _cv_next_reg_U35  ( .A1(cv_next_d[4]), .A2(_cv_next_reg_n250 ), .ZN(_cv_next_reg_N7 ) );
AND2_X2 _cv_next_reg_U34  ( .A1(cv_next_d[67]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N70 ) );
AND2_X2 _cv_next_reg_U33  ( .A1(cv_next_d[68]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N71 ) );
AND2_X2 _cv_next_reg_U32  ( .A1(cv_next_d[69]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N72 ) );
AND2_X2 _cv_next_reg_U31  ( .A1(cv_next_d[70]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N73 ) );
AND2_X2 _cv_next_reg_U30  ( .A1(cv_next_d[71]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N74 ) );
AND2_X2 _cv_next_reg_U29  ( .A1(cv_next_d[72]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N75 ) );
AND2_X2 _cv_next_reg_U28  ( .A1(cv_next_d[73]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N76 ) );
AND2_X2 _cv_next_reg_U27  ( .A1(cv_next_d[74]), .A2(_cv_next_reg_n250 ),.ZN(_cv_next_reg_N77 ) );
AND2_X2 _cv_next_reg_U26  ( .A1(cv_next_d[75]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N78 ) );
AND2_X2 _cv_next_reg_U25  ( .A1(cv_next_d[76]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N79 ) );
AND2_X2 _cv_next_reg_U24  ( .A1(cv_next_d[5]), .A2(_cv_next_reg_n240 ), .ZN(_cv_next_reg_N8 ) );
AND2_X2 _cv_next_reg_U23  ( .A1(cv_next_d[77]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N80 ) );
AND2_X2 _cv_next_reg_U22  ( .A1(cv_next_d[78]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N81 ) );
AND2_X2 _cv_next_reg_U21  ( .A1(cv_next_d[79]), .A2(_cv_next_reg_n240 ),.ZN(_cv_next_reg_N82 ) );
AND2_X2 _cv_next_reg_U13  ( .A1(cv_next_d[6]), .A2(_cv_next_reg_n240 ), .ZN(_cv_next_reg_N9 ) );
AND2_X2 _cv_next_reg_U3  ( .A1(cv_next_d[96]), .A2(_cv_next_reg_n240 ), .ZN(_cv_next_reg_N99 ) );
DFF_X2 _cv_next_reg_q_reg_0_  ( .D(_cv_next_reg_N3 ), .CK(clk), .Q(cv_next[0]), .QN() );
DFF_X2 _cv_next_reg_q_reg_1_  ( .D(_cv_next_reg_N4 ), .CK(clk), .Q(cv_next[1]), .QN() );
DFF_X2 _cv_next_reg_q_reg_2_  ( .D(_cv_next_reg_N5 ), .CK(clk), .Q(cv_next[2]), .QN() );
DFF_X2 _cv_next_reg_q_reg_3_  ( .D(_cv_next_reg_N6 ), .CK(clk), .Q(cv_next[3]), .QN() );
DFF_X2 _cv_next_reg_q_reg_4_  ( .D(_cv_next_reg_N7 ), .CK(clk), .Q(cv_next[4]), .QN() );
DFF_X2 _cv_next_reg_q_reg_5_  ( .D(_cv_next_reg_N8 ), .CK(clk), .Q(cv_next[5]), .QN() );
DFF_X2 _cv_next_reg_q_reg_6_  ( .D(_cv_next_reg_N9 ), .CK(clk), .Q(cv_next[6]), .QN() );
DFF_X2 _cv_next_reg_q_reg_7_  ( .D(_cv_next_reg_N10 ), .CK(clk), .Q(cv_next[7]), .QN() );
DFF_X2 _cv_next_reg_q_reg_8_  ( .D(_cv_next_reg_N11 ), .CK(clk), .Q(cv_next[8]), .QN() );
DFF_X2 _cv_next_reg_q_reg_9_  ( .D(_cv_next_reg_N12 ), .CK(clk), .Q(cv_next[9]), .QN() );
DFF_X2 _cv_next_reg_q_reg_10_  ( .D(_cv_next_reg_N13 ), .CK(clk), .Q(cv_next[10]), .QN() );
DFF_X2 _cv_next_reg_q_reg_11_  ( .D(_cv_next_reg_N14 ), .CK(clk), .Q(cv_next[11]), .QN() );
DFF_X2 _cv_next_reg_q_reg_12_  ( .D(_cv_next_reg_N15 ), .CK(clk), .Q(cv_next[12]), .QN() );
DFF_X2 _cv_next_reg_q_reg_13_  ( .D(_cv_next_reg_N16 ), .CK(clk), .Q(cv_next[13]), .QN() );
DFF_X2 _cv_next_reg_q_reg_14_  ( .D(_cv_next_reg_N17 ), .CK(clk), .Q(cv_next[14]), .QN() );
DFF_X2 _cv_next_reg_q_reg_15_  ( .D(_cv_next_reg_N18 ), .CK(clk), .Q(cv_next[15]), .QN() );
DFF_X2 _cv_next_reg_q_reg_16_  ( .D(_cv_next_reg_N19 ), .CK(clk), .Q(cv_next[16]), .QN() );
DFF_X2 _cv_next_reg_q_reg_17_  ( .D(_cv_next_reg_N20 ), .CK(clk), .Q(cv_next[17]), .QN() );
DFF_X2 _cv_next_reg_q_reg_18_  ( .D(_cv_next_reg_N21 ), .CK(clk), .Q(cv_next[18]), .QN() );
DFF_X2 _cv_next_reg_q_reg_19_  ( .D(_cv_next_reg_N22 ), .CK(clk), .Q(cv_next[19]), .QN() );
DFF_X2 _cv_next_reg_q_reg_20_  ( .D(_cv_next_reg_N23 ), .CK(clk), .Q(cv_next[20]), .QN() );
DFF_X2 _cv_next_reg_q_reg_21_  ( .D(_cv_next_reg_N24 ), .CK(clk), .Q(cv_next[21]), .QN() );
DFF_X2 _cv_next_reg_q_reg_22_  ( .D(_cv_next_reg_N25 ), .CK(clk), .Q(cv_next[22]), .QN() );
DFF_X2 _cv_next_reg_q_reg_23_  ( .D(_cv_next_reg_N26 ), .CK(clk), .Q(cv_next[23]), .QN() );
DFF_X2 _cv_next_reg_q_reg_24_  ( .D(_cv_next_reg_N27 ), .CK(clk), .Q(cv_next[24]), .QN() );
DFF_X2 _cv_next_reg_q_reg_25_  ( .D(_cv_next_reg_N28 ), .CK(clk), .Q(cv_next[25]), .QN() );
DFF_X2 _cv_next_reg_q_reg_26_  ( .D(_cv_next_reg_N29 ), .CK(clk), .Q(cv_next[26]), .QN() );
DFF_X2 _cv_next_reg_q_reg_27_  ( .D(_cv_next_reg_N30 ), .CK(clk), .Q(cv_next[27]), .QN() );
DFF_X2 _cv_next_reg_q_reg_28_  ( .D(_cv_next_reg_N31 ), .CK(clk), .Q(cv_next[28]), .QN() );
DFF_X2 _cv_next_reg_q_reg_29_  ( .D(_cv_next_reg_N32 ), .CK(clk), .Q(cv_next[29]), .QN() );
DFF_X2 _cv_next_reg_q_reg_30_  ( .D(_cv_next_reg_N33 ), .CK(clk), .Q(cv_next[30]), .QN() );
DFF_X2 _cv_next_reg_q_reg_31_  ( .D(_cv_next_reg_N34 ), .CK(clk), .Q(cv_next[31]), .QN() );
DFF_X2 _cv_next_reg_q_reg_32_  ( .D(_cv_next_reg_N35 ), .CK(clk), .Q(cv_next[32]), .QN() );
DFF_X2 _cv_next_reg_q_reg_33_  ( .D(_cv_next_reg_N36 ), .CK(clk), .Q(cv_next[33]), .QN() );
DFF_X2 _cv_next_reg_q_reg_34_  ( .D(_cv_next_reg_N37 ), .CK(clk), .Q(cv_next[34]), .QN() );
DFF_X2 _cv_next_reg_q_reg_35_  ( .D(_cv_next_reg_N38 ), .CK(clk), .Q(cv_next[35]), .QN() );
DFF_X2 _cv_next_reg_q_reg_36_  ( .D(_cv_next_reg_N39 ), .CK(clk), .Q(cv_next[36]), .QN() );
DFF_X2 _cv_next_reg_q_reg_37_  ( .D(_cv_next_reg_N40 ), .CK(clk), .Q(cv_next[37]), .QN() );
DFF_X2 _cv_next_reg_q_reg_38_  ( .D(_cv_next_reg_N41 ), .CK(clk), .Q(cv_next[38]), .QN() );
DFF_X2 _cv_next_reg_q_reg_39_  ( .D(_cv_next_reg_N42 ), .CK(clk), .Q(cv_next[39]), .QN() );
DFF_X2 _cv_next_reg_q_reg_40_  ( .D(_cv_next_reg_N43 ), .CK(clk), .Q(cv_next[40]), .QN() );
DFF_X2 _cv_next_reg_q_reg_41_  ( .D(_cv_next_reg_N44 ), .CK(clk), .Q(cv_next[41]), .QN() );
DFF_X2 _cv_next_reg_q_reg_42_  ( .D(_cv_next_reg_N45 ), .CK(clk), .Q(cv_next[42]), .QN() );
DFF_X2 _cv_next_reg_q_reg_43_  ( .D(_cv_next_reg_N46 ), .CK(clk), .Q(cv_next[43]), .QN() );
DFF_X2 _cv_next_reg_q_reg_44_  ( .D(_cv_next_reg_N47 ), .CK(clk), .Q(cv_next[44]), .QN() );
DFF_X2 _cv_next_reg_q_reg_45_  ( .D(_cv_next_reg_N48 ), .CK(clk), .Q(cv_next[45]), .QN() );
DFF_X2 _cv_next_reg_q_reg_46_  ( .D(_cv_next_reg_N49 ), .CK(clk), .Q(cv_next[46]), .QN() );
DFF_X2 _cv_next_reg_q_reg_47_  ( .D(_cv_next_reg_N50 ), .CK(clk), .Q(cv_next[47]), .QN() );
DFF_X2 _cv_next_reg_q_reg_48_  ( .D(_cv_next_reg_N51 ), .CK(clk), .Q(cv_next[48]), .QN() );
DFF_X2 _cv_next_reg_q_reg_49_  ( .D(_cv_next_reg_N52 ), .CK(clk), .Q(cv_next[49]), .QN() );
DFF_X2 _cv_next_reg_q_reg_50_  ( .D(_cv_next_reg_N53 ), .CK(clk), .Q(cv_next[50]), .QN() );
DFF_X2 _cv_next_reg_q_reg_51_  ( .D(_cv_next_reg_N54 ), .CK(clk), .Q(cv_next[51]), .QN() );
DFF_X2 _cv_next_reg_q_reg_52_  ( .D(_cv_next_reg_N55 ), .CK(clk), .Q(cv_next[52]), .QN() );
DFF_X2 _cv_next_reg_q_reg_53_  ( .D(_cv_next_reg_N56 ), .CK(clk), .Q(cv_next[53]), .QN() );
DFF_X2 _cv_next_reg_q_reg_54_  ( .D(_cv_next_reg_N57 ), .CK(clk), .Q(cv_next[54]), .QN() );
DFF_X2 _cv_next_reg_q_reg_55_  ( .D(_cv_next_reg_N58 ), .CK(clk), .Q(cv_next[55]), .QN() );
DFF_X2 _cv_next_reg_q_reg_56_  ( .D(_cv_next_reg_N59 ), .CK(clk), .Q(cv_next[56]), .QN() );
DFF_X2 _cv_next_reg_q_reg_57_  ( .D(_cv_next_reg_N60 ), .CK(clk), .Q(cv_next[57]), .QN() );
DFF_X2 _cv_next_reg_q_reg_58_  ( .D(_cv_next_reg_N61 ), .CK(clk), .Q(cv_next[58]), .QN() );
DFF_X2 _cv_next_reg_q_reg_59_  ( .D(_cv_next_reg_N62 ), .CK(clk), .Q(cv_next[59]), .QN() );
DFF_X2 _cv_next_reg_q_reg_60_  ( .D(_cv_next_reg_N63 ), .CK(clk), .Q(cv_next[60]), .QN() );
DFF_X2 _cv_next_reg_q_reg_61_  ( .D(_cv_next_reg_N64 ), .CK(clk), .Q(cv_next[61]), .QN() );
DFF_X2 _cv_next_reg_q_reg_62_  ( .D(_cv_next_reg_N65 ), .CK(clk), .Q(cv_next[62]), .QN() );
DFF_X2 _cv_next_reg_q_reg_63_  ( .D(_cv_next_reg_N66 ), .CK(clk), .Q(cv_next[63]), .QN() );
DFF_X2 _cv_next_reg_q_reg_64_  ( .D(_cv_next_reg_N67 ), .CK(clk), .Q(cv_next[64]), .QN() );
DFF_X2 _cv_next_reg_q_reg_65_  ( .D(_cv_next_reg_N68 ), .CK(clk), .Q(cv_next[65]), .QN() );
DFF_X2 _cv_next_reg_q_reg_66_  ( .D(_cv_next_reg_N69 ), .CK(clk), .Q(cv_next[66]), .QN() );
DFF_X2 _cv_next_reg_q_reg_67_  ( .D(_cv_next_reg_N70 ), .CK(clk), .Q(cv_next[67]), .QN() );
DFF_X2 _cv_next_reg_q_reg_68_  ( .D(_cv_next_reg_N71 ), .CK(clk), .Q(cv_next[68]), .QN() );
DFF_X2 _cv_next_reg_q_reg_69_  ( .D(_cv_next_reg_N72 ), .CK(clk), .Q(cv_next[69]), .QN() );
DFF_X2 _cv_next_reg_q_reg_70_  ( .D(_cv_next_reg_N73 ), .CK(clk), .Q(cv_next[70]), .QN() );
DFF_X2 _cv_next_reg_q_reg_71_  ( .D(_cv_next_reg_N74 ), .CK(clk), .Q(cv_next[71]), .QN() );
DFF_X2 _cv_next_reg_q_reg_72_  ( .D(_cv_next_reg_N75 ), .CK(clk), .Q(cv_next[72]), .QN() );
DFF_X2 _cv_next_reg_q_reg_73_  ( .D(_cv_next_reg_N76 ), .CK(clk), .Q(cv_next[73]), .QN() );
DFF_X2 _cv_next_reg_q_reg_74_  ( .D(_cv_next_reg_N77 ), .CK(clk), .Q(cv_next[74]), .QN() );
DFF_X2 _cv_next_reg_q_reg_75_  ( .D(_cv_next_reg_N78 ), .CK(clk), .Q(cv_next[75]), .QN() );
DFF_X2 _cv_next_reg_q_reg_76_  ( .D(_cv_next_reg_N79 ), .CK(clk), .Q(cv_next[76]), .QN() );
DFF_X2 _cv_next_reg_q_reg_77_  ( .D(_cv_next_reg_N80 ), .CK(clk), .Q(cv_next[77]), .QN() );
DFF_X2 _cv_next_reg_q_reg_78_  ( .D(_cv_next_reg_N81 ), .CK(clk), .Q(cv_next[78]), .QN() );
DFF_X2 _cv_next_reg_q_reg_79_  ( .D(_cv_next_reg_N82 ), .CK(clk), .Q(cv_next[79]), .QN() );
DFF_X2 _cv_next_reg_q_reg_80_  ( .D(_cv_next_reg_N83 ), .CK(clk), .Q(cv_next[80]), .QN() );
DFF_X2 _cv_next_reg_q_reg_81_  ( .D(_cv_next_reg_N84 ), .CK(clk), .Q(cv_next[81]), .QN() );
DFF_X2 _cv_next_reg_q_reg_82_  ( .D(_cv_next_reg_N85 ), .CK(clk), .Q(cv_next[82]), .QN() );
DFF_X2 _cv_next_reg_q_reg_83_  ( .D(_cv_next_reg_N86 ), .CK(clk), .Q(cv_next[83]), .QN() );
DFF_X2 _cv_next_reg_q_reg_84_  ( .D(_cv_next_reg_N87 ), .CK(clk), .Q(cv_next[84]), .QN() );
DFF_X2 _cv_next_reg_q_reg_85_  ( .D(_cv_next_reg_N88 ), .CK(clk), .Q(cv_next[85]), .QN() );
DFF_X2 _cv_next_reg_q_reg_86_  ( .D(_cv_next_reg_N89 ), .CK(clk), .Q(cv_next[86]), .QN() );
DFF_X2 _cv_next_reg_q_reg_87_  ( .D(_cv_next_reg_N90 ), .CK(clk), .Q(cv_next[87]), .QN() );
DFF_X2 _cv_next_reg_q_reg_88_  ( .D(_cv_next_reg_N91 ), .CK(clk), .Q(cv_next[88]), .QN() );
DFF_X2 _cv_next_reg_q_reg_89_  ( .D(_cv_next_reg_N92 ), .CK(clk), .Q(cv_next[89]), .QN() );
DFF_X2 _cv_next_reg_q_reg_90_  ( .D(_cv_next_reg_N93 ), .CK(clk), .Q(cv_next[90]), .QN() );
DFF_X2 _cv_next_reg_q_reg_91_  ( .D(_cv_next_reg_N94 ), .CK(clk), .Q(cv_next[91]), .QN() );
DFF_X2 _cv_next_reg_q_reg_92_  ( .D(_cv_next_reg_N95 ), .CK(clk), .Q(cv_next[92]), .QN() );
DFF_X2 _cv_next_reg_q_reg_93_  ( .D(_cv_next_reg_N96 ), .CK(clk), .Q(cv_next[93]), .QN() );
DFF_X2 _cv_next_reg_q_reg_94_  ( .D(_cv_next_reg_N97 ), .CK(clk), .Q(cv_next[94]), .QN() );
DFF_X2 _cv_next_reg_q_reg_95_  ( .D(_cv_next_reg_N98 ), .CK(clk), .Q(cv_next[95]), .QN() );
DFF_X2 _cv_next_reg_q_reg_96_  ( .D(_cv_next_reg_N99 ), .CK(clk), .Q(cv_next[96]), .QN() );
DFF_X2 _cv_next_reg_q_reg_97_  ( .D(_cv_next_reg_N100 ), .CK(clk), .Q(cv_next[97]), .QN() );
DFF_X2 _cv_next_reg_q_reg_98_  ( .D(_cv_next_reg_N101 ), .CK(clk), .Q(cv_next[98]), .QN() );
DFF_X2 _cv_next_reg_q_reg_99_  ( .D(_cv_next_reg_N102 ), .CK(clk), .Q(cv_next[99]), .QN() );
DFF_X2 _cv_next_reg_q_reg_100_  ( .D(_cv_next_reg_N103 ), .CK(clk), .Q(cv_next[100]), .QN() );
DFF_X2 _cv_next_reg_q_reg_101_  ( .D(_cv_next_reg_N104 ), .CK(clk), .Q(cv_next[101]), .QN() );
DFF_X2 _cv_next_reg_q_reg_102_  ( .D(_cv_next_reg_N105 ), .CK(clk), .Q(cv_next[102]), .QN() );
DFF_X2 _cv_next_reg_q_reg_103_  ( .D(_cv_next_reg_N106 ), .CK(clk), .Q(cv_next[103]), .QN() );
DFF_X2 _cv_next_reg_q_reg_104_  ( .D(_cv_next_reg_N107 ), .CK(clk), .Q(cv_next[104]), .QN() );
DFF_X2 _cv_next_reg_q_reg_105_  ( .D(_cv_next_reg_N108 ), .CK(clk), .Q(cv_next[105]), .QN() );
DFF_X2 _cv_next_reg_q_reg_106_  ( .D(_cv_next_reg_N109 ), .CK(clk), .Q(cv_next[106]), .QN() );
DFF_X2 _cv_next_reg_q_reg_107_  ( .D(_cv_next_reg_N110 ), .CK(clk), .Q(cv_next[107]), .QN() );
DFF_X2 _cv_next_reg_q_reg_108_  ( .D(_cv_next_reg_N111 ), .CK(clk), .Q(cv_next[108]), .QN() );
DFF_X2 _cv_next_reg_q_reg_109_  ( .D(_cv_next_reg_N112 ), .CK(clk), .Q(cv_next[109]), .QN() );
DFF_X2 _cv_next_reg_q_reg_110_  ( .D(_cv_next_reg_N113 ), .CK(clk), .Q(cv_next[110]), .QN() );
DFF_X2 _cv_next_reg_q_reg_111_  ( .D(_cv_next_reg_N114 ), .CK(clk), .Q(cv_next[111]), .QN() );
DFF_X2 _cv_next_reg_q_reg_112_  ( .D(_cv_next_reg_N115 ), .CK(clk), .Q(cv_next[112]), .QN() );
DFF_X2 _cv_next_reg_q_reg_113_  ( .D(_cv_next_reg_N116 ), .CK(clk), .Q(cv_next[113]), .QN() );
DFF_X2 _cv_next_reg_q_reg_114_  ( .D(_cv_next_reg_N117 ), .CK(clk), .Q(cv_next[114]), .QN() );
DFF_X2 _cv_next_reg_q_reg_115_  ( .D(_cv_next_reg_N118 ), .CK(clk), .Q(cv_next[115]), .QN() );
DFF_X2 _cv_next_reg_q_reg_116_  ( .D(_cv_next_reg_N119 ), .CK(clk), .Q(cv_next[116]), .QN() );
DFF_X2 _cv_next_reg_q_reg_117_  ( .D(_cv_next_reg_N120 ), .CK(clk), .Q(cv_next[117]), .QN() );
DFF_X2 _cv_next_reg_q_reg_118_  ( .D(_cv_next_reg_N121 ), .CK(clk), .Q(cv_next[118]), .QN() );
DFF_X2 _cv_next_reg_q_reg_119_  ( .D(_cv_next_reg_N122 ), .CK(clk), .Q(cv_next[119]), .QN() );
DFF_X2 _cv_next_reg_q_reg_120_  ( .D(_cv_next_reg_N123 ), .CK(clk), .Q(cv_next[120]), .QN() );
DFF_X2 _cv_next_reg_q_reg_121_  ( .D(_cv_next_reg_N124 ), .CK(clk), .Q(cv_next[121]), .QN() );
DFF_X2 _cv_next_reg_q_reg_122_  ( .D(_cv_next_reg_N125 ), .CK(clk), .Q(cv_next[122]), .QN() );
DFF_X2 _cv_next_reg_q_reg_123_  ( .D(_cv_next_reg_N126 ), .CK(clk), .Q(cv_next[123]), .QN() );
DFF_X2 _cv_next_reg_q_reg_124_  ( .D(_cv_next_reg_N127 ), .CK(clk), .Q(cv_next[124]), .QN() );
DFF_X2 _cv_next_reg_q_reg_125_  ( .D(_cv_next_reg_N128 ), .CK(clk), .Q(cv_next[125]), .QN() );
DFF_X2 _cv_next_reg_q_reg_126_  ( .D(_cv_next_reg_N129 ), .CK(clk), .Q(cv_next[126]), .QN() );
DFF_X2 _cv_next_reg_q_reg_127_  ( .D(_cv_next_reg_N130 ), .CK(clk), .Q(cv_next[127]), .QN() );
DFF_X2 _cv_next_reg_q_reg_128_  ( .D(_cv_next_reg_N131 ), .CK(clk), .Q(cv_next[128]), .QN() );
DFF_X2 _cv_next_reg_q_reg_129_  ( .D(_cv_next_reg_N132 ), .CK(clk), .Q(cv_next[129]), .QN() );
DFF_X2 _cv_next_reg_q_reg_130_  ( .D(_cv_next_reg_N133 ), .CK(clk), .Q(cv_next[130]), .QN() );
DFF_X2 _cv_next_reg_q_reg_131_  ( .D(_cv_next_reg_N134 ), .CK(clk), .Q(cv_next[131]), .QN() );
DFF_X2 _cv_next_reg_q_reg_132_  ( .D(_cv_next_reg_N135 ), .CK(clk), .Q(cv_next[132]), .QN() );
DFF_X2 _cv_next_reg_q_reg_133_  ( .D(_cv_next_reg_N136 ), .CK(clk), .Q(cv_next[133]), .QN() );
DFF_X2 _cv_next_reg_q_reg_134_  ( .D(_cv_next_reg_N137 ), .CK(clk), .Q(cv_next[134]), .QN() );
DFF_X2 _cv_next_reg_q_reg_135_  ( .D(_cv_next_reg_N138 ), .CK(clk), .Q(cv_next[135]), .QN() );
DFF_X2 _cv_next_reg_q_reg_136_  ( .D(_cv_next_reg_N139 ), .CK(clk), .Q(cv_next[136]), .QN() );
DFF_X2 _cv_next_reg_q_reg_137_  ( .D(_cv_next_reg_N140 ), .CK(clk), .Q(cv_next[137]), .QN() );
DFF_X2 _cv_next_reg_q_reg_138_  ( .D(_cv_next_reg_N141 ), .CK(clk), .Q(cv_next[138]), .QN() );
DFF_X2 _cv_next_reg_q_reg_139_  ( .D(_cv_next_reg_N142 ), .CK(clk), .Q(cv_next[139]), .QN() );
DFF_X2 _cv_next_reg_q_reg_140_  ( .D(_cv_next_reg_N143 ), .CK(clk), .Q(cv_next[140]), .QN() );
DFF_X2 _cv_next_reg_q_reg_141_  ( .D(_cv_next_reg_N144 ), .CK(clk), .Q(cv_next[141]), .QN() );
DFF_X2 _cv_next_reg_q_reg_142_  ( .D(_cv_next_reg_N145 ), .CK(clk), .Q(cv_next[142]), .QN() );
DFF_X2 _cv_next_reg_q_reg_143_  ( .D(_cv_next_reg_N146 ), .CK(clk), .Q(cv_next[143]), .QN() );
DFF_X2 _cv_next_reg_q_reg_144_  ( .D(_cv_next_reg_N147 ), .CK(clk), .Q(cv_next[144]), .QN() );
DFF_X2 _cv_next_reg_q_reg_145_  ( .D(_cv_next_reg_N148 ), .CK(clk), .Q(cv_next[145]), .QN() );
DFF_X2 _cv_next_reg_q_reg_146_  ( .D(_cv_next_reg_N149 ), .CK(clk), .Q(cv_next[146]), .QN() );
DFF_X2 _cv_next_reg_q_reg_147_  ( .D(_cv_next_reg_N150 ), .CK(clk), .Q(cv_next[147]), .QN() );
DFF_X2 _cv_next_reg_q_reg_148_  ( .D(_cv_next_reg_N151 ), .CK(clk), .Q(cv_next[148]), .QN() );
DFF_X2 _cv_next_reg_q_reg_149_  ( .D(_cv_next_reg_N152 ), .CK(clk), .Q(cv_next[149]), .QN() );
DFF_X2 _cv_next_reg_q_reg_150_  ( .D(_cv_next_reg_N153 ), .CK(clk), .Q(cv_next[150]), .QN() );
DFF_X2 _cv_next_reg_q_reg_151_  ( .D(_cv_next_reg_N154 ), .CK(clk), .Q(cv_next[151]), .QN() );
DFF_X2 _cv_next_reg_q_reg_152_  ( .D(_cv_next_reg_N155 ), .CK(clk), .Q(cv_next[152]), .QN() );
DFF_X2 _cv_next_reg_q_reg_153_  ( .D(_cv_next_reg_N156 ), .CK(clk), .Q(cv_next[153]), .QN() );
DFF_X2 _cv_next_reg_q_reg_154_  ( .D(_cv_next_reg_N157 ), .CK(clk), .Q(cv_next[154]), .QN() );
DFF_X2 _cv_next_reg_q_reg_155_  ( .D(_cv_next_reg_N158 ), .CK(clk), .Q(cv_next[155]), .QN() );
DFF_X2 _cv_next_reg_q_reg_156_  ( .D(_cv_next_reg_N159 ), .CK(clk), .Q(cv_next[156]), .QN() );
DFF_X2 _cv_next_reg_q_reg_157_  ( .D(_cv_next_reg_N160 ), .CK(clk), .Q(cv_next[157]), .QN() );
DFF_X2 _cv_next_reg_q_reg_158_  ( .D(_cv_next_reg_N161 ), .CK(clk), .Q(cv_next[158]), .QN() );
DFF_X2 _cv_next_reg_q_reg_159_  ( .D(_cv_next_reg_N162 ), .CK(clk), .Q(cv_next[159]), .QN() );
NAND2_X2 _add_98_2_U411  ( .A1(rnd_q[96]), .A2(cv_q[96]), .ZN(_add_98_2_n222 ) );
INV_X4 _add_98_2_U410  ( .A(_add_98_2_n343 ), .ZN(_add_98_2_n379 ) );
NAND2_X2 _add_98_2_U409  ( .A1(rnd_q[106]), .A2(cv_q[106]), .ZN(_add_98_2_n342 ) );
NAND2_X2 _add_98_2_U408  ( .A1(_add_98_2_n379 ), .A2(_add_98_2_n342 ), .ZN(_add_98_2_n359 ) );
NAND2_X2 _add_98_2_U407  ( .A1(rnd_q[104]), .A2(cv_q[104]), .ZN(_add_98_2_n52 ) );
NAND2_X2 _add_98_2_U406  ( .A1(rnd_q[97]), .A2(cv_q[97]), .ZN(_add_98_2_n375 ) );
NAND2_X2 _add_98_2_U405  ( .A1(_add_98_2_n375 ), .A2(_add_98_2_n222 ), .ZN(_add_98_2_n374 ) );
NAND2_X2 _add_98_2_U404  ( .A1(_add_98_2_n1 ), .A2(_add_98_2_n374 ), .ZN(_add_98_2_n370 ) );
NAND2_X2 _add_98_2_U403  ( .A1(cv_q[98]), .A2(rnd_q[98]), .ZN(_add_98_2_n373 ) );
INV_X4 _add_98_2_U402  ( .A(_add_98_2_n219 ), .ZN(_add_98_2_n371 ) );
NAND2_X2 _add_98_2_U401  ( .A1(rnd_q[99]), .A2(cv_q[99]), .ZN(_add_98_2_n217 ) );
INV_X4 _add_98_2_U400  ( .A(_add_98_2_n29 ), .ZN(_add_98_2_n369 ) );
NAND2_X2 _add_98_2_U399  ( .A1(rnd_q[103]), .A2(cv_q[103]), .ZN(_add_98_2_n56 ) );
NAND2_X2 _add_98_2_U398  ( .A1(rnd_q[102]), .A2(cv_q[102]), .ZN(_add_98_2_n368 ) );
NAND2_X2 _add_98_2_U397  ( .A1(rnd_q[100]), .A2(cv_q[100]), .ZN(_add_98_2_n66 ) );
NAND2_X2 _add_98_2_U396  ( .A1(rnd_q[101]), .A2(cv_q[101]), .ZN(_add_98_2_n63 ) );
NAND2_X2 _add_98_2_U395  ( .A1(_add_98_2_n66 ), .A2(_add_98_2_n63 ), .ZN(_add_98_2_n367 ) );
NAND2_X2 _add_98_2_U394  ( .A1(_add_98_2_n366 ), .A2(_add_98_2_n367 ), .ZN(_add_98_2_n365 ) );
NAND2_X2 _add_98_2_U393  ( .A1(_add_98_2_n35 ), .A2(_add_98_2_n365 ), .ZN(_add_98_2_n364 ) );
NAND2_X2 _add_98_2_U392  ( .A1(_add_98_2_n9 ), .A2(_add_98_2_n363 ), .ZN(_add_98_2_n362 ) );
XNOR2_X2 _add_98_2_U391  ( .A(_add_98_2_n359 ), .B(_add_98_2_n358 ), .ZN(N71) );
NAND2_X2 _add_98_2_U390  ( .A1(_add_98_2_n358 ), .A2(_add_98_2_n379 ), .ZN(_add_98_2_n357 ) );
NAND2_X2 _add_98_2_U389  ( .A1(_add_98_2_n357 ), .A2(_add_98_2_n342 ), .ZN(_add_98_2_n355 ) );
NAND2_X2 _add_98_2_U388  ( .A1(rnd_q[107]), .A2(cv_q[107]), .ZN(_add_98_2_n341 ) );
NAND2_X2 _add_98_2_U387  ( .A1(_add_98_2_n341 ), .A2(_add_98_2_n308 ), .ZN(_add_98_2_n356 ) );
XNOR2_X2 _add_98_2_U386  ( .A(_add_98_2_n355 ), .B(_add_98_2_n356 ), .ZN(N72) );
INV_X4 _add_98_2_U385  ( .A(_add_98_2_n43 ), .ZN(_add_98_2_n350 ) );
INV_X4 _add_98_2_U384  ( .A(_add_98_2_n46 ), .ZN(_add_98_2_n351 ) );
INV_X4 _add_98_2_U383  ( .A(_add_98_2_n308 ), .ZN(_add_98_2_n353 ) );
NAND2_X2 _add_98_2_U382  ( .A1(_add_98_2_n345 ), .A2(_add_98_2_n346 ), .ZN(_add_98_2_n337 ) );
NAND2_X2 _add_98_2_U381  ( .A1(cv_q[105]), .A2(rnd_q[105]), .ZN(_add_98_2_n344 ) );
INV_X4 _add_98_2_U380  ( .A(_add_98_2_n342 ), .ZN(_add_98_2_n339 ) );
INV_X4 _add_98_2_U379  ( .A(_add_98_2_n341 ), .ZN(_add_98_2_n340 ) );
NAND2_X2 _add_98_2_U378  ( .A1(_add_98_2_n309 ), .A2(_add_98_2_n308 ), .ZN(_add_98_2_n332 ) );
INV_X4 _add_98_2_U377  ( .A(_add_98_2_n332 ), .ZN(_add_98_2_n321 ) );
NAND2_X2 _add_98_2_U376  ( .A1(rnd_q[108]), .A2(cv_q[108]), .ZN(_add_98_2_n322 ) );
INV_X4 _add_98_2_U375  ( .A(_add_98_2_n322 ), .ZN(_add_98_2_n335 ) );
XNOR2_X2 _add_98_2_U374  ( .A(_add_98_2_n333 ), .B(_add_98_2_n334 ), .ZN(N73) );
NAND2_X2 _add_98_2_U373  ( .A1(_add_98_2_n328 ), .A2(_add_98_2_n4 ), .ZN(_add_98_2_n331 ) );
NAND2_X2 _add_98_2_U372  ( .A1(_add_98_2_n331 ), .A2(_add_98_2_n322 ), .ZN(_add_98_2_n329 ) );
NAND2_X2 _add_98_2_U371  ( .A1(rnd_q[109]), .A2(cv_q[109]), .ZN(_add_98_2_n323 ) );
NAND2_X2 _add_98_2_U370  ( .A1(_add_98_2_n323 ), .A2(_add_98_2_n6 ), .ZN(_add_98_2_n330 ) );
XNOR2_X2 _add_98_2_U369  ( .A(_add_98_2_n329 ), .B(_add_98_2_n330 ), .ZN(N74) );
NAND2_X2 _add_98_2_U368  ( .A1(rnd_q[110]), .A2(cv_q[110]), .ZN(_add_98_2_n324 ) );
NAND2_X2 _add_98_2_U367  ( .A1(_add_98_2_n11 ), .A2(_add_98_2_n324 ), .ZN(_add_98_2_n326 ) );
XNOR2_X2 _add_98_2_U366  ( .A(_add_98_2_n325 ), .B(_add_98_2_n326 ), .ZN(N75) );
INV_X4 _add_98_2_U365  ( .A(_add_98_2_n300 ), .ZN(_add_98_2_n311 ) );
INV_X4 _add_98_2_U364  ( .A(_add_98_2_n324 ), .ZN(_add_98_2_n306 ) );
NAND2_X2 _add_98_2_U363  ( .A1(_add_98_2_n322 ), .A2(_add_98_2_n323 ), .ZN(_add_98_2_n319 ) );
XNOR2_X2 _add_98_2_U362  ( .A(_add_98_2_n313 ), .B(_add_98_2_n314 ), .ZN(N76) );
NAND2_X2 _add_98_2_U361  ( .A1(rnd_q[112]), .A2(cv_q[112]), .ZN(_add_98_2_n280 ) );
NAND2_X2 _add_98_2_U360  ( .A1(_add_98_2_n280 ), .A2(_add_98_2_n282 ), .ZN(_add_98_2_n283 ) );
INV_X4 _add_98_2_U359  ( .A(_add_98_2_n133 ), .ZN(_add_98_2_n211 ) );
NAND2_X2 _add_98_2_U358  ( .A1(cv_q[109]), .A2(rnd_q[109]), .ZN(_add_98_2_n307 ) );
NAND2_X2 _add_98_2_U357  ( .A1(rnd_q[108]), .A2(cv_q[108]), .ZN(_add_98_2_n302 ) );
NAND2_X2 _add_98_2_U356  ( .A1(_add_98_2_n299 ), .A2(_add_98_2_n300 ), .ZN(_add_98_2_n132 ) );
INV_X4 _add_98_2_U355  ( .A(_add_98_2_n132 ), .ZN(_add_98_2_n210 ) );
INV_X4 _add_98_2_U354  ( .A(_add_98_2_n222 ), .ZN(_add_98_2_n298 ) );
NAND2_X2 _add_98_2_U353  ( .A1(rnd_q[97]), .A2(cv_q[97]), .ZN(_add_98_2_n138 ) );
INV_X4 _add_98_2_U352  ( .A(_add_98_2_n138 ), .ZN(_add_98_2_n260 ) );
INV_X4 _add_98_2_U351  ( .A(_add_98_2_n217 ), .ZN(_add_98_2_n77 ) );
NAND2_X2 _add_98_2_U350  ( .A1(_add_98_2_n296 ), .A2(_add_98_2_n297 ), .ZN(_add_98_2_n293 ) );
NAND2_X2 _add_98_2_U349  ( .A1(rnd_q[101]), .A2(cv_q[101]), .ZN(_add_98_2_n289 ) );
NAND2_X2 _add_98_2_U348  ( .A1(_add_98_2_n66 ), .A2(_add_98_2_n289 ), .ZN(_add_98_2_n288 ) );
NAND2_X2 _add_98_2_U347  ( .A1(_add_98_2_n227 ), .A2(_add_98_2_n288 ), .ZN(_add_98_2_n287 ) );
NAND2_X2 _add_98_2_U346  ( .A1(_add_98_2_n35 ), .A2(_add_98_2_n287 ), .ZN(_add_98_2_n285 ) );
NAND3_X2 _add_98_2_U345  ( .A1(_add_98_2_n285 ), .A2(_add_98_2_n3 ), .A3(_add_98_2_n286 ), .ZN(_add_98_2_n258 ) );
INV_X4 _add_98_2_U344  ( .A(_add_98_2_n258 ), .ZN(_add_98_2_n135 ) );
XNOR2_X2 _add_98_2_U343  ( .A(_add_98_2_n283 ), .B(_add_98_2_n88 ), .ZN(N77));
INV_X4 _add_98_2_U342  ( .A(_add_98_2_n274 ), .ZN(_add_98_2_n282 ) );
NAND2_X2 _add_98_2_U341  ( .A1(_add_98_2_n88 ), .A2(_add_98_2_n282 ), .ZN(_add_98_2_n281 ) );
NAND2_X2 _add_98_2_U340  ( .A1(_add_98_2_n280 ), .A2(_add_98_2_n281 ), .ZN(_add_98_2_n278 ) );
NAND2_X2 _add_98_2_U339  ( .A1(rnd_q[113]), .A2(cv_q[113]), .ZN(_add_98_2_n275 ) );
NAND2_X2 _add_98_2_U338  ( .A1(_add_98_2_n40 ), .A2(_add_98_2_n275 ), .ZN(_add_98_2_n279 ) );
XNOR2_X2 _add_98_2_U337  ( .A(_add_98_2_n278 ), .B(_add_98_2_n279 ), .ZN(N78) );
NAND2_X2 _add_98_2_U336  ( .A1(_add_98_2_n33 ), .A2(_add_98_2_n275 ), .ZN(_add_98_2_n265 ) );
INV_X4 _add_98_2_U335  ( .A(_add_98_2_n265 ), .ZN(_add_98_2_n271 ) );
NAND2_X2 _add_98_2_U334  ( .A1(_add_98_2_n268 ), .A2(_add_98_2_n88 ), .ZN(_add_98_2_n272 ) );
NAND2_X2 _add_98_2_U333  ( .A1(_add_98_2_n271 ), .A2(_add_98_2_n272 ), .ZN(_add_98_2_n269 ) );
NAND2_X2 _add_98_2_U332  ( .A1(rnd_q[114]), .A2(cv_q[114]), .ZN(_add_98_2_n264 ) );
NAND2_X2 _add_98_2_U331  ( .A1(_add_98_2_n264 ), .A2(_add_98_2_n266 ), .ZN(_add_98_2_n270 ) );
XNOR2_X2 _add_98_2_U330  ( .A(_add_98_2_n269 ), .B(_add_98_2_n270 ), .ZN(N79) );
INV_X4 _add_98_2_U329  ( .A(_add_98_2_n88 ), .ZN(_add_98_2_n267 ) );
NAND2_X2 _add_98_2_U328  ( .A1(_add_98_2_n268 ), .A2(_add_98_2_n266 ), .ZN(_add_98_2_n256 ) );
NAND2_X2 _add_98_2_U327  ( .A1(_add_98_2_n265 ), .A2(_add_98_2_n266 ), .ZN(_add_98_2_n263 ) );
NAND2_X2 _add_98_2_U326  ( .A1(_add_98_2_n263 ), .A2(_add_98_2_n264 ), .ZN(_add_98_2_n197 ) );
NAND2_X2 _add_98_2_U325  ( .A1(rnd_q[115]), .A2(cv_q[115]), .ZN(_add_98_2_n127 ) );
XNOR2_X2 _add_98_2_U324  ( .A(_add_98_2_n261 ), .B(_add_98_2_n23 ), .ZN(N80));
XNOR2_X2 _add_98_2_U323  ( .A(_add_98_2_n222 ), .B(_add_98_2_n259 ), .ZN(N62) );
INV_X4 _add_98_2_U322  ( .A(_add_98_2_n256 ), .ZN(_add_98_2_n255 ) );
NAND2_X2 _add_98_2_U321  ( .A1(_add_98_2_n255 ), .A2(_add_98_2_n196 ), .ZN(_add_98_2_n129 ) );
NAND2_X2 _add_98_2_U320  ( .A1(_add_98_2_n197 ), .A2(_add_98_2_n196 ), .ZN(_add_98_2_n126 ) );
NAND2_X2 _add_98_2_U319  ( .A1(_add_98_2_n126 ), .A2(_add_98_2_n127 ), .ZN(_add_98_2_n253 ) );
XNOR2_X2 _add_98_2_U318  ( .A(_add_98_2_n235 ), .B(_add_98_2_n251 ), .ZN(N81) );
NAND2_X2 _add_98_2_U317  ( .A1(rnd_q[117]), .A2(cv_q[117]), .ZN(_add_98_2_n202 ) );
INV_X4 _add_98_2_U316  ( .A(_add_98_2_n202 ), .ZN(_add_98_2_n248 ) );
XNOR2_X2 _add_98_2_U315  ( .A(_add_98_2_n246 ), .B(_add_98_2_n247 ), .ZN(N82) );
INV_X4 _add_98_2_U314  ( .A(_add_98_2_n236 ), .ZN(_add_98_2_n243 ) );
INV_X4 _add_98_2_U313  ( .A(_add_98_2_n242 ), .ZN(_add_98_2_n241 ) );
NAND2_X2 _add_98_2_U312  ( .A1(_add_98_2_n203 ), .A2(_add_98_2_n202 ), .ZN(_add_98_2_n240 ) );
NAND2_X2 _add_98_2_U311  ( .A1(rnd_q[118]), .A2(cv_q[118]), .ZN(_add_98_2_n204 ) );
XNOR2_X2 _add_98_2_U310  ( .A(_add_98_2_n238 ), .B(_add_98_2_n26 ), .ZN(N83));
NAND2_X2 _add_98_2_U309  ( .A1(_add_98_2_n203 ), .A2(_add_98_2_n202 ), .ZN(_add_98_2_n237 ) );
NAND2_X2 _add_98_2_U308  ( .A1(_add_98_2_n237 ), .A2(_add_98_2_n199 ), .ZN(_add_98_2_n234 ) );
NAND2_X2 _add_98_2_U307  ( .A1(_add_98_2_n236 ), .A2(_add_98_2_n199 ), .ZN(_add_98_2_n231 ) );
NAND2_X2 _add_98_2_U306  ( .A1(rnd_q[119]), .A2(cv_q[119]), .ZN(_add_98_2_n152 ) );
NAND2_X2 _add_98_2_U305  ( .A1(_add_98_2_n200 ), .A2(_add_98_2_n152 ), .ZN(_add_98_2_n233 ) );
XNOR2_X2 _add_98_2_U304  ( .A(_add_98_2_n232 ), .B(_add_98_2_n233 ), .ZN(N84) );
INV_X4 _add_98_2_U303  ( .A(_add_98_2_n231 ), .ZN(_add_98_2_n230 ) );
NAND2_X2 _add_98_2_U302  ( .A1(_add_98_2_n230 ), .A2(_add_98_2_n200 ), .ZN(_add_98_2_n147 ) );
NAND2_X2 _add_98_2_U301  ( .A1(rnd_q[101]), .A2(cv_q[101]), .ZN(_add_98_2_n229 ) );
NAND2_X2 _add_98_2_U300  ( .A1(_add_98_2_n66 ), .A2(_add_98_2_n229 ), .ZN(_add_98_2_n228 ) );
NAND2_X2 _add_98_2_U299  ( .A1(_add_98_2_n227 ), .A2(_add_98_2_n228 ), .ZN(_add_98_2_n226 ) );
NAND2_X2 _add_98_2_U298  ( .A1(_add_98_2_n35 ), .A2(_add_98_2_n226 ), .ZN(_add_98_2_n223 ) );
INV_X4 _add_98_2_U297  ( .A(_add_98_2_n215 ), .ZN(_add_98_2_n224 ) );
INV_X4 _add_98_2_U296  ( .A(_add_98_2_n216 ), .ZN(_add_98_2_n225 ) );
NAND4_X2 _add_98_2_U295  ( .A1(_add_98_2_n223 ), .A2(_add_98_2_n3 ), .A3(_add_98_2_n224 ), .A4(_add_98_2_n225 ), .ZN(_add_98_2_n207 ) );
NAND2_X2 _add_98_2_U294  ( .A1(rnd_q[97]), .A2(cv_q[97]), .ZN(_add_98_2_n221 ) );
NAND2_X2 _add_98_2_U293  ( .A1(_add_98_2_n221 ), .A2(_add_98_2_n222 ), .ZN(_add_98_2_n220 ) );
NAND2_X2 _add_98_2_U292  ( .A1(_add_98_2_n1 ), .A2(_add_98_2_n220 ), .ZN(_add_98_2_n218 ) );
INV_X4 _add_98_2_U291  ( .A(_add_98_2_n49 ), .ZN(_add_98_2_n214 ) );
NAND2_X2 _add_98_2_U290  ( .A1(_add_98_2_n205 ), .A2(_add_98_2_n206 ), .ZN(_add_98_2_n189 ) );
INV_X4 _add_98_2_U289  ( .A(_add_98_2_n146 ), .ZN(_add_98_2_n198 ) );
NAND2_X2 _add_98_2_U288  ( .A1(_add_98_2_n198 ), .A2(_add_98_2_n152 ), .ZN(_add_98_2_n191 ) );
INV_X4 _add_98_2_U287  ( .A(_add_98_2_n197 ), .ZN(_add_98_2_n194 ) );
INV_X4 _add_98_2_U286  ( .A(_add_98_2_n196 ), .ZN(_add_98_2_n195 ) );
NAND2_X2 _add_98_2_U285  ( .A1(_add_98_2_n189 ), .A2(_add_98_2_n190 ), .ZN(_add_98_2_n163 ) );
NAND2_X2 _add_98_2_U284  ( .A1(rnd_q[120]), .A2(cv_q[120]), .ZN(_add_98_2_n187 ) );
NAND2_X2 _add_98_2_U283  ( .A1(_add_98_2_n187 ), .A2(_add_98_2_n172 ), .ZN(_add_98_2_n188 ) );
XNOR2_X2 _add_98_2_U282  ( .A(_add_98_2_n163 ), .B(_add_98_2_n188 ), .ZN(N85) );
INV_X4 _add_98_2_U281  ( .A(_add_98_2_n181 ), .ZN(_add_98_2_n172 ) );
NAND2_X2 _add_98_2_U280  ( .A1(_add_98_2_n172 ), .A2(_add_98_2_n163 ), .ZN(_add_98_2_n186 ) );
NAND2_X2 _add_98_2_U279  ( .A1(_add_98_2_n186 ), .A2(_add_98_2_n187 ), .ZN(_add_98_2_n182 ) );
NAND2_X2 _add_98_2_U278  ( .A1(rnd_q[121]), .A2(cv_q[121]), .ZN(_add_98_2_n161 ) );
INV_X4 _add_98_2_U277  ( .A(rnd_q[121]), .ZN(_add_98_2_n184 ) );
INV_X4 _add_98_2_U276  ( .A(cv_q[121]), .ZN(_add_98_2_n185 ) );
NAND2_X2 _add_98_2_U275  ( .A1(_add_98_2_n184 ), .A2(_add_98_2_n185 ), .ZN(_add_98_2_n171 ) );
NAND2_X2 _add_98_2_U274  ( .A1(_add_98_2_n161 ), .A2(_add_98_2_n171 ), .ZN(_add_98_2_n183 ) );
XNOR2_X2 _add_98_2_U273  ( .A(_add_98_2_n182 ), .B(_add_98_2_n183 ), .ZN(N86) );
INV_X4 _add_98_2_U272  ( .A(_add_98_2_n163 ), .ZN(_add_98_2_n180 ) );
INV_X4 _add_98_2_U271  ( .A(_add_98_2_n171 ), .ZN(_add_98_2_n178 ) );
NAND2_X2 _add_98_2_U270  ( .A1(cv_q[120]), .A2(rnd_q[120]), .ZN(_add_98_2_n179 ) );
NAND2_X2 _add_98_2_U269  ( .A1(_add_98_2_n10 ), .A2(_add_98_2_n161 ), .ZN(_add_98_2_n177 ) );
INV_X4 _add_98_2_U268  ( .A(rnd_q[122]), .ZN(_add_98_2_n174 ) );
INV_X4 _add_98_2_U267  ( .A(cv_q[122]), .ZN(_add_98_2_n175 ) );
NAND2_X2 _add_98_2_U266  ( .A1(_add_98_2_n174 ), .A2(_add_98_2_n175 ), .ZN(_add_98_2_n159 ) );
NAND2_X2 _add_98_2_U265  ( .A1(rnd_q[122]), .A2(cv_q[122]), .ZN(_add_98_2_n162 ) );
XNOR2_X2 _add_98_2_U264  ( .A(_add_98_2_n173 ), .B(_add_98_2_n24 ), .ZN(N87));
NAND2_X2 _add_98_2_U263  ( .A1(_add_98_2_n30 ), .A2(_add_98_2_n163 ), .ZN(_add_98_2_n168 ) );
NAND2_X2 _add_98_2_U262  ( .A1(_add_98_2_n170 ), .A2(_add_98_2_n159 ), .ZN(_add_98_2_n169 ) );
NAND2_X2 _add_98_2_U261  ( .A1(_add_98_2_n168 ), .A2(_add_98_2_n169 ), .ZN(_add_98_2_n164 ) );
INV_X4 _add_98_2_U260  ( .A(rnd_q[123]), .ZN(_add_98_2_n166 ) );
INV_X4 _add_98_2_U259  ( .A(cv_q[123]), .ZN(_add_98_2_n167 ) );
NAND2_X2 _add_98_2_U258  ( .A1(_add_98_2_n166 ), .A2(_add_98_2_n167 ), .ZN(_add_98_2_n150 ) );
NAND2_X2 _add_98_2_U257  ( .A1(rnd_q[123]), .A2(cv_q[123]), .ZN(_add_98_2_n158 ) );
NAND2_X2 _add_98_2_U256  ( .A1(_add_98_2_n150 ), .A2(_add_98_2_n158 ), .ZN(_add_98_2_n165 ) );
XNOR2_X2 _add_98_2_U255  ( .A(_add_98_2_n164 ), .B(_add_98_2_n165 ), .ZN(N88) );
NAND2_X2 _add_98_2_U254  ( .A1(_add_98_2_n157 ), .A2(_add_98_2_n158 ), .ZN(_add_98_2_n153 ) );
INV_X4 _add_98_2_U253  ( .A(rnd_q[124]), .ZN(_add_98_2_n155 ) );
INV_X4 _add_98_2_U252  ( .A(cv_q[124]), .ZN(_add_98_2_n156 ) );
NAND2_X2 _add_98_2_U251  ( .A1(_add_98_2_n155 ), .A2(_add_98_2_n156 ), .ZN(_add_98_2_n151 ) );
NAND2_X2 _add_98_2_U250  ( .A1(rnd_q[124]), .A2(cv_q[124]), .ZN(_add_98_2_n101 ) );
XNOR2_X2 _add_98_2_U249  ( .A(_add_98_2_n154 ), .B(_add_98_2_n25 ), .ZN(N89));
INV_X4 _add_98_2_U248  ( .A(_add_98_2_n152 ), .ZN(_add_98_2_n149 ) );
INV_X4 _add_98_2_U247  ( .A(_add_98_2_n122 ), .ZN(_add_98_2_n104 ) );
INV_X4 _add_98_2_U246  ( .A(_add_98_2_n101 ), .ZN(_add_98_2_n148 ) );
INV_X4 _add_98_2_U245  ( .A(_add_98_2_n147 ), .ZN(_add_98_2_n103 ) );
INV_X4 _add_98_2_U244  ( .A(_add_98_2_n129 ), .ZN(_add_98_2_n87 ) );
NAND2_X2 _add_98_2_U243  ( .A1(_add_98_2_n126 ), .A2(_add_98_2_n127 ), .ZN(_add_98_2_n102 ) );
NAND2_X2 _add_98_2_U242  ( .A1(_add_98_2_n102 ), .A2(_add_98_2_n14 ), .ZN(_add_98_2_n145 ) );
NAND2_X2 _add_98_2_U241  ( .A1(_add_98_2_n146 ), .A2(_add_98_2_n104 ), .ZN(_add_98_2_n93 ) );
NAND4_X2 _add_98_2_U240  ( .A1(_add_98_2_n143 ), .A2(_add_98_2_n144 ), .A3(_add_98_2_n145 ), .A4(_add_98_2_n93 ), .ZN(_add_98_2_n139 ) );
NAND2_X2 _add_98_2_U239  ( .A1(rnd_q[125]), .A2(cv_q[125]), .ZN(_add_98_2_n91 ) );
INV_X4 _add_98_2_U238  ( .A(rnd_q[125]), .ZN(_add_98_2_n141 ) );
INV_X4 _add_98_2_U237  ( .A(cv_q[125]), .ZN(_add_98_2_n142 ) );
NAND2_X2 _add_98_2_U236  ( .A1(_add_98_2_n141 ), .A2(_add_98_2_n142 ), .ZN(_add_98_2_n117 ) );
NAND2_X2 _add_98_2_U235  ( .A1(_add_98_2_n91 ), .A2(_add_98_2_n117 ), .ZN(_add_98_2_n140 ) );
XNOR2_X2 _add_98_2_U234  ( .A(_add_98_2_n139 ), .B(_add_98_2_n140 ), .ZN(N90) );
XNOR2_X2 _add_98_2_U233  ( .A(_add_98_2_n80 ), .B(_add_98_2_n136 ), .ZN(N63));
INV_X4 _add_98_2_U232  ( .A(_add_98_2_n134 ), .ZN(_add_98_2_n130 ) );
NAND2_X2 _add_98_2_U231  ( .A1(_add_98_2_n132 ), .A2(_add_98_2_n133 ), .ZN(_add_98_2_n131 ) );
NAND2_X2 _add_98_2_U230  ( .A1(_add_98_2_n126 ), .A2(_add_98_2_n127 ), .ZN(_add_98_2_n125 ) );
NAND2_X2 _add_98_2_U229  ( .A1(_add_98_2_n103 ), .A2(_add_98_2_n117 ), .ZN(_add_98_2_n123 ) );
NAND2_X2 _add_98_2_U228  ( .A1(_add_98_2_n12 ), .A2(_add_98_2_n117 ), .ZN(_add_98_2_n113 ) );
INV_X4 _add_98_2_U227  ( .A(_add_98_2_n93 ), .ZN(_add_98_2_n120 ) );
NAND2_X2 _add_98_2_U226  ( .A1(_add_98_2_n120 ), .A2(_add_98_2_n117 ), .ZN(_add_98_2_n114 ) );
INV_X4 _add_98_2_U225  ( .A(_add_98_2_n91 ), .ZN(_add_98_2_n118 ) );
INV_X4 _add_98_2_U224  ( .A(_add_98_2_n117 ), .ZN(_add_98_2_n105 ) );
NAND2_X2 _add_98_2_U223  ( .A1(_add_98_2_n19 ), .A2(_add_98_2_n117 ), .ZN(_add_98_2_n116 ) );
NAND4_X2 _add_98_2_U222  ( .A1(_add_98_2_n113 ), .A2(_add_98_2_n114 ), .A3(_add_98_2_n115 ), .A4(_add_98_2_n116 ), .ZN(_add_98_2_n112 ) );
INV_X4 _add_98_2_U221  ( .A(rnd_q[126]), .ZN(_add_98_2_n109 ) );
INV_X4 _add_98_2_U220  ( .A(cv_q[126]), .ZN(_add_98_2_n110 ) );
NAND2_X2 _add_98_2_U219  ( .A1(rnd_q[126]), .A2(cv_q[126]), .ZN(_add_98_2_n100 ) );
INV_X4 _add_98_2_U218  ( .A(_add_98_2_n100 ), .ZN(_add_98_2_n108 ) );
XNOR2_X2 _add_98_2_U217  ( .A(_add_98_2_n106 ), .B(_add_98_2_n107 ), .ZN(N91) );
NAND2_X2 _add_98_2_U216  ( .A1(_add_98_2_n13 ), .A2(_add_98_2_n102 ), .ZN(_add_98_2_n83 ) );
NAND2_X2 _add_98_2_U215  ( .A1(_add_98_2_n94 ), .A2(_add_98_2_n148 ), .ZN(_add_98_2_n99 ) );
NAND2_X2 _add_98_2_U214  ( .A1(_add_98_2_n99 ), .A2(_add_98_2_n100 ), .ZN(_add_98_2_n95 ) );
NAND2_X2 _add_98_2_U213  ( .A1(_add_98_2_n12 ), .A2(_add_98_2_n94 ), .ZN(_add_98_2_n97 ) );
NAND2_X2 _add_98_2_U212  ( .A1(_add_98_2_n19 ), .A2(_add_98_2_n94 ), .ZN(_add_98_2_n98 ) );
NAND2_X2 _add_98_2_U211  ( .A1(_add_98_2_n97 ), .A2(_add_98_2_n98 ), .ZN(_add_98_2_n96 ) );
INV_X4 _add_98_2_U210  ( .A(_add_98_2_n94 ), .ZN(_add_98_2_n92 ) );
NAND4_X2 _add_98_2_U209  ( .A1(_add_98_2_n83 ), .A2(_add_98_2_n84 ), .A3(_add_98_2_n85 ), .A4(_add_98_2_n86 ), .ZN(_add_98_2_n81 ) );
XNOR2_X2 _add_98_2_U208  ( .A(rnd_q[127]), .B(cv_q[127]), .ZN(_add_98_2_n82 ) );
XNOR2_X2 _add_98_2_U207  ( .A(_add_98_2_n81 ), .B(_add_98_2_n82 ), .ZN(N92));
XNOR2_X2 _add_98_2_U206  ( .A(_add_98_2_n74 ), .B(_add_98_2_n75 ), .ZN(N64));
INV_X4 _add_98_2_U205  ( .A(_add_98_2_n66 ), .ZN(_add_98_2_n72 ) );
XNOR2_X2 _add_98_2_U204  ( .A(_add_98_2_n29 ), .B(_add_98_2_n73 ), .ZN(N65));
INV_X4 _add_98_2_U203  ( .A(_add_98_2_n63 ), .ZN(_add_98_2_n70 ) );
XNOR2_X2 _add_98_2_U202  ( .A(_add_98_2_n68 ), .B(_add_98_2_n69 ), .ZN(N66));
NAND2_X2 _add_98_2_U201  ( .A1(rnd_q[102]), .A2(cv_q[102]), .ZN(_add_98_2_n58 ) );
NAND2_X2 _add_98_2_U200  ( .A1(_add_98_2_n58 ), .A2(_add_98_2_n7 ), .ZN(_add_98_2_n61 ) );
NAND2_X2 _add_98_2_U199  ( .A1(_add_98_2_n29 ), .A2(_add_98_2_n66 ), .ZN(_add_98_2_n65 ) );
NAND2_X2 _add_98_2_U198  ( .A1(_add_98_2_n64 ), .A2(_add_98_2_n65 ), .ZN(_add_98_2_n62 ) );
NAND2_X2 _add_98_2_U197  ( .A1(_add_98_2_n62 ), .A2(_add_98_2_n63 ), .ZN(_add_98_2_n59 ) );
XNOR2_X2 _add_98_2_U196  ( .A(_add_98_2_n61 ), .B(_add_98_2_n59 ), .ZN(N67));
NAND2_X2 _add_98_2_U195  ( .A1(_add_98_2_n59 ), .A2(_add_98_2_n7 ), .ZN(_add_98_2_n57 ) );
NAND2_X2 _add_98_2_U194  ( .A1(_add_98_2_n57 ), .A2(_add_98_2_n58 ), .ZN(_add_98_2_n54 ) );
NAND2_X2 _add_98_2_U193  ( .A1(_add_98_2_n56 ), .A2(_add_98_2_n3 ), .ZN(_add_98_2_n55 ) );
XNOR2_X2 _add_98_2_U192  ( .A(_add_98_2_n54 ), .B(_add_98_2_n55 ), .ZN(N68));
INV_X4 _add_98_2_U191  ( .A(_add_98_2_n52 ), .ZN(_add_98_2_n45 ) );
XNOR2_X2 _add_98_2_U190  ( .A(_add_98_2_n50 ), .B(_add_98_2_n51 ), .ZN(N69));
XNOR2_X2 _add_98_2_U189  ( .A(_add_98_2_n41 ), .B(_add_98_2_n42 ), .ZN(N70));
NAND2_X2 _add_98_2_U188  ( .A1(_add_98_2_n258 ), .A2(_add_98_2_n134 ), .ZN(_add_98_2_n257 ) );
NOR2_X2 _add_98_2_U187  ( .A1(_add_98_2_n20 ), .A2(_add_98_2_n108 ), .ZN(_add_98_2_n107 ) );
NOR2_X2 _add_98_2_U186  ( .A1(_add_98_2_n242 ), .A2(_add_98_2_n248 ), .ZN(_add_98_2_n247 ) );
NOR2_X2 _add_98_2_U185  ( .A1(_add_98_2_n38 ), .A2(_add_98_2_n43 ), .ZN(_add_98_2_n42 ) );
NOR2_X2 _add_98_2_U184  ( .A1(_add_98_2_n70 ), .A2(_add_98_2_n67 ), .ZN(_add_98_2_n69 ) );
NOR2_X2 _add_98_2_U183  ( .A1(_add_98_2_n36 ), .A2(_add_98_2_n72 ), .ZN(_add_98_2_n73 ) );
NOR2_X2 _add_98_2_U182  ( .A1(_add_98_2_n39 ), .A2(_add_98_2_n79 ), .ZN(_add_98_2_n136 ) );
NOR2_X2 _add_98_2_U181  ( .A1(_add_98_2_n260 ), .A2(_add_98_2_n137 ), .ZN(_add_98_2_n259 ) );
AND2_X2 _add_98_2_U180  ( .A1(cv_q[104]), .A2(rnd_q[104]), .ZN(_add_98_2_n345 ) );
NOR2_X1 _add_98_2_U179  ( .A1(cv_q[105]), .A2(rnd_q[105]), .ZN(_add_98_2_n347 ) );
NOR2_X1 _add_98_2_U178  ( .A1(cv_q[106]), .A2(rnd_q[106]), .ZN(_add_98_2_n348 ) );
NOR2_X2 _add_98_2_U177  ( .A1(_add_98_2_n347 ), .A2(_add_98_2_n348 ), .ZN(_add_98_2_n346 ) );
NOR2_X2 _add_98_2_U176  ( .A1(_add_98_2_n311 ), .A2(_add_98_2_n34 ), .ZN(_add_98_2_n313 ) );
NOR2_X2 _add_98_2_U175  ( .A1(_add_98_2_n335 ), .A2(_add_98_2_n312 ), .ZN(_add_98_2_n334 ) );
NOR2_X2 _add_98_2_U174  ( .A1(_add_98_2_n76 ), .A2(_add_98_2_n77 ), .ZN(_add_98_2_n75 ) );
AND2_X2 _add_98_2_U173  ( .A1(rnd_q[98]), .A2(cv_q[98]), .ZN(_add_98_2_n39 ));
AND2_X2 _add_98_2_U172  ( .A1(rnd_q[105]), .A2(cv_q[105]), .ZN(_add_98_2_n38 ) );
AND2_X2 _add_98_2_U171  ( .A1(rnd_q[116]), .A2(cv_q[116]), .ZN(_add_98_2_n37 ) );
NOR2_X1 _add_98_2_U170  ( .A1(cv_q[113]), .A2(rnd_q[113]), .ZN(_add_98_2_n273 ) );
NOR2_X2 _add_98_2_U169  ( .A1(_add_98_2_n273 ), .A2(_add_98_2_n274 ), .ZN(_add_98_2_n268 ) );
NOR2_X1 _add_98_2_U168  ( .A1(cv_q[101]), .A2(rnd_q[101]), .ZN(_add_98_2_n290 ) );
NOR2_X1 _add_98_2_U167  ( .A1(cv_q[102]), .A2(rnd_q[102]), .ZN(_add_98_2_n291 ) );
NOR2_X2 _add_98_2_U166  ( .A1(_add_98_2_n290 ), .A2(_add_98_2_n291 ), .ZN(_add_98_2_n227 ) );
AND2_X2 _add_98_2_U165  ( .A1(_add_98_2_n56 ), .A2(_add_98_2_n368 ), .ZN(_add_98_2_n35 ) );
AND2_X2 _add_98_2_U164  ( .A1(rnd_q[111]), .A2(cv_q[111]), .ZN(_add_98_2_n34 ) );
NOR2_X1 _add_98_2_U163  ( .A1(cv_q[113]), .A2(rnd_q[113]), .ZN(_add_98_2_n276 ) );
NOR2_X2 _add_98_2_U162  ( .A1(_add_98_2_n46 ), .A2(_add_98_2_n45 ), .ZN(_add_98_2_n51 ) );
NOR2_X2 _add_98_2_U161  ( .A1(_add_98_2_n37 ), .A2(_add_98_2_n250 ), .ZN(_add_98_2_n251 ) );
NOR2_X1 _add_98_2_U160  ( .A1(cv_q[116]), .A2(rnd_q[116]), .ZN(_add_98_2_n245 ) );
NOR2_X1 _add_98_2_U159  ( .A1(cv_q[117]), .A2(rnd_q[117]), .ZN(_add_98_2_n244 ) );
NOR2_X2 _add_98_2_U158  ( .A1(_add_98_2_n244 ), .A2(_add_98_2_n245 ), .ZN(_add_98_2_n236 ) );
NOR2_X1 _add_98_2_U157  ( .A1(cv_q[101]), .A2(rnd_q[101]), .ZN(_add_98_2_n377 ) );
NOR2_X1 _add_98_2_U156  ( .A1(cv_q[117]), .A2(rnd_q[117]), .ZN(_add_98_2_n242 ) );
OR2_X2 _add_98_2_U155  ( .A1(_add_98_2_n276 ), .A2(_add_98_2_n277 ), .ZN(_add_98_2_n33 ) );
NOR2_X1 _add_98_2_U154  ( .A1(cv_q[99]), .A2(rnd_q[99]), .ZN(_add_98_2_n76 ));
NOR2_X1 _add_98_2_U153  ( .A1(cv_q[98]), .A2(rnd_q[98]), .ZN(_add_98_2_n79 ));
NOR2_X1 _add_98_2_U152  ( .A1(cv_q[97]), .A2(rnd_q[97]), .ZN(_add_98_2_n137 ) );
NAND3_X1 _add_98_2_U151  ( .A1(cv_q[116]), .A2(rnd_q[116]), .A3(_add_98_2_n241 ), .ZN(_add_98_2_n203 ) );
NOR2_X1 _add_98_2_U150  ( .A1(cv_q[116]), .A2(rnd_q[116]), .ZN(_add_98_2_n250 ) );
OR2_X2 _add_98_2_U149  ( .A1(rnd_q[119]), .A2(cv_q[119]), .ZN(_add_98_2_n200 ) );
NOR2_X1 _add_98_2_U148  ( .A1(cv_q[112]), .A2(rnd_q[112]), .ZN(_add_98_2_n274 ) );
NOR2_X1 _add_98_2_U147  ( .A1(cv_q[102]), .A2(rnd_q[102]), .ZN(_add_98_2_n60 ) );
NOR2_X2 _add_98_2_U146  ( .A1(cv_q[120]), .A2(rnd_q[120]), .ZN(_add_98_2_n181 ) );
NOR2_X1 _add_98_2_U145  ( .A1(cv_q[101]), .A2(rnd_q[101]), .ZN(_add_98_2_n67 ) );
NOR2_X2 _add_98_2_U144  ( .A1(_add_98_2_n76 ), .A2(_add_98_2_n373 ), .ZN(_add_98_2_n219 ) );
NOR2_X2 _add_98_2_U143  ( .A1(_add_98_2_n303 ), .A2(_add_98_2_n307 ), .ZN(_add_98_2_n305 ) );
NOR3_X2 _add_98_2_U142  ( .A1(_add_98_2_n302 ), .A2(_add_98_2_n303 ), .A3(_add_98_2_n304 ), .ZN(_add_98_2_n301 ) );
NOR2_X2 _add_98_2_U141  ( .A1(_add_98_2_n298 ), .A2(_add_98_2_n219 ), .ZN(_add_98_2_n296 ) );
NAND3_X2 _add_98_2_U140  ( .A1(_add_98_2_n214 ), .A2(_add_98_2_n363 ), .A3(_add_98_2_n369 ), .ZN(_add_98_2_n361 ) );
NOR2_X2 _add_98_2_U139  ( .A1(_add_98_2_n38 ), .A2(_add_98_2_n378 ), .ZN(_add_98_2_n360 ) );
NAND3_X2 _add_98_2_U138  ( .A1(_add_98_2_n360 ), .A2(_add_98_2_n361 ), .A3(_add_98_2_n362 ), .ZN(_add_98_2_n358 ) );
NAND3_X2 _add_98_2_U137  ( .A1(_add_98_2_n328 ), .A2(_add_98_2_n6 ), .A3(_add_98_2_n4 ), .ZN(_add_98_2_n327 ) );
NAND3_X2 _add_98_2_U136  ( .A1(_add_98_2_n22 ), .A2(_add_98_2_n323 ), .A3(_add_98_2_n327 ), .ZN(_add_98_2_n325 ) );
NOR2_X2 _add_98_2_U135  ( .A1(_add_98_2_n79 ), .A2(_add_98_2_n80 ), .ZN(_add_98_2_n78 ) );
NOR2_X2 _add_98_2_U134  ( .A1(_add_98_2_n78 ), .A2(_add_98_2_n39 ), .ZN(_add_98_2_n74 ) );
NOR2_X2 _add_98_2_U133  ( .A1(_add_98_2_n18 ), .A2(_add_98_2_n153 ), .ZN(_add_98_2_n154 ) );
NOR2_X2 _add_98_2_U132  ( .A1(_add_98_2_n29 ), .A2(_add_98_2_n49 ), .ZN(_add_98_2_n48 ) );
NOR2_X2 _add_98_2_U131  ( .A1(_add_98_2_n48 ), .A2(_add_98_2_n9 ), .ZN(_add_98_2_n47 ) );
NOR2_X2 _add_98_2_U130  ( .A1(_add_98_2_n46 ), .A2(_add_98_2_n47 ), .ZN(_add_98_2_n44 ) );
NOR2_X2 _add_98_2_U129  ( .A1(_add_98_2_n44 ), .A2(_add_98_2_n45 ), .ZN(_add_98_2_n41 ) );
NOR2_X2 _add_98_2_U128  ( .A1(_add_98_2_n29 ), .A2(_add_98_2_n36 ), .ZN(_add_98_2_n71 ) );
NOR2_X2 _add_98_2_U127  ( .A1(_add_98_2_n71 ), .A2(_add_98_2_n72 ), .ZN(_add_98_2_n68 ) );
NOR2_X2 _add_98_2_U126  ( .A1(_add_98_2_n60 ), .A2(_add_98_2_n67 ), .ZN(_add_98_2_n366 ) );
NOR2_X2 _add_98_2_U125  ( .A1(_add_98_2_n235 ), .A2(_add_98_2_n243 ), .ZN(_add_98_2_n239 ) );
NOR2_X2 _add_98_2_U124  ( .A1(_add_98_2_n239 ), .A2(_add_98_2_n240 ), .ZN(_add_98_2_n238 ) );
NOR2_X2 _add_98_2_U123  ( .A1(_add_98_2_n36 ), .A2(_add_98_2_n67 ), .ZN(_add_98_2_n64 ) );
NOR2_X2 _add_98_2_U122  ( .A1(_add_98_2_n20 ), .A2(_add_98_2_n91 ), .ZN(_add_98_2_n90 ) );
NAND3_X2 _add_98_2_U121  ( .A1(_add_98_2_n202 ), .A2(_add_98_2_n203 ), .A3(_add_98_2_n204 ), .ZN(_add_98_2_n201 ) );
AND2_X4 _add_98_2_U120  ( .A1(_add_98_2_n199 ), .A2(_add_98_2_n200 ), .ZN(_add_98_2_n32 ) );
AND2_X2 _add_98_2_U119  ( .A1(_add_98_2_n201 ), .A2(_add_98_2_n32 ), .ZN(_add_98_2_n146 ) );
OR2_X4 _add_98_2_U118  ( .A1(_add_98_2_n137 ), .A2(_add_98_2_n222 ), .ZN(_add_98_2_n31 ) );
AND2_X2 _add_98_2_U117  ( .A1(_add_98_2_n138 ), .A2(_add_98_2_n31 ), .ZN(_add_98_2_n80 ) );
NOR2_X2 _add_98_2_U116  ( .A1(_add_98_2_n105 ), .A2(_add_98_2_n101 ), .ZN(_add_98_2_n119 ) );
NOR2_X2 _add_98_2_U115  ( .A1(_add_98_2_n250 ), .A2(_add_98_2_n235 ), .ZN(_add_98_2_n249 ) );
NOR2_X2 _add_98_2_U114  ( .A1(_add_98_2_n249 ), .A2(_add_98_2_n37 ), .ZN(_add_98_2_n246 ) );
NOR3_X2 _add_98_2_U113  ( .A1(_add_98_2_n135 ), .A2(_add_98_2_n130 ), .A3(_add_98_2_n131 ), .ZN(_add_98_2_n128 ) );
NOR2_X2 _add_98_2_U112  ( .A1(_add_98_2_n128 ), .A2(_add_98_2_n129 ), .ZN(_add_98_2_n124 ) );
NOR2_X2 _add_98_2_U111  ( .A1(_add_98_2_n124 ), .A2(_add_98_2_n125 ), .ZN(_add_98_2_n121 ) );
NOR2_X2 _add_98_2_U110  ( .A1(_add_98_2_n312 ), .A2(_add_98_2_n15 ), .ZN(_add_98_2_n318 ) );
NOR2_X2 _add_98_2_U109  ( .A1(_add_98_2_n43 ), .A2(_add_98_2_n52 ), .ZN(_add_98_2_n378 ) );
NOR2_X2 _add_98_2_U108  ( .A1(_add_98_2_n147 ), .A2(_add_98_2_n127 ), .ZN(_add_98_2_n193 ) );
AND3_X2 _add_98_2_U107  ( .A1(_add_98_2_n171 ), .A2(_add_98_2_n159 ), .A3(_add_98_2_n172 ), .ZN(_add_98_2_n30 ) );
NAND3_X2 _add_98_2_U106  ( .A1(_add_98_2_n150 ), .A2(_add_98_2_n151 ), .A3(_add_98_2_n30 ), .ZN(_add_98_2_n122 ) );
NOR3_X2 _add_98_2_U105  ( .A1(_add_98_2_n194 ), .A2(_add_98_2_n147 ), .A3(_add_98_2_n195 ), .ZN(_add_98_2_n192 ) );
NOR2_X2 _add_98_2_U104  ( .A1(_add_98_2_n312 ), .A2(_add_98_2_n15 ), .ZN(_add_98_2_n328 ) );
NOR2_X2 _add_98_2_U103  ( .A1(_add_98_2_n46 ), .A2(_add_98_2_n43 ), .ZN(_add_98_2_n363 ) );
NAND3_X2 _add_98_2_U102  ( .A1(_add_98_2_n217 ), .A2(_add_98_2_n218 ), .A3(_add_98_2_n371 ), .ZN(_add_98_2_n212 ) );
NAND3_X2 _add_98_2_U101  ( .A1(_add_98_2_n161 ), .A2(_add_98_2_n10 ), .A3(_add_98_2_n162 ), .ZN(_add_98_2_n160 ) );
NAND3_X2 _add_98_2_U100  ( .A1(_add_98_2_n159 ), .A2(_add_98_2_n150 ), .A3(_add_98_2_n160 ), .ZN(_add_98_2_n157 ) );
NOR2_X2 _add_98_2_U99  ( .A1(_add_98_2_n36 ), .A2(_add_98_2_n377 ), .ZN(_add_98_2_n376 ) );
NAND3_X2 _add_98_2_U98  ( .A1(_add_98_2_n3 ), .A2(_add_98_2_n7 ), .A3(_add_98_2_n376 ), .ZN(_add_98_2_n49 ) );
NOR2_X2 _add_98_2_U97  ( .A1(_add_98_2_n20 ), .A2(_add_98_2_n105 ), .ZN(_add_98_2_n94 ) );
AND3_X2 _add_98_2_U96  ( .A1(_add_98_2_n371 ), .A2(_add_98_2_n217 ), .A3(_add_98_2_n370 ), .ZN(_add_98_2_n29 ) );
OR3_X4 _add_98_2_U95  ( .A1(_add_98_2_n305 ), .A2(_add_98_2_n306 ), .A3(_add_98_2_n34 ), .ZN(_add_98_2_n28 ) );
OR2_X2 _add_98_2_U94  ( .A1(_add_98_2_n28 ), .A2(_add_98_2_n301 ), .ZN(_add_98_2_n299 ) );
NOR2_X2 _add_98_2_U93  ( .A1(_add_98_2_n210 ), .A2(_add_98_2_n211 ), .ZN(_add_98_2_n209 ) );
NAND3_X2 _add_98_2_U92  ( .A1(_add_98_2_n212 ), .A2(_add_98_2_n213 ), .A3(_add_98_2_n214 ), .ZN(_add_98_2_n208 ) );
NAND3_X2 _add_98_2_U91  ( .A1(_add_98_2_n208 ), .A2(_add_98_2_n209 ), .A3(_add_98_2_n207 ), .ZN(_add_98_2_n206 ) );
NAND3_X2 _add_98_2_U90  ( .A1(_add_98_2_n234 ), .A2(_add_98_2_n204 ), .A3(_add_98_2_n17 ), .ZN(_add_98_2_n232 ) );
NOR3_X2 _add_98_2_U89  ( .A1(_add_98_2_n180 ), .A2(_add_98_2_n178 ), .A3(_add_98_2_n181 ), .ZN(_add_98_2_n176 ) );
NOR2_X2 _add_98_2_U88  ( .A1(_add_98_2_n176 ), .A2(_add_98_2_n177 ), .ZN(_add_98_2_n173 ) );
NOR2_X2 _add_98_2_U87  ( .A1(_add_98_2_n339 ), .A2(_add_98_2_n340 ), .ZN(_add_98_2_n338 ) );
NAND3_X2 _add_98_2_U86  ( .A1(_add_98_2_n337 ), .A2(_add_98_2_n16 ), .A3(_add_98_2_n338 ), .ZN(_add_98_2_n309 ) );
NAND3_X2 _add_98_2_U85  ( .A1(_add_98_2_n224 ), .A2(_add_98_2_n308 ), .A3(_add_98_2_n309 ), .ZN(_add_98_2_n133 ) );
NAND3_X2 _add_98_2_U84  ( .A1(_add_98_2_n162 ), .A2(_add_98_2_n10 ), .A3(_add_98_2_n161 ), .ZN(_add_98_2_n170 ) );
NOR2_X2 _add_98_2_U83  ( .A1(_add_98_2_n311 ), .A2(_add_98_2_n312 ), .ZN(_add_98_2_n310 ) );
NAND3_X2 _add_98_2_U82  ( .A1(_add_98_2_n6 ), .A2(_add_98_2_n11 ), .A3(_add_98_2_n310 ), .ZN(_add_98_2_n215 ) );
NOR3_X2 _add_98_2_U81  ( .A1(_add_98_2_n257 ), .A2(_add_98_2_n211 ), .A3(_add_98_2_n210 ), .ZN(_add_98_2_n254 ) );
NOR2_X2 _add_98_2_U80  ( .A1(_add_98_2_n254 ), .A2(_add_98_2_n129 ), .ZN(_add_98_2_n252 ) );
NOR2_X2 _add_98_2_U79  ( .A1(_add_98_2_n252 ), .A2(_add_98_2_n253 ), .ZN(_add_98_2_n235 ) );
NOR3_X2 _add_98_2_U78  ( .A1(_add_98_2_n219 ), .A2(_add_98_2_n77 ), .A3(_add_98_2_n1 ), .ZN(_add_98_2_n295 ) );
NOR2_X2 _add_98_2_U77  ( .A1(_add_98_2_n343 ), .A2(_add_98_2_n353 ), .ZN(_add_98_2_n352 ) );
NAND3_X2 _add_98_2_U76  ( .A1(_add_98_2_n350 ), .A2(_add_98_2_n351 ), .A3(_add_98_2_n352 ), .ZN(_add_98_2_n216 ) );
NOR2_X2 _add_98_2_U75  ( .A1(_add_98_2_n215 ), .A2(_add_98_2_n216 ), .ZN(_add_98_2_n286 ) );
NOR3_X2 _add_98_2_U74  ( .A1(_add_98_2_n191 ), .A2(_add_98_2_n192 ), .A3(_add_98_2_n193 ), .ZN(_add_98_2_n190 ) );
NOR2_X2 _add_98_2_U73  ( .A1(_add_98_2_n267 ), .A2(_add_98_2_n256 ), .ZN(_add_98_2_n262 ) );
NOR2_X2 _add_98_2_U72  ( .A1(_add_98_2_n262 ), .A2(_add_98_2_n197 ), .ZN(_add_98_2_n261 ) );
NOR2_X2 _add_98_2_U71  ( .A1(_add_98_2_n118 ), .A2(_add_98_2_n119 ), .ZN(_add_98_2_n115 ) );
NOR3_X2 _add_98_2_U70  ( .A1(_add_98_2_n121 ), .A2(_add_98_2_n122 ), .A3(_add_98_2_n123 ), .ZN(_add_98_2_n111 ) );
NOR2_X2 _add_98_2_U69  ( .A1(_add_98_2_n111 ), .A2(_add_98_2_n112 ), .ZN(_add_98_2_n106 ) );
NOR2_X2 _add_98_2_U68  ( .A1(_add_98_2_n29 ), .A2(_add_98_2_n49 ), .ZN(_add_98_2_n53 ) );
NOR2_X2 _add_98_2_U67  ( .A1(_add_98_2_n53 ), .A2(_add_98_2_n9 ), .ZN(_add_98_2_n50 ) );
NOR2_X2 _add_98_2_U66  ( .A1(_add_98_2_n129 ), .A2(_add_98_2_n147 ), .ZN(_add_98_2_n205 ) );
NOR2_X2 _add_98_2_U65  ( .A1(_add_98_2_n92 ), .A2(_add_98_2_n93 ), .ZN(_add_98_2_n89 ) );
NOR2_X2 _add_98_2_U64  ( .A1(_add_98_2_n29 ), .A2(_add_98_2_n49 ), .ZN(_add_98_2_n354 ) );
NOR2_X2 _add_98_2_U63  ( .A1(_add_98_2_n354 ), .A2(_add_98_2_n9 ), .ZN(_add_98_2_n349 ) );
NOR2_X2 _add_98_2_U62  ( .A1(_add_98_2_n349 ), .A2(_add_98_2_n216 ), .ZN(_add_98_2_n336 ) );
NOR2_X2 _add_98_2_U61  ( .A1(_add_98_2_n336 ), .A2(_add_98_2_n321 ), .ZN(_add_98_2_n333 ) );
NOR2_X2 _add_98_2_U60  ( .A1(_add_98_2_n215 ), .A2(_add_98_2_n216 ), .ZN(_add_98_2_n213 ) );
NOR2_X2 _add_98_2_U59  ( .A1(_add_98_2_n318 ), .A2(_add_98_2_n319 ), .ZN(_add_98_2_n317 ) );
NOR3_X2 _add_98_2_U58  ( .A1(_add_98_2_n316 ), .A2(_add_98_2_n317 ), .A3(_add_98_2_n21 ), .ZN(_add_98_2_n315 ) );
NOR2_X2 _add_98_2_U57  ( .A1(_add_98_2_n306 ), .A2(_add_98_2_n315 ), .ZN(_add_98_2_n314 ) );
NOR2_X2 _add_98_2_U56  ( .A1(_add_98_2_n29 ), .A2(_add_98_2_n49 ), .ZN(_add_98_2_n320 ) );
NAND3_X2 _add_98_2_U55  ( .A1(_add_98_2_n88 ), .A2(_add_98_2_n14 ), .A3(_add_98_2_n87 ), .ZN(_add_98_2_n144 ) );
NOR3_X2 _add_98_2_U54  ( .A1(_add_98_2_n19 ), .A2(_add_98_2_n12 ), .A3(_add_98_2_n148 ), .ZN(_add_98_2_n143 ) );
NOR2_X2 _add_98_2_U53  ( .A1(_add_98_2_n95 ), .A2(_add_98_2_n96 ), .ZN(_add_98_2_n84 ) );
NOR2_X2 _add_98_2_U52  ( .A1(_add_98_2_n89 ), .A2(_add_98_2_n90 ), .ZN(_add_98_2_n85 ) );
NOR4_X2 _add_98_2_U51  ( .A1(_add_98_2_n320 ), .A2(_add_98_2_n321 ), .A3(_add_98_2_n9 ), .A4(_add_98_2_n319 ), .ZN(_add_98_2_n316 ) );
NOR2_X2 _add_98_2_U50  ( .A1(_add_98_2_n260 ), .A2(_add_98_2_n77 ), .ZN(_add_98_2_n297 ) );
NOR2_X2 _add_98_2_U49  ( .A1(_add_98_2_n49 ), .A2(_add_98_2_n295 ), .ZN(_add_98_2_n294 ) );
NOR2_X2 _add_98_2_U48  ( .A1(_add_98_2_n215 ), .A2(_add_98_2_n216 ), .ZN(_add_98_2_n292 ) );
NAND3_X2 _add_98_2_U47  ( .A1(_add_98_2_n292 ), .A2(_add_98_2_n293 ), .A3(_add_98_2_n294 ), .ZN(_add_98_2_n134 ) );
NAND3_X2 _add_98_2_U46  ( .A1(_add_98_2_n87 ), .A2(_add_98_2_n88 ), .A3(_add_98_2_n13 ), .ZN(_add_98_2_n86 ) );
NOR2_X2 _add_98_2_U45  ( .A1(_add_98_2_n211 ), .A2(_add_98_2_n210 ), .ZN(_add_98_2_n284 ) );
NAND3_X2 _add_98_2_U44  ( .A1(_add_98_2_n284 ), .A2(_add_98_2_n134 ), .A3(_add_98_2_n258 ), .ZN(_add_98_2_n88 ) );
OR2_X4 _add_98_2_U43  ( .A1(rnd_q[96]), .A2(cv_q[96]), .ZN(_add_98_2_n372 ));
OR2_X1 _add_98_2_U42  ( .A1(cv_q[113]), .A2(rnd_q[113]), .ZN(_add_98_2_n40 ));
OR2_X4 _add_98_2_U41  ( .A1(rnd_q[114]), .A2(cv_q[114]), .ZN(_add_98_2_n266 ) );
NAND2_X1 _add_98_2_U40  ( .A1(cv_q[112]), .A2(rnd_q[112]), .ZN(_add_98_2_n277 ) );
OR2_X4 _add_98_2_U39  ( .A1(rnd_q[118]), .A2(cv_q[118]), .ZN(_add_98_2_n199 ) );
OR2_X4 _add_98_2_U38  ( .A1(rnd_q[115]), .A2(cv_q[115]), .ZN(_add_98_2_n196 ) );
OR2_X4 _add_98_2_U37  ( .A1(rnd_q[111]), .A2(cv_q[111]), .ZN(_add_98_2_n300 ) );
OR2_X4 _add_98_2_U36  ( .A1(rnd_q[107]), .A2(cv_q[107]), .ZN(_add_98_2_n308 ) );
NOR2_X1 _add_98_2_U35  ( .A1(cv_q[108]), .A2(rnd_q[108]), .ZN(_add_98_2_n312 ) );
NOR2_X1 _add_98_2_U34  ( .A1(rnd_q[100]), .A2(cv_q[100]), .ZN(_add_98_2_n36 ) );
NOR2_X1 _add_98_2_U33  ( .A1(cv_q[105]), .A2(rnd_q[105]), .ZN(_add_98_2_n43 ) );
NOR2_X1 _add_98_2_U32  ( .A1(cv_q[104]), .A2(rnd_q[104]), .ZN(_add_98_2_n46 ) );
NOR2_X1 _add_98_2_U31  ( .A1(cv_q[110]), .A2(rnd_q[110]), .ZN(_add_98_2_n303 ) );
NOR2_X1 _add_98_2_U30  ( .A1(cv_q[106]), .A2(rnd_q[106]), .ZN(_add_98_2_n343 ) );
NOR2_X1 _add_98_2_U29  ( .A1(cv_q[109]), .A2(rnd_q[109]), .ZN(_add_98_2_n304 ) );
AND2_X4 _add_98_2_U28  ( .A1(_add_98_2_n372 ), .A2(_add_98_2_n222 ), .ZN(N61) );
AND2_X4 _add_98_2_U27  ( .A1(_add_98_2_n199 ), .A2(_add_98_2_n204 ), .ZN(_add_98_2_n26 ) );
AND2_X4 _add_98_2_U26  ( .A1(_add_98_2_n151 ), .A2(_add_98_2_n101 ), .ZN(_add_98_2_n25 ) );
AND2_X4 _add_98_2_U25  ( .A1(_add_98_2_n159 ), .A2(_add_98_2_n162 ), .ZN(_add_98_2_n24 ) );
AND2_X4 _add_98_2_U24  ( .A1(_add_98_2_n127 ), .A2(_add_98_2_n196 ), .ZN(_add_98_2_n23 ) );
OR2_X4 _add_98_2_U23  ( .A1(_add_98_2_n304 ), .A2(_add_98_2_n322 ), .ZN(_add_98_2_n22 ) );
OR2_X4 _add_98_2_U22  ( .A1(_add_98_2_n303 ), .A2(_add_98_2_n304 ), .ZN(_add_98_2_n21 ) );
AND2_X4 _add_98_2_U21  ( .A1(_add_98_2_n109 ), .A2(_add_98_2_n110 ), .ZN(_add_98_2_n20 ) );
AND2_X4 _add_98_2_U20  ( .A1(_add_98_2_n153 ), .A2(_add_98_2_n151 ), .ZN(_add_98_2_n19 ) );
AND3_X4 _add_98_2_U19  ( .A1(_add_98_2_n30 ), .A2(_add_98_2_n150 ), .A3(_add_98_2_n163 ), .ZN(_add_98_2_n18 ) );
OR2_X4 _add_98_2_U18  ( .A1(_add_98_2_n235 ), .A2(_add_98_2_n231 ), .ZN(_add_98_2_n17 ) );
OR2_X4 _add_98_2_U17  ( .A1(_add_98_2_n343 ), .A2(_add_98_2_n344 ), .ZN(_add_98_2_n16 ) );
AND2_X4 _add_98_2_U16  ( .A1(_add_98_2_n216 ), .A2(_add_98_2_n332 ), .ZN(_add_98_2_n15 ) );
AND2_X4 _add_98_2_U15  ( .A1(_add_98_2_n103 ), .A2(_add_98_2_n104 ), .ZN(_add_98_2_n14 ) );
AND3_X4 _add_98_2_U14  ( .A1(_add_98_2_n103 ), .A2(_add_98_2_n94 ), .A3(_add_98_2_n104 ), .ZN(_add_98_2_n13 ) );
AND2_X4 _add_98_2_U13  ( .A1(_add_98_2_n149 ), .A2(_add_98_2_n104 ), .ZN(_add_98_2_n12 ) );
OR2_X4 _add_98_2_U12  ( .A1(cv_q[110]), .A2(rnd_q[110]), .ZN(_add_98_2_n11 ));
OR2_X4 _add_98_2_U11  ( .A1(_add_98_2_n178 ), .A2(_add_98_2_n179 ), .ZN(_add_98_2_n10 ) );
AND2_X4 _add_98_2_U10  ( .A1(_add_98_2_n364 ), .A2(_add_98_2_n3 ), .ZN(_add_98_2_n9 ) );
OR2_X4 _add_98_2_U9  ( .A1(cv_q[99]), .A2(rnd_q[99]), .ZN(_add_98_2_n8 ) );
OR2_X4 _add_98_2_U8  ( .A1(cv_q[102]), .A2(rnd_q[102]), .ZN(_add_98_2_n7 ));
OR2_X4 _add_98_2_U7  ( .A1(cv_q[109]), .A2(rnd_q[109]), .ZN(_add_98_2_n6 ));
OR2_X4 _add_98_2_U6  ( .A1(cv_q[98]), .A2(rnd_q[98]), .ZN(_add_98_2_n5 ) );
OR3_X4 _add_98_2_U5  ( .A1(_add_98_2_n320 ), .A2(_add_98_2_n9 ), .A3(_add_98_2_n321 ), .ZN(_add_98_2_n4 ) );
OR2_X4 _add_98_2_U4  ( .A1(cv_q[103]), .A2(rnd_q[103]), .ZN(_add_98_2_n3 ));
OR2_X4 _add_98_2_U3  ( .A1(cv_q[97]), .A2(rnd_q[97]), .ZN(_add_98_2_n2 ) );
AND3_X4 _add_98_2_U2  ( .A1(_add_98_2_n5 ), .A2(_add_98_2_n8 ), .A3(_add_98_2_n2 ), .ZN(_add_98_2_n1 ) );
NAND2_X2 _add_98_3_U413  ( .A1(rnd_q[64]), .A2(cv_q[64]), .ZN(_add_98_3_n222 ) );
INV_X4 _add_98_3_U412  ( .A(_add_98_3_n345 ), .ZN(_add_98_3_n381 ) );
NAND2_X2 _add_98_3_U411  ( .A1(rnd_q[74]), .A2(cv_q[74]), .ZN(_add_98_3_n344 ) );
NAND2_X2 _add_98_3_U410  ( .A1(_add_98_3_n381 ), .A2(_add_98_3_n344 ), .ZN(_add_98_3_n361 ) );
NAND2_X2 _add_98_3_U409  ( .A1(rnd_q[72]), .A2(cv_q[72]), .ZN(_add_98_3_n52 ) );
NAND2_X2 _add_98_3_U408  ( .A1(rnd_q[65]), .A2(cv_q[65]), .ZN(_add_98_3_n377 ) );
NAND2_X2 _add_98_3_U407  ( .A1(_add_98_3_n377 ), .A2(_add_98_3_n222 ), .ZN(_add_98_3_n376 ) );
NAND2_X2 _add_98_3_U406  ( .A1(_add_98_3_n1 ), .A2(_add_98_3_n376 ), .ZN(_add_98_3_n372 ) );
NAND2_X2 _add_98_3_U405  ( .A1(cv_q[66]), .A2(rnd_q[66]), .ZN(_add_98_3_n375 ) );
INV_X4 _add_98_3_U404  ( .A(_add_98_3_n219 ), .ZN(_add_98_3_n373 ) );
NAND2_X2 _add_98_3_U403  ( .A1(rnd_q[67]), .A2(cv_q[67]), .ZN(_add_98_3_n217 ) );
INV_X4 _add_98_3_U402  ( .A(_add_98_3_n29 ), .ZN(_add_98_3_n371 ) );
NAND2_X2 _add_98_3_U401  ( .A1(rnd_q[71]), .A2(cv_q[71]), .ZN(_add_98_3_n56 ) );
NAND2_X2 _add_98_3_U400  ( .A1(rnd_q[70]), .A2(cv_q[70]), .ZN(_add_98_3_n370 ) );
NAND2_X2 _add_98_3_U399  ( .A1(rnd_q[68]), .A2(cv_q[68]), .ZN(_add_98_3_n66 ) );
NAND2_X2 _add_98_3_U398  ( .A1(rnd_q[69]), .A2(cv_q[69]), .ZN(_add_98_3_n63 ) );
NAND2_X2 _add_98_3_U397  ( .A1(_add_98_3_n66 ), .A2(_add_98_3_n63 ), .ZN(_add_98_3_n369 ) );
NAND2_X2 _add_98_3_U396  ( .A1(_add_98_3_n368 ), .A2(_add_98_3_n369 ), .ZN(_add_98_3_n367 ) );
NAND2_X2 _add_98_3_U395  ( .A1(_add_98_3_n40 ), .A2(_add_98_3_n367 ), .ZN(_add_98_3_n366 ) );
NAND2_X2 _add_98_3_U394  ( .A1(_add_98_3_n9 ), .A2(_add_98_3_n365 ), .ZN(_add_98_3_n364 ) );
XNOR2_X2 _add_98_3_U393  ( .A(_add_98_3_n361 ), .B(_add_98_3_n360 ), .ZN(N103) );
NAND2_X2 _add_98_3_U392  ( .A1(_add_98_3_n360 ), .A2(_add_98_3_n381 ), .ZN(_add_98_3_n359 ) );
NAND2_X2 _add_98_3_U391  ( .A1(_add_98_3_n359 ), .A2(_add_98_3_n344 ), .ZN(_add_98_3_n357 ) );
NAND2_X2 _add_98_3_U390  ( .A1(rnd_q[75]), .A2(cv_q[75]), .ZN(_add_98_3_n343 ) );
NAND2_X2 _add_98_3_U389  ( .A1(_add_98_3_n343 ), .A2(_add_98_3_n310 ), .ZN(_add_98_3_n358 ) );
XNOR2_X2 _add_98_3_U388  ( .A(_add_98_3_n357 ), .B(_add_98_3_n358 ), .ZN(N104) );
INV_X4 _add_98_3_U387  ( .A(_add_98_3_n43 ), .ZN(_add_98_3_n352 ) );
INV_X4 _add_98_3_U386  ( .A(_add_98_3_n46 ), .ZN(_add_98_3_n353 ) );
INV_X4 _add_98_3_U385  ( .A(_add_98_3_n310 ), .ZN(_add_98_3_n355 ) );
NAND2_X2 _add_98_3_U384  ( .A1(_add_98_3_n347 ), .A2(_add_98_3_n348 ), .ZN(_add_98_3_n339 ) );
NAND2_X2 _add_98_3_U383  ( .A1(cv_q[73]), .A2(rnd_q[73]), .ZN(_add_98_3_n346 ) );
INV_X4 _add_98_3_U382  ( .A(_add_98_3_n344 ), .ZN(_add_98_3_n341 ) );
INV_X4 _add_98_3_U381  ( .A(_add_98_3_n343 ), .ZN(_add_98_3_n342 ) );
NAND2_X2 _add_98_3_U380  ( .A1(_add_98_3_n311 ), .A2(_add_98_3_n310 ), .ZN(_add_98_3_n334 ) );
INV_X4 _add_98_3_U379  ( .A(_add_98_3_n334 ), .ZN(_add_98_3_n323 ) );
NAND2_X2 _add_98_3_U378  ( .A1(rnd_q[76]), .A2(cv_q[76]), .ZN(_add_98_3_n324 ) );
INV_X4 _add_98_3_U377  ( .A(_add_98_3_n324 ), .ZN(_add_98_3_n337 ) );
XNOR2_X2 _add_98_3_U376  ( .A(_add_98_3_n335 ), .B(_add_98_3_n336 ), .ZN(N105) );
NAND2_X2 _add_98_3_U375  ( .A1(_add_98_3_n330 ), .A2(_add_98_3_n5 ), .ZN(_add_98_3_n333 ) );
NAND2_X2 _add_98_3_U374  ( .A1(_add_98_3_n333 ), .A2(_add_98_3_n324 ), .ZN(_add_98_3_n331 ) );
NAND2_X2 _add_98_3_U373  ( .A1(rnd_q[77]), .A2(cv_q[77]), .ZN(_add_98_3_n325 ) );
NAND2_X2 _add_98_3_U372  ( .A1(_add_98_3_n325 ), .A2(_add_98_3_n6 ), .ZN(_add_98_3_n332 ) );
XNOR2_X2 _add_98_3_U371  ( .A(_add_98_3_n331 ), .B(_add_98_3_n332 ), .ZN(N106) );
NAND2_X2 _add_98_3_U370  ( .A1(rnd_q[78]), .A2(cv_q[78]), .ZN(_add_98_3_n326 ) );
NAND2_X2 _add_98_3_U369  ( .A1(_add_98_3_n11 ), .A2(_add_98_3_n326 ), .ZN(_add_98_3_n328 ) );
XNOR2_X2 _add_98_3_U368  ( .A(_add_98_3_n327 ), .B(_add_98_3_n328 ), .ZN(N107) );
INV_X4 _add_98_3_U367  ( .A(_add_98_3_n302 ), .ZN(_add_98_3_n313 ) );
INV_X4 _add_98_3_U366  ( .A(_add_98_3_n326 ), .ZN(_add_98_3_n308 ) );
NAND2_X2 _add_98_3_U365  ( .A1(_add_98_3_n324 ), .A2(_add_98_3_n325 ), .ZN(_add_98_3_n321 ) );
XNOR2_X2 _add_98_3_U364  ( .A(_add_98_3_n315 ), .B(_add_98_3_n316 ), .ZN(N108) );
NAND2_X2 _add_98_3_U363  ( .A1(rnd_q[80]), .A2(cv_q[80]), .ZN(_add_98_3_n282 ) );
NAND2_X2 _add_98_3_U362  ( .A1(_add_98_3_n282 ), .A2(_add_98_3_n284 ), .ZN(_add_98_3_n285 ) );
INV_X4 _add_98_3_U361  ( .A(_add_98_3_n133 ), .ZN(_add_98_3_n211 ) );
NAND2_X2 _add_98_3_U360  ( .A1(cv_q[77]), .A2(rnd_q[77]), .ZN(_add_98_3_n309 ) );
NAND2_X2 _add_98_3_U359  ( .A1(rnd_q[76]), .A2(cv_q[76]), .ZN(_add_98_3_n304 ) );
NAND2_X2 _add_98_3_U358  ( .A1(_add_98_3_n301 ), .A2(_add_98_3_n302 ), .ZN(_add_98_3_n132 ) );
INV_X4 _add_98_3_U357  ( .A(_add_98_3_n132 ), .ZN(_add_98_3_n210 ) );
INV_X4 _add_98_3_U356  ( .A(_add_98_3_n222 ), .ZN(_add_98_3_n300 ) );
NAND2_X2 _add_98_3_U355  ( .A1(rnd_q[65]), .A2(cv_q[65]), .ZN(_add_98_3_n138 ) );
INV_X4 _add_98_3_U354  ( .A(_add_98_3_n138 ), .ZN(_add_98_3_n262 ) );
INV_X4 _add_98_3_U353  ( .A(_add_98_3_n217 ), .ZN(_add_98_3_n77 ) );
NAND2_X2 _add_98_3_U352  ( .A1(_add_98_3_n298 ), .A2(_add_98_3_n299 ), .ZN(_add_98_3_n295 ) );
NAND2_X2 _add_98_3_U351  ( .A1(rnd_q[69]), .A2(cv_q[69]), .ZN(_add_98_3_n291 ) );
NAND2_X2 _add_98_3_U350  ( .A1(_add_98_3_n66 ), .A2(_add_98_3_n291 ), .ZN(_add_98_3_n290 ) );
NAND2_X2 _add_98_3_U349  ( .A1(_add_98_3_n227 ), .A2(_add_98_3_n290 ), .ZN(_add_98_3_n289 ) );
NAND2_X2 _add_98_3_U348  ( .A1(_add_98_3_n40 ), .A2(_add_98_3_n289 ), .ZN(_add_98_3_n287 ) );
NAND3_X2 _add_98_3_U347  ( .A1(_add_98_3_n287 ), .A2(_add_98_3_n3 ), .A3(_add_98_3_n288 ), .ZN(_add_98_3_n260 ) );
INV_X4 _add_98_3_U346  ( .A(_add_98_3_n260 ), .ZN(_add_98_3_n135 ) );
XNOR2_X2 _add_98_3_U345  ( .A(_add_98_3_n285 ), .B(_add_98_3_n88 ), .ZN(N109) );
INV_X4 _add_98_3_U344  ( .A(_add_98_3_n276 ), .ZN(_add_98_3_n284 ) );
NAND2_X2 _add_98_3_U343  ( .A1(_add_98_3_n88 ), .A2(_add_98_3_n284 ), .ZN(_add_98_3_n283 ) );
NAND2_X2 _add_98_3_U342  ( .A1(_add_98_3_n282 ), .A2(_add_98_3_n283 ), .ZN(_add_98_3_n280 ) );
NAND2_X2 _add_98_3_U341  ( .A1(rnd_q[81]), .A2(cv_q[81]), .ZN(_add_98_3_n277 ) );
NAND2_X2 _add_98_3_U340  ( .A1(_add_98_3_n33 ), .A2(_add_98_3_n277 ), .ZN(_add_98_3_n281 ) );
XNOR2_X2 _add_98_3_U339  ( .A(_add_98_3_n280 ), .B(_add_98_3_n281 ), .ZN(N110) );
NAND2_X2 _add_98_3_U338  ( .A1(_add_98_3_n39 ), .A2(_add_98_3_n277 ), .ZN(_add_98_3_n267 ) );
INV_X4 _add_98_3_U337  ( .A(_add_98_3_n267 ), .ZN(_add_98_3_n273 ) );
NAND2_X2 _add_98_3_U336  ( .A1(_add_98_3_n270 ), .A2(_add_98_3_n88 ), .ZN(_add_98_3_n274 ) );
NAND2_X2 _add_98_3_U335  ( .A1(_add_98_3_n273 ), .A2(_add_98_3_n274 ), .ZN(_add_98_3_n271 ) );
NAND2_X2 _add_98_3_U334  ( .A1(rnd_q[82]), .A2(cv_q[82]), .ZN(_add_98_3_n266 ) );
NAND2_X2 _add_98_3_U333  ( .A1(_add_98_3_n266 ), .A2(_add_98_3_n268 ), .ZN(_add_98_3_n272 ) );
XNOR2_X2 _add_98_3_U332  ( .A(_add_98_3_n271 ), .B(_add_98_3_n272 ), .ZN(N111) );
INV_X4 _add_98_3_U331  ( .A(_add_98_3_n88 ), .ZN(_add_98_3_n269 ) );
NAND2_X2 _add_98_3_U330  ( .A1(_add_98_3_n270 ), .A2(_add_98_3_n268 ), .ZN(_add_98_3_n258 ) );
NAND2_X2 _add_98_3_U329  ( .A1(_add_98_3_n267 ), .A2(_add_98_3_n268 ), .ZN(_add_98_3_n265 ) );
NAND2_X2 _add_98_3_U328  ( .A1(_add_98_3_n265 ), .A2(_add_98_3_n266 ), .ZN(_add_98_3_n197 ) );
NAND2_X2 _add_98_3_U327  ( .A1(rnd_q[83]), .A2(cv_q[83]), .ZN(_add_98_3_n127 ) );
XNOR2_X2 _add_98_3_U326  ( .A(_add_98_3_n263 ), .B(_add_98_3_n23 ), .ZN(N112) );
XNOR2_X2 _add_98_3_U325  ( .A(_add_98_3_n222 ), .B(_add_98_3_n261 ), .ZN(N94) );
INV_X4 _add_98_3_U324  ( .A(_add_98_3_n258 ), .ZN(_add_98_3_n257 ) );
NAND2_X2 _add_98_3_U323  ( .A1(_add_98_3_n257 ), .A2(_add_98_3_n196 ), .ZN(_add_98_3_n129 ) );
NAND2_X2 _add_98_3_U322  ( .A1(_add_98_3_n197 ), .A2(_add_98_3_n196 ), .ZN(_add_98_3_n126 ) );
NAND2_X2 _add_98_3_U321  ( .A1(_add_98_3_n126 ), .A2(_add_98_3_n127 ), .ZN(_add_98_3_n255 ) );
XNOR2_X2 _add_98_3_U320  ( .A(_add_98_3_n237 ), .B(_add_98_3_n253 ), .ZN(N113) );
NAND2_X2 _add_98_3_U319  ( .A1(rnd_q[85]), .A2(cv_q[85]), .ZN(_add_98_3_n202 ) );
INV_X4 _add_98_3_U318  ( .A(_add_98_3_n202 ), .ZN(_add_98_3_n250 ) );
XNOR2_X2 _add_98_3_U317  ( .A(_add_98_3_n248 ), .B(_add_98_3_n249 ), .ZN(N114) );
INV_X4 _add_98_3_U316  ( .A(_add_98_3_n238 ), .ZN(_add_98_3_n245 ) );
INV_X4 _add_98_3_U315  ( .A(_add_98_3_n244 ), .ZN(_add_98_3_n243 ) );
NAND2_X2 _add_98_3_U314  ( .A1(_add_98_3_n203 ), .A2(_add_98_3_n202 ), .ZN(_add_98_3_n242 ) );
NAND2_X2 _add_98_3_U313  ( .A1(rnd_q[86]), .A2(cv_q[86]), .ZN(_add_98_3_n204 ) );
XNOR2_X2 _add_98_3_U312  ( .A(_add_98_3_n240 ), .B(_add_98_3_n26 ), .ZN(N115) );
NAND2_X2 _add_98_3_U311  ( .A1(_add_98_3_n203 ), .A2(_add_98_3_n202 ), .ZN(_add_98_3_n239 ) );
NAND2_X2 _add_98_3_U310  ( .A1(_add_98_3_n239 ), .A2(_add_98_3_n199 ), .ZN(_add_98_3_n236 ) );
NAND2_X2 _add_98_3_U309  ( .A1(_add_98_3_n238 ), .A2(_add_98_3_n199 ), .ZN(_add_98_3_n231 ) );
INV_X4 _add_98_3_U308  ( .A(rnd_q[87]), .ZN(_add_98_3_n234 ) );
INV_X4 _add_98_3_U307  ( .A(cv_q[87]), .ZN(_add_98_3_n235 ) );
NAND2_X2 _add_98_3_U306  ( .A1(_add_98_3_n234 ), .A2(_add_98_3_n235 ), .ZN(_add_98_3_n200 ) );
NAND2_X2 _add_98_3_U305  ( .A1(rnd_q[87]), .A2(cv_q[87]), .ZN(_add_98_3_n152 ) );
NAND2_X2 _add_98_3_U304  ( .A1(_add_98_3_n200 ), .A2(_add_98_3_n152 ), .ZN(_add_98_3_n233 ) );
XNOR2_X2 _add_98_3_U303  ( .A(_add_98_3_n232 ), .B(_add_98_3_n233 ), .ZN(N116) );
INV_X4 _add_98_3_U302  ( .A(_add_98_3_n231 ), .ZN(_add_98_3_n230 ) );
NAND2_X2 _add_98_3_U301  ( .A1(_add_98_3_n230 ), .A2(_add_98_3_n200 ), .ZN(_add_98_3_n147 ) );
NAND2_X2 _add_98_3_U300  ( .A1(rnd_q[69]), .A2(cv_q[69]), .ZN(_add_98_3_n229 ) );
NAND2_X2 _add_98_3_U299  ( .A1(_add_98_3_n66 ), .A2(_add_98_3_n229 ), .ZN(_add_98_3_n228 ) );
NAND2_X2 _add_98_3_U298  ( .A1(_add_98_3_n227 ), .A2(_add_98_3_n228 ), .ZN(_add_98_3_n226 ) );
NAND2_X2 _add_98_3_U297  ( .A1(_add_98_3_n40 ), .A2(_add_98_3_n226 ), .ZN(_add_98_3_n223 ) );
INV_X4 _add_98_3_U296  ( .A(_add_98_3_n215 ), .ZN(_add_98_3_n224 ) );
INV_X4 _add_98_3_U295  ( .A(_add_98_3_n216 ), .ZN(_add_98_3_n225 ) );
NAND4_X2 _add_98_3_U294  ( .A1(_add_98_3_n223 ), .A2(_add_98_3_n3 ), .A3(_add_98_3_n224 ), .A4(_add_98_3_n225 ), .ZN(_add_98_3_n207 ) );
NAND2_X2 _add_98_3_U293  ( .A1(rnd_q[65]), .A2(cv_q[65]), .ZN(_add_98_3_n221 ) );
NAND2_X2 _add_98_3_U292  ( .A1(_add_98_3_n221 ), .A2(_add_98_3_n222 ), .ZN(_add_98_3_n220 ) );
NAND2_X2 _add_98_3_U291  ( .A1(_add_98_3_n1 ), .A2(_add_98_3_n220 ), .ZN(_add_98_3_n218 ) );
INV_X4 _add_98_3_U290  ( .A(_add_98_3_n49 ), .ZN(_add_98_3_n214 ) );
NAND2_X2 _add_98_3_U289  ( .A1(_add_98_3_n205 ), .A2(_add_98_3_n206 ), .ZN(_add_98_3_n189 ) );
INV_X4 _add_98_3_U288  ( .A(_add_98_3_n146 ), .ZN(_add_98_3_n198 ) );
NAND2_X2 _add_98_3_U287  ( .A1(_add_98_3_n198 ), .A2(_add_98_3_n152 ), .ZN(_add_98_3_n191 ) );
INV_X4 _add_98_3_U286  ( .A(_add_98_3_n197 ), .ZN(_add_98_3_n194 ) );
INV_X4 _add_98_3_U285  ( .A(_add_98_3_n196 ), .ZN(_add_98_3_n195 ) );
NAND2_X2 _add_98_3_U284  ( .A1(_add_98_3_n189 ), .A2(_add_98_3_n190 ), .ZN(_add_98_3_n163 ) );
NAND2_X2 _add_98_3_U283  ( .A1(rnd_q[88]), .A2(cv_q[88]), .ZN(_add_98_3_n187 ) );
NAND2_X2 _add_98_3_U282  ( .A1(_add_98_3_n187 ), .A2(_add_98_3_n172 ), .ZN(_add_98_3_n188 ) );
XNOR2_X2 _add_98_3_U281  ( .A(_add_98_3_n163 ), .B(_add_98_3_n188 ), .ZN(N117) );
INV_X4 _add_98_3_U280  ( .A(_add_98_3_n181 ), .ZN(_add_98_3_n172 ) );
NAND2_X2 _add_98_3_U279  ( .A1(_add_98_3_n172 ), .A2(_add_98_3_n163 ), .ZN(_add_98_3_n186 ) );
NAND2_X2 _add_98_3_U278  ( .A1(_add_98_3_n186 ), .A2(_add_98_3_n187 ), .ZN(_add_98_3_n182 ) );
NAND2_X2 _add_98_3_U277  ( .A1(rnd_q[89]), .A2(cv_q[89]), .ZN(_add_98_3_n161 ) );
INV_X4 _add_98_3_U276  ( .A(rnd_q[89]), .ZN(_add_98_3_n184 ) );
INV_X4 _add_98_3_U275  ( .A(cv_q[89]), .ZN(_add_98_3_n185 ) );
NAND2_X2 _add_98_3_U274  ( .A1(_add_98_3_n184 ), .A2(_add_98_3_n185 ), .ZN(_add_98_3_n171 ) );
NAND2_X2 _add_98_3_U273  ( .A1(_add_98_3_n161 ), .A2(_add_98_3_n171 ), .ZN(_add_98_3_n183 ) );
XNOR2_X2 _add_98_3_U272  ( .A(_add_98_3_n182 ), .B(_add_98_3_n183 ), .ZN(N118) );
INV_X4 _add_98_3_U271  ( .A(_add_98_3_n163 ), .ZN(_add_98_3_n180 ) );
INV_X4 _add_98_3_U270  ( .A(_add_98_3_n171 ), .ZN(_add_98_3_n178 ) );
NAND2_X2 _add_98_3_U269  ( .A1(cv_q[88]), .A2(rnd_q[88]), .ZN(_add_98_3_n179 ) );
NAND2_X2 _add_98_3_U268  ( .A1(_add_98_3_n10 ), .A2(_add_98_3_n161 ), .ZN(_add_98_3_n177 ) );
INV_X4 _add_98_3_U267  ( .A(rnd_q[90]), .ZN(_add_98_3_n174 ) );
INV_X4 _add_98_3_U266  ( .A(cv_q[90]), .ZN(_add_98_3_n175 ) );
NAND2_X2 _add_98_3_U265  ( .A1(_add_98_3_n174 ), .A2(_add_98_3_n175 ), .ZN(_add_98_3_n159 ) );
NAND2_X2 _add_98_3_U264  ( .A1(rnd_q[90]), .A2(cv_q[90]), .ZN(_add_98_3_n162 ) );
XNOR2_X2 _add_98_3_U263  ( .A(_add_98_3_n173 ), .B(_add_98_3_n24 ), .ZN(N119) );
NAND2_X2 _add_98_3_U262  ( .A1(_add_98_3_n30 ), .A2(_add_98_3_n163 ), .ZN(_add_98_3_n168 ) );
NAND2_X2 _add_98_3_U261  ( .A1(_add_98_3_n170 ), .A2(_add_98_3_n159 ), .ZN(_add_98_3_n169 ) );
NAND2_X2 _add_98_3_U260  ( .A1(_add_98_3_n168 ), .A2(_add_98_3_n169 ), .ZN(_add_98_3_n164 ) );
INV_X4 _add_98_3_U259  ( .A(rnd_q[91]), .ZN(_add_98_3_n166 ) );
INV_X4 _add_98_3_U258  ( .A(cv_q[91]), .ZN(_add_98_3_n167 ) );
NAND2_X2 _add_98_3_U257  ( .A1(_add_98_3_n166 ), .A2(_add_98_3_n167 ), .ZN(_add_98_3_n150 ) );
NAND2_X2 _add_98_3_U256  ( .A1(rnd_q[91]), .A2(cv_q[91]), .ZN(_add_98_3_n158 ) );
NAND2_X2 _add_98_3_U255  ( .A1(_add_98_3_n150 ), .A2(_add_98_3_n158 ), .ZN(_add_98_3_n165 ) );
XNOR2_X2 _add_98_3_U254  ( .A(_add_98_3_n164 ), .B(_add_98_3_n165 ), .ZN(N120) );
NAND2_X2 _add_98_3_U253  ( .A1(_add_98_3_n157 ), .A2(_add_98_3_n158 ), .ZN(_add_98_3_n153 ) );
INV_X4 _add_98_3_U252  ( .A(rnd_q[92]), .ZN(_add_98_3_n155 ) );
INV_X4 _add_98_3_U251  ( .A(cv_q[92]), .ZN(_add_98_3_n156 ) );
NAND2_X2 _add_98_3_U250  ( .A1(_add_98_3_n155 ), .A2(_add_98_3_n156 ), .ZN(_add_98_3_n151 ) );
NAND2_X2 _add_98_3_U249  ( .A1(rnd_q[92]), .A2(cv_q[92]), .ZN(_add_98_3_n101 ) );
XNOR2_X2 _add_98_3_U248  ( .A(_add_98_3_n154 ), .B(_add_98_3_n25 ), .ZN(N121) );
INV_X4 _add_98_3_U247  ( .A(_add_98_3_n152 ), .ZN(_add_98_3_n149 ) );
INV_X4 _add_98_3_U246  ( .A(_add_98_3_n122 ), .ZN(_add_98_3_n104 ) );
INV_X4 _add_98_3_U245  ( .A(_add_98_3_n101 ), .ZN(_add_98_3_n148 ) );
INV_X4 _add_98_3_U244  ( .A(_add_98_3_n147 ), .ZN(_add_98_3_n103 ) );
INV_X4 _add_98_3_U243  ( .A(_add_98_3_n129 ), .ZN(_add_98_3_n87 ) );
NAND2_X2 _add_98_3_U242  ( .A1(_add_98_3_n126 ), .A2(_add_98_3_n127 ), .ZN(_add_98_3_n102 ) );
NAND2_X2 _add_98_3_U241  ( .A1(_add_98_3_n102 ), .A2(_add_98_3_n14 ), .ZN(_add_98_3_n145 ) );
NAND2_X2 _add_98_3_U240  ( .A1(_add_98_3_n146 ), .A2(_add_98_3_n104 ), .ZN(_add_98_3_n93 ) );
NAND4_X2 _add_98_3_U239  ( .A1(_add_98_3_n143 ), .A2(_add_98_3_n144 ), .A3(_add_98_3_n145 ), .A4(_add_98_3_n93 ), .ZN(_add_98_3_n139 ) );
NAND2_X2 _add_98_3_U238  ( .A1(rnd_q[93]), .A2(cv_q[93]), .ZN(_add_98_3_n91 ) );
INV_X4 _add_98_3_U237  ( .A(rnd_q[93]), .ZN(_add_98_3_n141 ) );
INV_X4 _add_98_3_U236  ( .A(cv_q[93]), .ZN(_add_98_3_n142 ) );
NAND2_X2 _add_98_3_U235  ( .A1(_add_98_3_n141 ), .A2(_add_98_3_n142 ), .ZN(_add_98_3_n117 ) );
NAND2_X2 _add_98_3_U234  ( .A1(_add_98_3_n91 ), .A2(_add_98_3_n117 ), .ZN(_add_98_3_n140 ) );
XNOR2_X2 _add_98_3_U233  ( .A(_add_98_3_n139 ), .B(_add_98_3_n140 ), .ZN(N122) );
XNOR2_X2 _add_98_3_U232  ( .A(_add_98_3_n80 ), .B(_add_98_3_n136 ), .ZN(N95));
INV_X4 _add_98_3_U231  ( .A(_add_98_3_n134 ), .ZN(_add_98_3_n130 ) );
NAND2_X2 _add_98_3_U230  ( .A1(_add_98_3_n132 ), .A2(_add_98_3_n133 ), .ZN(_add_98_3_n131 ) );
NAND2_X2 _add_98_3_U229  ( .A1(_add_98_3_n126 ), .A2(_add_98_3_n127 ), .ZN(_add_98_3_n125 ) );
NAND2_X2 _add_98_3_U228  ( .A1(_add_98_3_n103 ), .A2(_add_98_3_n117 ), .ZN(_add_98_3_n123 ) );
NAND2_X2 _add_98_3_U227  ( .A1(_add_98_3_n12 ), .A2(_add_98_3_n117 ), .ZN(_add_98_3_n113 ) );
INV_X4 _add_98_3_U226  ( .A(_add_98_3_n93 ), .ZN(_add_98_3_n120 ) );
NAND2_X2 _add_98_3_U225  ( .A1(_add_98_3_n120 ), .A2(_add_98_3_n117 ), .ZN(_add_98_3_n114 ) );
INV_X4 _add_98_3_U224  ( .A(_add_98_3_n91 ), .ZN(_add_98_3_n118 ) );
INV_X4 _add_98_3_U223  ( .A(_add_98_3_n117 ), .ZN(_add_98_3_n105 ) );
NAND2_X2 _add_98_3_U222  ( .A1(_add_98_3_n19 ), .A2(_add_98_3_n117 ), .ZN(_add_98_3_n116 ) );
NAND4_X2 _add_98_3_U221  ( .A1(_add_98_3_n113 ), .A2(_add_98_3_n114 ), .A3(_add_98_3_n115 ), .A4(_add_98_3_n116 ), .ZN(_add_98_3_n112 ) );
INV_X4 _add_98_3_U220  ( .A(rnd_q[94]), .ZN(_add_98_3_n109 ) );
INV_X4 _add_98_3_U219  ( .A(cv_q[94]), .ZN(_add_98_3_n110 ) );
NAND2_X2 _add_98_3_U218  ( .A1(rnd_q[94]), .A2(cv_q[94]), .ZN(_add_98_3_n100 ) );
INV_X4 _add_98_3_U217  ( .A(_add_98_3_n100 ), .ZN(_add_98_3_n108 ) );
XNOR2_X2 _add_98_3_U216  ( .A(_add_98_3_n106 ), .B(_add_98_3_n107 ), .ZN(N123) );
NAND2_X2 _add_98_3_U215  ( .A1(_add_98_3_n13 ), .A2(_add_98_3_n102 ), .ZN(_add_98_3_n83 ) );
NAND2_X2 _add_98_3_U214  ( .A1(_add_98_3_n94 ), .A2(_add_98_3_n148 ), .ZN(_add_98_3_n99 ) );
NAND2_X2 _add_98_3_U213  ( .A1(_add_98_3_n99 ), .A2(_add_98_3_n100 ), .ZN(_add_98_3_n95 ) );
NAND2_X2 _add_98_3_U212  ( .A1(_add_98_3_n12 ), .A2(_add_98_3_n94 ), .ZN(_add_98_3_n97 ) );
NAND2_X2 _add_98_3_U211  ( .A1(_add_98_3_n19 ), .A2(_add_98_3_n94 ), .ZN(_add_98_3_n98 ) );
NAND2_X2 _add_98_3_U210  ( .A1(_add_98_3_n97 ), .A2(_add_98_3_n98 ), .ZN(_add_98_3_n96 ) );
INV_X4 _add_98_3_U209  ( .A(_add_98_3_n94 ), .ZN(_add_98_3_n92 ) );
NAND4_X2 _add_98_3_U208  ( .A1(_add_98_3_n83 ), .A2(_add_98_3_n84 ), .A3(_add_98_3_n85 ), .A4(_add_98_3_n86 ), .ZN(_add_98_3_n81 ) );
XNOR2_X2 _add_98_3_U207  ( .A(rnd_q[95]), .B(cv_q[95]), .ZN(_add_98_3_n82 ));
XNOR2_X2 _add_98_3_U206  ( .A(_add_98_3_n81 ), .B(_add_98_3_n82 ), .ZN(N124));
XNOR2_X2 _add_98_3_U205  ( .A(_add_98_3_n74 ), .B(_add_98_3_n75 ), .ZN(N96));
INV_X4 _add_98_3_U204  ( .A(_add_98_3_n66 ), .ZN(_add_98_3_n72 ) );
XNOR2_X2 _add_98_3_U203  ( .A(_add_98_3_n29 ), .B(_add_98_3_n73 ), .ZN(N97));
INV_X4 _add_98_3_U202  ( .A(_add_98_3_n63 ), .ZN(_add_98_3_n70 ) );
XNOR2_X2 _add_98_3_U201  ( .A(_add_98_3_n68 ), .B(_add_98_3_n69 ), .ZN(N98));
NAND2_X2 _add_98_3_U200  ( .A1(rnd_q[70]), .A2(cv_q[70]), .ZN(_add_98_3_n58 ) );
NAND2_X2 _add_98_3_U199  ( .A1(_add_98_3_n58 ), .A2(_add_98_3_n7 ), .ZN(_add_98_3_n61 ) );
NAND2_X2 _add_98_3_U198  ( .A1(_add_98_3_n29 ), .A2(_add_98_3_n66 ), .ZN(_add_98_3_n65 ) );
NAND2_X2 _add_98_3_U197  ( .A1(_add_98_3_n64 ), .A2(_add_98_3_n65 ), .ZN(_add_98_3_n62 ) );
NAND2_X2 _add_98_3_U196  ( .A1(_add_98_3_n62 ), .A2(_add_98_3_n63 ), .ZN(_add_98_3_n59 ) );
XNOR2_X2 _add_98_3_U195  ( .A(_add_98_3_n61 ), .B(_add_98_3_n59 ), .ZN(N99));
NAND2_X2 _add_98_3_U194  ( .A1(_add_98_3_n59 ), .A2(_add_98_3_n7 ), .ZN(_add_98_3_n57 ) );
NAND2_X2 _add_98_3_U193  ( .A1(_add_98_3_n57 ), .A2(_add_98_3_n58 ), .ZN(_add_98_3_n54 ) );
NAND2_X2 _add_98_3_U192  ( .A1(_add_98_3_n56 ), .A2(_add_98_3_n3 ), .ZN(_add_98_3_n55 ) );
XNOR2_X2 _add_98_3_U191  ( .A(_add_98_3_n54 ), .B(_add_98_3_n55 ), .ZN(N100));
INV_X4 _add_98_3_U190  ( .A(_add_98_3_n52 ), .ZN(_add_98_3_n45 ) );
XNOR2_X2 _add_98_3_U189  ( .A(_add_98_3_n50 ), .B(_add_98_3_n51 ), .ZN(N101));
XNOR2_X2 _add_98_3_U188  ( .A(_add_98_3_n41 ), .B(_add_98_3_n42 ), .ZN(N102));
NAND2_X2 _add_98_3_U187  ( .A1(_add_98_3_n260 ), .A2(_add_98_3_n134 ), .ZN(_add_98_3_n259 ) );
NOR2_X2 _add_98_3_U186  ( .A1(_add_98_3_n313 ), .A2(_add_98_3_n38 ), .ZN(_add_98_3_n315 ) );
NOR2_X2 _add_98_3_U185  ( .A1(_add_98_3_n70 ), .A2(_add_98_3_n67 ), .ZN(_add_98_3_n69 ) );
NOR2_X2 _add_98_3_U184  ( .A1(_add_98_3_n34 ), .A2(_add_98_3_n72 ), .ZN(_add_98_3_n73 ) );
NOR2_X2 _add_98_3_U183  ( .A1(_add_98_3_n36 ), .A2(_add_98_3_n79 ), .ZN(_add_98_3_n136 ) );
AND2_X2 _add_98_3_U182  ( .A1(cv_q[72]), .A2(rnd_q[72]), .ZN(_add_98_3_n347 ) );
AND2_X2 _add_98_3_U181  ( .A1(_add_98_3_n56 ), .A2(_add_98_3_n370 ), .ZN(_add_98_3_n40 ) );
NOR2_X2 _add_98_3_U180  ( .A1(_add_98_3_n20 ), .A2(_add_98_3_n108 ), .ZN(_add_98_3_n107 ) );
NOR2_X2 _add_98_3_U179  ( .A1(_add_98_3_n244 ), .A2(_add_98_3_n250 ), .ZN(_add_98_3_n249 ) );
NOR2_X2 _add_98_3_U178  ( .A1(_add_98_3_n46 ), .A2(_add_98_3_n45 ), .ZN(_add_98_3_n51 ) );
NOR2_X2 _add_98_3_U177  ( .A1(_add_98_3_n76 ), .A2(_add_98_3_n77 ), .ZN(_add_98_3_n75 ) );
NOR2_X2 _add_98_3_U176  ( .A1(_add_98_3_n262 ), .A2(_add_98_3_n137 ), .ZN(_add_98_3_n261 ) );
OR2_X2 _add_98_3_U175  ( .A1(_add_98_3_n278 ), .A2(_add_98_3_n279 ), .ZN(_add_98_3_n39 ) );
AND2_X2 _add_98_3_U174  ( .A1(rnd_q[79]), .A2(cv_q[79]), .ZN(_add_98_3_n38 ));
AND2_X2 _add_98_3_U173  ( .A1(rnd_q[73]), .A2(cv_q[73]), .ZN(_add_98_3_n37 ));
AND2_X2 _add_98_3_U172  ( .A1(rnd_q[66]), .A2(cv_q[66]), .ZN(_add_98_3_n36 ));
AND2_X2 _add_98_3_U171  ( .A1(rnd_q[84]), .A2(cv_q[84]), .ZN(_add_98_3_n35 ));
NOR2_X2 _add_98_3_U170  ( .A1(_add_98_3_n275 ), .A2(_add_98_3_n276 ), .ZN(_add_98_3_n270 ) );
NOR2_X1 _add_98_3_U169  ( .A1(cv_q[73]), .A2(rnd_q[73]), .ZN(_add_98_3_n349 ) );
NOR2_X1 _add_98_3_U168  ( .A1(cv_q[74]), .A2(rnd_q[74]), .ZN(_add_98_3_n350 ) );
NOR2_X2 _add_98_3_U167  ( .A1(_add_98_3_n349 ), .A2(_add_98_3_n350 ), .ZN(_add_98_3_n348 ) );
NOR2_X2 _add_98_3_U166  ( .A1(_add_98_3_n246 ), .A2(_add_98_3_n247 ), .ZN(_add_98_3_n238 ) );
NOR2_X2 _add_98_3_U165  ( .A1(_add_98_3_n35 ), .A2(_add_98_3_n252 ), .ZN(_add_98_3_n253 ) );
NOR2_X2 _add_98_3_U164  ( .A1(_add_98_3_n337 ), .A2(_add_98_3_n314 ), .ZN(_add_98_3_n336 ) );
NOR2_X2 _add_98_3_U163  ( .A1(_add_98_3_n37 ), .A2(_add_98_3_n43 ), .ZN(_add_98_3_n42 ) );
NOR2_X1 _add_98_3_U162  ( .A1(cv_q[69]), .A2(rnd_q[69]), .ZN(_add_98_3_n292 ) );
NOR2_X1 _add_98_3_U161  ( .A1(cv_q[70]), .A2(rnd_q[70]), .ZN(_add_98_3_n293 ) );
NOR2_X2 _add_98_3_U160  ( .A1(_add_98_3_n292 ), .A2(_add_98_3_n293 ), .ZN(_add_98_3_n227 ) );
NOR2_X1 _add_98_3_U159  ( .A1(cv_q[69]), .A2(rnd_q[69]), .ZN(_add_98_3_n379 ) );
NOR2_X1 _add_98_3_U158  ( .A1(cv_q[67]), .A2(rnd_q[67]), .ZN(_add_98_3_n76 ));
NOR2_X1 _add_98_3_U157  ( .A1(cv_q[66]), .A2(rnd_q[66]), .ZN(_add_98_3_n79 ));
NOR2_X2 _add_98_3_U156  ( .A1(cv_q[88]), .A2(rnd_q[88]), .ZN(_add_98_3_n181 ) );
NOR2_X1 _add_98_3_U155  ( .A1(cv_q[70]), .A2(rnd_q[70]), .ZN(_add_98_3_n60 ));
NOR2_X1 _add_98_3_U154  ( .A1(cv_q[69]), .A2(rnd_q[69]), .ZN(_add_98_3_n67 ));
NOR2_X2 _add_98_3_U153  ( .A1(_add_98_3_n76 ), .A2(_add_98_3_n375 ), .ZN(_add_98_3_n219 ) );
NOR2_X2 _add_98_3_U152  ( .A1(_add_98_3_n305 ), .A2(_add_98_3_n309 ), .ZN(_add_98_3_n307 ) );
NOR3_X2 _add_98_3_U151  ( .A1(_add_98_3_n304 ), .A2(_add_98_3_n305 ), .A3(_add_98_3_n306 ), .ZN(_add_98_3_n303 ) );
NAND3_X2 _add_98_3_U150  ( .A1(_add_98_3_n202 ), .A2(_add_98_3_n203 ), .A3(_add_98_3_n204 ), .ZN(_add_98_3_n201 ) );
AND2_X4 _add_98_3_U149  ( .A1(_add_98_3_n199 ), .A2(_add_98_3_n200 ), .ZN(_add_98_3_n32 ) );
AND2_X2 _add_98_3_U148  ( .A1(_add_98_3_n201 ), .A2(_add_98_3_n32 ), .ZN(_add_98_3_n146 ) );
NOR2_X2 _add_98_3_U147  ( .A1(_add_98_3_n300 ), .A2(_add_98_3_n219 ), .ZN(_add_98_3_n298 ) );
NAND3_X2 _add_98_3_U146  ( .A1(_add_98_3_n214 ), .A2(_add_98_3_n365 ), .A3(_add_98_3_n371 ), .ZN(_add_98_3_n363 ) );
NOR2_X2 _add_98_3_U145  ( .A1(_add_98_3_n37 ), .A2(_add_98_3_n380 ), .ZN(_add_98_3_n362 ) );
NAND3_X2 _add_98_3_U144  ( .A1(_add_98_3_n362 ), .A2(_add_98_3_n363 ), .A3(_add_98_3_n364 ), .ZN(_add_98_3_n360 ) );
NAND3_X2 _add_98_3_U143  ( .A1(_add_98_3_n330 ), .A2(_add_98_3_n6 ), .A3(_add_98_3_n5 ), .ZN(_add_98_3_n329 ) );
NAND3_X2 _add_98_3_U142  ( .A1(_add_98_3_n22 ), .A2(_add_98_3_n325 ), .A3(_add_98_3_n329 ), .ZN(_add_98_3_n327 ) );
NOR2_X2 _add_98_3_U141  ( .A1(_add_98_3_n79 ), .A2(_add_98_3_n80 ), .ZN(_add_98_3_n78 ) );
NOR2_X2 _add_98_3_U140  ( .A1(_add_98_3_n78 ), .A2(_add_98_3_n36 ), .ZN(_add_98_3_n74 ) );
NOR2_X2 _add_98_3_U139  ( .A1(_add_98_3_n18 ), .A2(_add_98_3_n153 ), .ZN(_add_98_3_n154 ) );
NOR2_X2 _add_98_3_U138  ( .A1(_add_98_3_n237 ), .A2(_add_98_3_n245 ), .ZN(_add_98_3_n241 ) );
NOR2_X2 _add_98_3_U137  ( .A1(_add_98_3_n241 ), .A2(_add_98_3_n242 ), .ZN(_add_98_3_n240 ) );
NOR2_X2 _add_98_3_U136  ( .A1(_add_98_3_n29 ), .A2(_add_98_3_n49 ), .ZN(_add_98_3_n48 ) );
NOR2_X2 _add_98_3_U135  ( .A1(_add_98_3_n48 ), .A2(_add_98_3_n9 ), .ZN(_add_98_3_n47 ) );
NOR2_X2 _add_98_3_U134  ( .A1(_add_98_3_n46 ), .A2(_add_98_3_n47 ), .ZN(_add_98_3_n44 ) );
NOR2_X2 _add_98_3_U133  ( .A1(_add_98_3_n44 ), .A2(_add_98_3_n45 ), .ZN(_add_98_3_n41 ) );
NOR2_X2 _add_98_3_U132  ( .A1(_add_98_3_n29 ), .A2(_add_98_3_n34 ), .ZN(_add_98_3_n71 ) );
NOR2_X2 _add_98_3_U131  ( .A1(_add_98_3_n71 ), .A2(_add_98_3_n72 ), .ZN(_add_98_3_n68 ) );
NOR3_X2 _add_98_3_U130  ( .A1(_add_98_3_n180 ), .A2(_add_98_3_n178 ), .A3(_add_98_3_n181 ), .ZN(_add_98_3_n176 ) );
NOR2_X2 _add_98_3_U129  ( .A1(_add_98_3_n176 ), .A2(_add_98_3_n177 ), .ZN(_add_98_3_n173 ) );
NOR2_X2 _add_98_3_U128  ( .A1(_add_98_3_n60 ), .A2(_add_98_3_n67 ), .ZN(_add_98_3_n368 ) );
NOR2_X2 _add_98_3_U127  ( .A1(_add_98_3_n341 ), .A2(_add_98_3_n342 ), .ZN(_add_98_3_n340 ) );
NAND3_X2 _add_98_3_U126  ( .A1(_add_98_3_n339 ), .A2(_add_98_3_n16 ), .A3(_add_98_3_n340 ), .ZN(_add_98_3_n311 ) );
NOR2_X2 _add_98_3_U125  ( .A1(_add_98_3_n34 ), .A2(_add_98_3_n67 ), .ZN(_add_98_3_n64 ) );
NOR2_X2 _add_98_3_U124  ( .A1(_add_98_3_n20 ), .A2(_add_98_3_n91 ), .ZN(_add_98_3_n90 ) );
NOR2_X2 _add_98_3_U123  ( .A1(_add_98_3_n105 ), .A2(_add_98_3_n101 ), .ZN(_add_98_3_n119 ) );
OR2_X4 _add_98_3_U122  ( .A1(_add_98_3_n137 ), .A2(_add_98_3_n222 ), .ZN(_add_98_3_n31 ) );
AND2_X2 _add_98_3_U121  ( .A1(_add_98_3_n138 ), .A2(_add_98_3_n31 ), .ZN(_add_98_3_n80 ) );
NOR2_X2 _add_98_3_U120  ( .A1(_add_98_3_n252 ), .A2(_add_98_3_n237 ), .ZN(_add_98_3_n251 ) );
NOR2_X2 _add_98_3_U119  ( .A1(_add_98_3_n251 ), .A2(_add_98_3_n35 ), .ZN(_add_98_3_n248 ) );
NOR2_X2 _add_98_3_U118  ( .A1(_add_98_3_n314 ), .A2(_add_98_3_n15 ), .ZN(_add_98_3_n320 ) );
NOR3_X2 _add_98_3_U117  ( .A1(_add_98_3_n135 ), .A2(_add_98_3_n130 ), .A3(_add_98_3_n131 ), .ZN(_add_98_3_n128 ) );
NOR2_X2 _add_98_3_U116  ( .A1(_add_98_3_n128 ), .A2(_add_98_3_n129 ), .ZN(_add_98_3_n124 ) );
NOR2_X2 _add_98_3_U115  ( .A1(_add_98_3_n124 ), .A2(_add_98_3_n125 ), .ZN(_add_98_3_n121 ) );
NOR2_X2 _add_98_3_U114  ( .A1(_add_98_3_n43 ), .A2(_add_98_3_n52 ), .ZN(_add_98_3_n380 ) );
NOR2_X2 _add_98_3_U113  ( .A1(_add_98_3_n147 ), .A2(_add_98_3_n127 ), .ZN(_add_98_3_n193 ) );
NAND3_X2 _add_98_3_U112  ( .A1(_add_98_3_n217 ), .A2(_add_98_3_n218 ), .A3(_add_98_3_n373 ), .ZN(_add_98_3_n212 ) );
AND3_X2 _add_98_3_U111  ( .A1(_add_98_3_n171 ), .A2(_add_98_3_n159 ), .A3(_add_98_3_n172 ), .ZN(_add_98_3_n30 ) );
NAND3_X2 _add_98_3_U110  ( .A1(_add_98_3_n150 ), .A2(_add_98_3_n151 ), .A3(_add_98_3_n30 ), .ZN(_add_98_3_n122 ) );
NOR3_X2 _add_98_3_U109  ( .A1(_add_98_3_n194 ), .A2(_add_98_3_n147 ), .A3(_add_98_3_n195 ), .ZN(_add_98_3_n192 ) );
NOR2_X2 _add_98_3_U108  ( .A1(_add_98_3_n314 ), .A2(_add_98_3_n15 ), .ZN(_add_98_3_n330 ) );
NOR2_X2 _add_98_3_U107  ( .A1(_add_98_3_n46 ), .A2(_add_98_3_n43 ), .ZN(_add_98_3_n365 ) );
AND3_X2 _add_98_3_U106  ( .A1(_add_98_3_n373 ), .A2(_add_98_3_n217 ), .A3(_add_98_3_n372 ), .ZN(_add_98_3_n29 ) );
NAND3_X2 _add_98_3_U105  ( .A1(_add_98_3_n161 ), .A2(_add_98_3_n10 ), .A3(_add_98_3_n162 ), .ZN(_add_98_3_n160 ) );
NAND3_X2 _add_98_3_U104  ( .A1(_add_98_3_n159 ), .A2(_add_98_3_n150 ), .A3(_add_98_3_n160 ), .ZN(_add_98_3_n157 ) );
NOR2_X2 _add_98_3_U103  ( .A1(_add_98_3_n34 ), .A2(_add_98_3_n379 ), .ZN(_add_98_3_n378 ) );
NAND3_X2 _add_98_3_U102  ( .A1(_add_98_3_n3 ), .A2(_add_98_3_n7 ), .A3(_add_98_3_n378 ), .ZN(_add_98_3_n49 ) );
NOR2_X2 _add_98_3_U101  ( .A1(_add_98_3_n20 ), .A2(_add_98_3_n105 ), .ZN(_add_98_3_n94 ) );
OR3_X4 _add_98_3_U100  ( .A1(_add_98_3_n307 ), .A2(_add_98_3_n308 ), .A3(_add_98_3_n38 ), .ZN(_add_98_3_n28 ) );
OR2_X2 _add_98_3_U99  ( .A1(_add_98_3_n28 ), .A2(_add_98_3_n303 ), .ZN(_add_98_3_n301 ) );
NOR2_X2 _add_98_3_U98  ( .A1(_add_98_3_n210 ), .A2(_add_98_3_n211 ), .ZN(_add_98_3_n209 ) );
NAND3_X2 _add_98_3_U97  ( .A1(_add_98_3_n212 ), .A2(_add_98_3_n213 ), .A3(_add_98_3_n214 ), .ZN(_add_98_3_n208 ) );
NAND3_X2 _add_98_3_U96  ( .A1(_add_98_3_n208 ), .A2(_add_98_3_n209 ), .A3(_add_98_3_n207 ), .ZN(_add_98_3_n206 ) );
NAND3_X2 _add_98_3_U95  ( .A1(_add_98_3_n236 ), .A2(_add_98_3_n204 ), .A3(_add_98_3_n17 ), .ZN(_add_98_3_n232 ) );
NAND3_X2 _add_98_3_U94  ( .A1(_add_98_3_n224 ), .A2(_add_98_3_n310 ), .A3(_add_98_3_n311 ), .ZN(_add_98_3_n133 ) );
NOR2_X2 _add_98_3_U93  ( .A1(_add_98_3_n215 ), .A2(_add_98_3_n216 ), .ZN(_add_98_3_n288 ) );
NAND3_X2 _add_98_3_U92  ( .A1(_add_98_3_n162 ), .A2(_add_98_3_n10 ), .A3(_add_98_3_n161 ), .ZN(_add_98_3_n170 ) );
NOR2_X2 _add_98_3_U91  ( .A1(_add_98_3_n313 ), .A2(_add_98_3_n314 ), .ZN(_add_98_3_n312 ) );
NAND3_X2 _add_98_3_U90  ( .A1(_add_98_3_n6 ), .A2(_add_98_3_n11 ), .A3(_add_98_3_n312 ), .ZN(_add_98_3_n215 ) );
NOR3_X2 _add_98_3_U89  ( .A1(_add_98_3_n259 ), .A2(_add_98_3_n211 ), .A3(_add_98_3_n210 ), .ZN(_add_98_3_n256 ) );
NOR2_X2 _add_98_3_U88  ( .A1(_add_98_3_n256 ), .A2(_add_98_3_n129 ), .ZN(_add_98_3_n254 ) );
NOR2_X2 _add_98_3_U87  ( .A1(_add_98_3_n254 ), .A2(_add_98_3_n255 ), .ZN(_add_98_3_n237 ) );
NOR3_X2 _add_98_3_U86  ( .A1(_add_98_3_n219 ), .A2(_add_98_3_n77 ), .A3(_add_98_3_n1 ), .ZN(_add_98_3_n297 ) );
NOR2_X2 _add_98_3_U85  ( .A1(_add_98_3_n345 ), .A2(_add_98_3_n355 ), .ZN(_add_98_3_n354 ) );
NAND3_X2 _add_98_3_U84  ( .A1(_add_98_3_n352 ), .A2(_add_98_3_n353 ), .A3(_add_98_3_n354 ), .ZN(_add_98_3_n216 ) );
NOR3_X2 _add_98_3_U83  ( .A1(_add_98_3_n191 ), .A2(_add_98_3_n192 ), .A3(_add_98_3_n193 ), .ZN(_add_98_3_n190 ) );
NOR2_X2 _add_98_3_U82  ( .A1(_add_98_3_n269 ), .A2(_add_98_3_n258 ), .ZN(_add_98_3_n264 ) );
NOR2_X2 _add_98_3_U81  ( .A1(_add_98_3_n264 ), .A2(_add_98_3_n197 ), .ZN(_add_98_3_n263 ) );
NOR2_X2 _add_98_3_U80  ( .A1(_add_98_3_n118 ), .A2(_add_98_3_n119 ), .ZN(_add_98_3_n115 ) );
NOR3_X2 _add_98_3_U79  ( .A1(_add_98_3_n121 ), .A2(_add_98_3_n122 ), .A3(_add_98_3_n123 ), .ZN(_add_98_3_n111 ) );
NOR2_X2 _add_98_3_U78  ( .A1(_add_98_3_n111 ), .A2(_add_98_3_n112 ), .ZN(_add_98_3_n106 ) );
NOR2_X2 _add_98_3_U77  ( .A1(_add_98_3_n29 ), .A2(_add_98_3_n49 ), .ZN(_add_98_3_n53 ) );
NOR2_X2 _add_98_3_U76  ( .A1(_add_98_3_n53 ), .A2(_add_98_3_n9 ), .ZN(_add_98_3_n50 ) );
NOR2_X2 _add_98_3_U75  ( .A1(_add_98_3_n129 ), .A2(_add_98_3_n147 ), .ZN(_add_98_3_n205 ) );
NOR2_X2 _add_98_3_U74  ( .A1(_add_98_3_n29 ), .A2(_add_98_3_n49 ), .ZN(_add_98_3_n356 ) );
NOR2_X2 _add_98_3_U73  ( .A1(_add_98_3_n356 ), .A2(_add_98_3_n9 ), .ZN(_add_98_3_n351 ) );
NOR2_X2 _add_98_3_U72  ( .A1(_add_98_3_n351 ), .A2(_add_98_3_n216 ), .ZN(_add_98_3_n338 ) );
NOR2_X2 _add_98_3_U71  ( .A1(_add_98_3_n338 ), .A2(_add_98_3_n323 ), .ZN(_add_98_3_n335 ) );
NOR2_X2 _add_98_3_U70  ( .A1(_add_98_3_n92 ), .A2(_add_98_3_n93 ), .ZN(_add_98_3_n89 ) );
NOR2_X2 _add_98_3_U69  ( .A1(_add_98_3_n215 ), .A2(_add_98_3_n216 ), .ZN(_add_98_3_n213 ) );
NOR2_X2 _add_98_3_U68  ( .A1(_add_98_3_n320 ), .A2(_add_98_3_n321 ), .ZN(_add_98_3_n319 ) );
NOR3_X2 _add_98_3_U67  ( .A1(_add_98_3_n318 ), .A2(_add_98_3_n319 ), .A3(_add_98_3_n21 ), .ZN(_add_98_3_n317 ) );
NOR2_X2 _add_98_3_U66  ( .A1(_add_98_3_n308 ), .A2(_add_98_3_n317 ), .ZN(_add_98_3_n316 ) );
NOR2_X2 _add_98_3_U65  ( .A1(_add_98_3_n29 ), .A2(_add_98_3_n49 ), .ZN(_add_98_3_n322 ) );
NAND3_X2 _add_98_3_U64  ( .A1(_add_98_3_n88 ), .A2(_add_98_3_n14 ), .A3(_add_98_3_n87 ), .ZN(_add_98_3_n144 ) );
NOR3_X2 _add_98_3_U63  ( .A1(_add_98_3_n19 ), .A2(_add_98_3_n12 ), .A3(_add_98_3_n148 ), .ZN(_add_98_3_n143 ) );
NOR2_X2 _add_98_3_U62  ( .A1(_add_98_3_n95 ), .A2(_add_98_3_n96 ), .ZN(_add_98_3_n84 ) );
NOR2_X2 _add_98_3_U61  ( .A1(_add_98_3_n89 ), .A2(_add_98_3_n90 ), .ZN(_add_98_3_n85 ) );
NOR4_X2 _add_98_3_U60  ( .A1(_add_98_3_n322 ), .A2(_add_98_3_n323 ), .A3(_add_98_3_n9 ), .A4(_add_98_3_n321 ), .ZN(_add_98_3_n318 ) );
NOR2_X2 _add_98_3_U59  ( .A1(_add_98_3_n262 ), .A2(_add_98_3_n77 ), .ZN(_add_98_3_n299 ) );
NOR2_X2 _add_98_3_U58  ( .A1(_add_98_3_n49 ), .A2(_add_98_3_n297 ), .ZN(_add_98_3_n296 ) );
NOR2_X2 _add_98_3_U57  ( .A1(_add_98_3_n215 ), .A2(_add_98_3_n216 ), .ZN(_add_98_3_n294 ) );
NAND3_X2 _add_98_3_U56  ( .A1(_add_98_3_n294 ), .A2(_add_98_3_n295 ), .A3(_add_98_3_n296 ), .ZN(_add_98_3_n134 ) );
NAND3_X2 _add_98_3_U55  ( .A1(_add_98_3_n87 ), .A2(_add_98_3_n88 ), .A3(_add_98_3_n13 ), .ZN(_add_98_3_n86 ) );
NOR2_X2 _add_98_3_U54  ( .A1(_add_98_3_n211 ), .A2(_add_98_3_n210 ), .ZN(_add_98_3_n286 ) );
NAND3_X2 _add_98_3_U53  ( .A1(_add_98_3_n286 ), .A2(_add_98_3_n134 ), .A3(_add_98_3_n260 ), .ZN(_add_98_3_n88 ) );
NAND3_X1 _add_98_3_U52  ( .A1(cv_q[84]), .A2(rnd_q[84]), .A3(_add_98_3_n243 ), .ZN(_add_98_3_n203 ) );
OR2_X4 _add_98_3_U51  ( .A1(rnd_q[64]), .A2(cv_q[64]), .ZN(_add_98_3_n374 ));
OR2_X1 _add_98_3_U50  ( .A1(cv_q[81]), .A2(rnd_q[81]), .ZN(_add_98_3_n33 ));
NOR2_X1 _add_98_3_U49  ( .A1(cv_q[81]), .A2(rnd_q[81]), .ZN(_add_98_3_n278 ));
OR2_X4 _add_98_3_U48  ( .A1(rnd_q[82]), .A2(cv_q[82]), .ZN(_add_98_3_n268 ));
NAND2_X1 _add_98_3_U47  ( .A1(cv_q[80]), .A2(rnd_q[80]), .ZN(_add_98_3_n279 ) );
NOR2_X1 _add_98_3_U46  ( .A1(cv_q[65]), .A2(rnd_q[65]), .ZN(_add_98_3_n137 ));
NOR2_X1 _add_98_3_U45  ( .A1(cv_q[81]), .A2(rnd_q[81]), .ZN(_add_98_3_n275 ));
NOR2_X1 _add_98_3_U44  ( .A1(cv_q[84]), .A2(rnd_q[84]), .ZN(_add_98_3_n252 ));
OR2_X4 _add_98_3_U43  ( .A1(rnd_q[86]), .A2(cv_q[86]), .ZN(_add_98_3_n199 ));
NOR2_X1 _add_98_3_U42  ( .A1(cv_q[84]), .A2(rnd_q[84]), .ZN(_add_98_3_n247 ));
NOR2_X1 _add_98_3_U41  ( .A1(cv_q[85]), .A2(rnd_q[85]), .ZN(_add_98_3_n246 ));
NOR2_X1 _add_98_3_U40  ( .A1(cv_q[85]), .A2(rnd_q[85]), .ZN(_add_98_3_n244 ));
OR2_X4 _add_98_3_U39  ( .A1(rnd_q[83]), .A2(cv_q[83]), .ZN(_add_98_3_n196 ));
NOR2_X1 _add_98_3_U38  ( .A1(cv_q[80]), .A2(rnd_q[80]), .ZN(_add_98_3_n276 ));
OR2_X4 _add_98_3_U37  ( .A1(rnd_q[79]), .A2(cv_q[79]), .ZN(_add_98_3_n302 ));
OR2_X4 _add_98_3_U36  ( .A1(rnd_q[75]), .A2(cv_q[75]), .ZN(_add_98_3_n310 ));
NOR2_X1 _add_98_3_U35  ( .A1(cv_q[76]), .A2(rnd_q[76]), .ZN(_add_98_3_n314 ));
NOR2_X1 _add_98_3_U34  ( .A1(rnd_q[68]), .A2(cv_q[68]), .ZN(_add_98_3_n34 ));
NOR2_X1 _add_98_3_U33  ( .A1(cv_q[73]), .A2(rnd_q[73]), .ZN(_add_98_3_n43 ));
NOR2_X1 _add_98_3_U32  ( .A1(cv_q[72]), .A2(rnd_q[72]), .ZN(_add_98_3_n46 ));
NOR2_X1 _add_98_3_U31  ( .A1(cv_q[78]), .A2(rnd_q[78]), .ZN(_add_98_3_n305 ));
NOR2_X1 _add_98_3_U30  ( .A1(cv_q[74]), .A2(rnd_q[74]), .ZN(_add_98_3_n345 ));
NOR2_X1 _add_98_3_U29  ( .A1(cv_q[77]), .A2(rnd_q[77]), .ZN(_add_98_3_n306 ));
AND2_X4 _add_98_3_U28  ( .A1(_add_98_3_n374 ), .A2(_add_98_3_n222 ), .ZN(N93) );
AND2_X4 _add_98_3_U27  ( .A1(_add_98_3_n199 ), .A2(_add_98_3_n204 ), .ZN(_add_98_3_n26 ) );
AND2_X4 _add_98_3_U26  ( .A1(_add_98_3_n151 ), .A2(_add_98_3_n101 ), .ZN(_add_98_3_n25 ) );
AND2_X4 _add_98_3_U25  ( .A1(_add_98_3_n159 ), .A2(_add_98_3_n162 ), .ZN(_add_98_3_n24 ) );
AND2_X4 _add_98_3_U24  ( .A1(_add_98_3_n127 ), .A2(_add_98_3_n196 ), .ZN(_add_98_3_n23 ) );
OR2_X4 _add_98_3_U23  ( .A1(_add_98_3_n306 ), .A2(_add_98_3_n324 ), .ZN(_add_98_3_n22 ) );
OR2_X4 _add_98_3_U22  ( .A1(_add_98_3_n305 ), .A2(_add_98_3_n306 ), .ZN(_add_98_3_n21 ) );
AND2_X4 _add_98_3_U21  ( .A1(_add_98_3_n109 ), .A2(_add_98_3_n110 ), .ZN(_add_98_3_n20 ) );
AND2_X4 _add_98_3_U20  ( .A1(_add_98_3_n153 ), .A2(_add_98_3_n151 ), .ZN(_add_98_3_n19 ) );
AND3_X4 _add_98_3_U19  ( .A1(_add_98_3_n30 ), .A2(_add_98_3_n150 ), .A3(_add_98_3_n163 ), .ZN(_add_98_3_n18 ) );
OR2_X4 _add_98_3_U18  ( .A1(_add_98_3_n237 ), .A2(_add_98_3_n231 ), .ZN(_add_98_3_n17 ) );
OR2_X4 _add_98_3_U17  ( .A1(_add_98_3_n345 ), .A2(_add_98_3_n346 ), .ZN(_add_98_3_n16 ) );
AND2_X4 _add_98_3_U16  ( .A1(_add_98_3_n216 ), .A2(_add_98_3_n334 ), .ZN(_add_98_3_n15 ) );
AND2_X4 _add_98_3_U15  ( .A1(_add_98_3_n103 ), .A2(_add_98_3_n104 ), .ZN(_add_98_3_n14 ) );
AND3_X4 _add_98_3_U14  ( .A1(_add_98_3_n103 ), .A2(_add_98_3_n94 ), .A3(_add_98_3_n104 ), .ZN(_add_98_3_n13 ) );
AND2_X4 _add_98_3_U13  ( .A1(_add_98_3_n149 ), .A2(_add_98_3_n104 ), .ZN(_add_98_3_n12 ) );
OR2_X4 _add_98_3_U12  ( .A1(cv_q[78]), .A2(rnd_q[78]), .ZN(_add_98_3_n11 ));
OR2_X4 _add_98_3_U11  ( .A1(_add_98_3_n178 ), .A2(_add_98_3_n179 ), .ZN(_add_98_3_n10 ) );
AND2_X4 _add_98_3_U10  ( .A1(_add_98_3_n366 ), .A2(_add_98_3_n3 ), .ZN(_add_98_3_n9 ) );
OR2_X4 _add_98_3_U9  ( .A1(cv_q[67]), .A2(rnd_q[67]), .ZN(_add_98_3_n8 ) );
OR2_X4 _add_98_3_U8  ( .A1(cv_q[70]), .A2(rnd_q[70]), .ZN(_add_98_3_n7 ) );
OR2_X4 _add_98_3_U7  ( .A1(cv_q[77]), .A2(rnd_q[77]), .ZN(_add_98_3_n6 ) );
OR3_X4 _add_98_3_U6  ( .A1(_add_98_3_n322 ), .A2(_add_98_3_n9 ), .A3(_add_98_3_n323 ), .ZN(_add_98_3_n5 ) );
OR2_X4 _add_98_3_U5  ( .A1(cv_q[66]), .A2(rnd_q[66]), .ZN(_add_98_3_n4 ) );
OR2_X4 _add_98_3_U4  ( .A1(cv_q[71]), .A2(rnd_q[71]), .ZN(_add_98_3_n3 ) );
OR2_X4 _add_98_3_U3  ( .A1(cv_q[65]), .A2(rnd_q[65]), .ZN(_add_98_3_n2 ) );
AND3_X4 _add_98_3_U2  ( .A1(_add_98_3_n4 ), .A2(_add_98_3_n8 ), .A3(_add_98_3_n2 ), .ZN(_add_98_3_n1 ) );
INV_X4 _add_98_5_U424  ( .A(rnd_q[0]), .ZN(_add_98_5_n391 ) );
INV_X4 _add_98_5_U423  ( .A(cv_q[0]), .ZN(_add_98_5_n392 ) );
NAND2_X2 _add_98_5_U422  ( .A1(_add_98_5_n391 ), .A2(_add_98_5_n392 ), .ZN(_add_98_5_n381 ) );
NAND2_X2 _add_98_5_U421  ( .A1(rnd_q[0]), .A2(cv_q[0]), .ZN(_add_98_5_n221 ));
INV_X4 _add_98_5_U420  ( .A(_add_98_5_n352 ), .ZN(_add_98_5_n390 ) );
NAND2_X2 _add_98_5_U419  ( .A1(rnd_q[10]), .A2(cv_q[10]), .ZN(_add_98_5_n351 ) );
NAND2_X2 _add_98_5_U418  ( .A1(_add_98_5_n390 ), .A2(_add_98_5_n351 ), .ZN(_add_98_5_n368 ) );
NAND2_X2 _add_98_5_U417  ( .A1(rnd_q[8]), .A2(cv_q[8]), .ZN(_add_98_5_n53 ));
INV_X4 _add_98_5_U416  ( .A(rnd_q[4]), .ZN(_add_98_5_n387 ) );
INV_X4 _add_98_5_U415  ( .A(cv_q[4]), .ZN(_add_98_5_n388 ) );
INV_X4 _add_98_5_U414  ( .A(_add_98_5_n50 ), .ZN(_add_98_5_n378 ) );
NAND2_X2 _add_98_5_U413  ( .A1(rnd_q[1]), .A2(cv_q[1]), .ZN(_add_98_5_n384 ));
NAND2_X2 _add_98_5_U412  ( .A1(_add_98_5_n384 ), .A2(_add_98_5_n221 ), .ZN(_add_98_5_n383 ) );
NAND2_X2 _add_98_5_U411  ( .A1(_add_98_5_n1 ), .A2(_add_98_5_n383 ), .ZN(_add_98_5_n380 ) );
NAND2_X2 _add_98_5_U410  ( .A1(cv_q[2]), .A2(rnd_q[2]), .ZN(_add_98_5_n382 ));
NAND2_X2 _add_98_5_U409  ( .A1(rnd_q[3]), .A2(cv_q[3]), .ZN(_add_98_5_n215 ));
INV_X4 _add_98_5_U408  ( .A(_add_98_5_n33 ), .ZN(_add_98_5_n379 ) );
NAND2_X2 _add_98_5_U407  ( .A1(rnd_q[7]), .A2(cv_q[7]), .ZN(_add_98_5_n57 ));
NAND2_X2 _add_98_5_U406  ( .A1(rnd_q[6]), .A2(cv_q[6]), .ZN(_add_98_5_n377 ));
NAND2_X2 _add_98_5_U405  ( .A1(rnd_q[4]), .A2(cv_q[4]), .ZN(_add_98_5_n67 ));
NAND2_X2 _add_98_5_U404  ( .A1(rnd_q[5]), .A2(cv_q[5]), .ZN(_add_98_5_n64 ));
NAND2_X2 _add_98_5_U403  ( .A1(_add_98_5_n67 ), .A2(_add_98_5_n64 ), .ZN(_add_98_5_n376 ) );
NAND2_X2 _add_98_5_U402  ( .A1(_add_98_5_n375 ), .A2(_add_98_5_n376 ), .ZN(_add_98_5_n374 ) );
NAND2_X2 _add_98_5_U401  ( .A1(_add_98_5_n38 ), .A2(_add_98_5_n374 ), .ZN(_add_98_5_n373 ) );
NAND2_X2 _add_98_5_U400  ( .A1(_add_98_5_n19 ), .A2(_add_98_5_n372 ), .ZN(_add_98_5_n371 ) );
XNOR2_X2 _add_98_5_U399  ( .A(_add_98_5_n368 ), .B(_add_98_5_n367 ), .ZN(N167) );
NAND2_X2 _add_98_5_U398  ( .A1(_add_98_5_n367 ), .A2(_add_98_5_n390 ), .ZN(_add_98_5_n366 ) );
NAND2_X2 _add_98_5_U397  ( .A1(_add_98_5_n366 ), .A2(_add_98_5_n351 ), .ZN(_add_98_5_n364 ) );
NAND2_X2 _add_98_5_U396  ( .A1(rnd_q[11]), .A2(cv_q[11]), .ZN(_add_98_5_n350 ) );
NAND2_X2 _add_98_5_U395  ( .A1(_add_98_5_n350 ), .A2(_add_98_5_n315 ), .ZN(_add_98_5_n365 ) );
XNOR2_X2 _add_98_5_U394  ( .A(_add_98_5_n364 ), .B(_add_98_5_n365 ), .ZN(N168) );
INV_X4 _add_98_5_U393  ( .A(_add_98_5_n44 ), .ZN(_add_98_5_n359 ) );
INV_X4 _add_98_5_U392  ( .A(_add_98_5_n47 ), .ZN(_add_98_5_n360 ) );
INV_X4 _add_98_5_U391  ( .A(_add_98_5_n315 ), .ZN(_add_98_5_n362 ) );
NAND2_X2 _add_98_5_U390  ( .A1(_add_98_5_n354 ), .A2(_add_98_5_n355 ), .ZN(_add_98_5_n346 ) );
NAND2_X2 _add_98_5_U389  ( .A1(cv_q[9]), .A2(rnd_q[9]), .ZN(_add_98_5_n353 ));
INV_X4 _add_98_5_U388  ( .A(_add_98_5_n351 ), .ZN(_add_98_5_n348 ) );
INV_X4 _add_98_5_U387  ( .A(_add_98_5_n350 ), .ZN(_add_98_5_n349 ) );
NAND2_X2 _add_98_5_U386  ( .A1(_add_98_5_n316 ), .A2(_add_98_5_n315 ), .ZN(_add_98_5_n341 ) );
INV_X4 _add_98_5_U385  ( .A(_add_98_5_n341 ), .ZN(_add_98_5_n328 ) );
NAND2_X2 _add_98_5_U384  ( .A1(rnd_q[12]), .A2(cv_q[12]), .ZN(_add_98_5_n329 ) );
INV_X4 _add_98_5_U383  ( .A(_add_98_5_n329 ), .ZN(_add_98_5_n344 ) );
XNOR2_X2 _add_98_5_U382  ( .A(_add_98_5_n342 ), .B(_add_98_5_n343 ), .ZN(N169) );
NAND2_X2 _add_98_5_U381  ( .A1(_add_98_5_n337 ), .A2(_add_98_5_n6 ), .ZN(_add_98_5_n340 ) );
NAND2_X2 _add_98_5_U380  ( .A1(_add_98_5_n340 ), .A2(_add_98_5_n329 ), .ZN(_add_98_5_n338 ) );
NAND2_X2 _add_98_5_U379  ( .A1(rnd_q[13]), .A2(cv_q[13]), .ZN(_add_98_5_n330 ) );
NAND2_X2 _add_98_5_U378  ( .A1(_add_98_5_n330 ), .A2(_add_98_5_n4 ), .ZN(_add_98_5_n339 ) );
XNOR2_X2 _add_98_5_U377  ( .A(_add_98_5_n338 ), .B(_add_98_5_n339 ), .ZN(N170) );
NAND2_X2 _add_98_5_U376  ( .A1(rnd_q[14]), .A2(cv_q[14]), .ZN(_add_98_5_n331 ) );
NAND2_X2 _add_98_5_U375  ( .A1(_add_98_5_n9 ), .A2(_add_98_5_n331 ), .ZN(_add_98_5_n335 ) );
XNOR2_X2 _add_98_5_U374  ( .A(_add_98_5_n334 ), .B(_add_98_5_n335 ), .ZN(N171) );
INV_X4 _add_98_5_U373  ( .A(rnd_q[15]), .ZN(_add_98_5_n332 ) );
INV_X4 _add_98_5_U372  ( .A(cv_q[15]), .ZN(_add_98_5_n333 ) );
NAND2_X2 _add_98_5_U371  ( .A1(_add_98_5_n332 ), .A2(_add_98_5_n333 ), .ZN(_add_98_5_n306 ) );
INV_X4 _add_98_5_U370  ( .A(_add_98_5_n306 ), .ZN(_add_98_5_n318 ) );
INV_X4 _add_98_5_U369  ( .A(_add_98_5_n331 ), .ZN(_add_98_5_n312 ) );
NAND2_X2 _add_98_5_U368  ( .A1(_add_98_5_n329 ), .A2(_add_98_5_n330 ), .ZN(_add_98_5_n326 ) );
XNOR2_X2 _add_98_5_U367  ( .A(_add_98_5_n320 ), .B(_add_98_5_n321 ), .ZN(N172) );
NAND2_X2 _add_98_5_U366  ( .A1(rnd_q[16]), .A2(cv_q[16]), .ZN(_add_98_5_n287 ) );
NAND2_X2 _add_98_5_U365  ( .A1(_add_98_5_n287 ), .A2(_add_98_5_n289 ), .ZN(_add_98_5_n290 ) );
INV_X4 _add_98_5_U364  ( .A(_add_98_5_n213 ), .ZN(_add_98_5_n314 ) );
INV_X4 _add_98_5_U363  ( .A(_add_98_5_n132 ), .ZN(_add_98_5_n210 ) );
NAND2_X2 _add_98_5_U362  ( .A1(cv_q[13]), .A2(rnd_q[13]), .ZN(_add_98_5_n313 ) );
NAND2_X2 _add_98_5_U361  ( .A1(rnd_q[12]), .A2(cv_q[12]), .ZN(_add_98_5_n308 ) );
NAND2_X2 _add_98_5_U360  ( .A1(_add_98_5_n305 ), .A2(_add_98_5_n306 ), .ZN(_add_98_5_n131 ) );
INV_X4 _add_98_5_U359  ( .A(_add_98_5_n131 ), .ZN(_add_98_5_n209 ) );
NAND2_X2 _add_98_5_U358  ( .A1(rnd_q[1]), .A2(cv_q[1]), .ZN(_add_98_5_n137 ));
INV_X4 _add_98_5_U357  ( .A(_add_98_5_n137 ), .ZN(_add_98_5_n262 ) );
INV_X4 _add_98_5_U356  ( .A(_add_98_5_n215 ), .ZN(_add_98_5_n78 ) );
NAND2_X2 _add_98_5_U355  ( .A1(_add_98_5_n303 ), .A2(_add_98_5_n304 ), .ZN(_add_98_5_n300 ) );
NAND2_X2 _add_98_5_U354  ( .A1(rnd_q[5]), .A2(cv_q[5]), .ZN(_add_98_5_n296 ));
NAND2_X2 _add_98_5_U353  ( .A1(_add_98_5_n67 ), .A2(_add_98_5_n296 ), .ZN(_add_98_5_n295 ) );
NAND2_X2 _add_98_5_U352  ( .A1(_add_98_5_n225 ), .A2(_add_98_5_n295 ), .ZN(_add_98_5_n294 ) );
NAND2_X2 _add_98_5_U351  ( .A1(_add_98_5_n38 ), .A2(_add_98_5_n294 ), .ZN(_add_98_5_n292 ) );
NAND3_X2 _add_98_5_U350  ( .A1(_add_98_5_n292 ), .A2(_add_98_5_n3 ), .A3(_add_98_5_n293 ), .ZN(_add_98_5_n260 ) );
INV_X4 _add_98_5_U349  ( .A(_add_98_5_n260 ), .ZN(_add_98_5_n134 ) );
XNOR2_X2 _add_98_5_U348  ( .A(_add_98_5_n290 ), .B(_add_98_5_n89 ), .ZN(N173) );
INV_X4 _add_98_5_U347  ( .A(_add_98_5_n281 ), .ZN(_add_98_5_n289 ) );
NAND2_X2 _add_98_5_U346  ( .A1(_add_98_5_n89 ), .A2(_add_98_5_n289 ), .ZN(_add_98_5_n288 ) );
NAND2_X2 _add_98_5_U345  ( .A1(_add_98_5_n287 ), .A2(_add_98_5_n288 ), .ZN(_add_98_5_n285 ) );
NAND2_X2 _add_98_5_U344  ( .A1(rnd_q[17]), .A2(cv_q[17]), .ZN(_add_98_5_n282 ) );
NAND2_X2 _add_98_5_U343  ( .A1(_add_98_5_n39 ), .A2(_add_98_5_n282 ), .ZN(_add_98_5_n286 ) );
XNOR2_X2 _add_98_5_U342  ( .A(_add_98_5_n285 ), .B(_add_98_5_n286 ), .ZN(N174) );
NAND2_X2 _add_98_5_U341  ( .A1(cv_q[16]), .A2(rnd_q[16]), .ZN(_add_98_5_n284 ) );
NAND2_X2 _add_98_5_U340  ( .A1(_add_98_5_n31 ), .A2(_add_98_5_n282 ), .ZN(_add_98_5_n270 ) );
INV_X4 _add_98_5_U339  ( .A(_add_98_5_n270 ), .ZN(_add_98_5_n278 ) );
NAND2_X2 _add_98_5_U338  ( .A1(_add_98_5_n273 ), .A2(_add_98_5_n89 ), .ZN(_add_98_5_n279 ) );
NAND2_X2 _add_98_5_U337  ( .A1(_add_98_5_n278 ), .A2(_add_98_5_n279 ), .ZN(_add_98_5_n274 ) );
NAND2_X2 _add_98_5_U336  ( .A1(rnd_q[18]), .A2(cv_q[18]), .ZN(_add_98_5_n269 ) );
INV_X4 _add_98_5_U335  ( .A(rnd_q[18]), .ZN(_add_98_5_n276 ) );
INV_X4 _add_98_5_U334  ( .A(cv_q[18]), .ZN(_add_98_5_n277 ) );
NAND2_X2 _add_98_5_U333  ( .A1(_add_98_5_n276 ), .A2(_add_98_5_n277 ), .ZN(_add_98_5_n271 ) );
NAND2_X2 _add_98_5_U332  ( .A1(_add_98_5_n269 ), .A2(_add_98_5_n271 ), .ZN(_add_98_5_n275 ) );
XNOR2_X2 _add_98_5_U331  ( .A(_add_98_5_n274 ), .B(_add_98_5_n275 ), .ZN(N175) );
INV_X4 _add_98_5_U330  ( .A(_add_98_5_n89 ), .ZN(_add_98_5_n272 ) );
NAND2_X2 _add_98_5_U329  ( .A1(_add_98_5_n273 ), .A2(_add_98_5_n271 ), .ZN(_add_98_5_n258 ) );
NAND2_X2 _add_98_5_U328  ( .A1(_add_98_5_n270 ), .A2(_add_98_5_n271 ), .ZN(_add_98_5_n268 ) );
NAND2_X2 _add_98_5_U327  ( .A1(_add_98_5_n268 ), .A2(_add_98_5_n269 ), .ZN(_add_98_5_n196 ) );
NAND2_X2 _add_98_5_U326  ( .A1(rnd_q[19]), .A2(cv_q[19]), .ZN(_add_98_5_n126 ) );
INV_X4 _add_98_5_U325  ( .A(rnd_q[19]), .ZN(_add_98_5_n265 ) );
INV_X4 _add_98_5_U324  ( .A(cv_q[19]), .ZN(_add_98_5_n266 ) );
NAND2_X2 _add_98_5_U323  ( .A1(_add_98_5_n265 ), .A2(_add_98_5_n266 ), .ZN(_add_98_5_n195 ) );
XNOR2_X2 _add_98_5_U322  ( .A(_add_98_5_n264 ), .B(_add_98_5_n25 ), .ZN(N176) );
INV_X4 _add_98_5_U321  ( .A(_add_98_5_n221 ), .ZN(_add_98_5_n263 ) );
XNOR2_X2 _add_98_5_U320  ( .A(_add_98_5_n221 ), .B(_add_98_5_n261 ), .ZN(N158) );
INV_X4 _add_98_5_U319  ( .A(_add_98_5_n258 ), .ZN(_add_98_5_n257 ) );
NAND2_X2 _add_98_5_U318  ( .A1(_add_98_5_n257 ), .A2(_add_98_5_n195 ), .ZN(_add_98_5_n128 ) );
NAND2_X2 _add_98_5_U317  ( .A1(_add_98_5_n196 ), .A2(_add_98_5_n195 ), .ZN(_add_98_5_n125 ) );
NAND2_X2 _add_98_5_U316  ( .A1(_add_98_5_n125 ), .A2(_add_98_5_n126 ), .ZN(_add_98_5_n255 ) );
XNOR2_X2 _add_98_5_U315  ( .A(_add_98_5_n235 ), .B(_add_98_5_n253 ), .ZN(N177) );
NAND2_X2 _add_98_5_U314  ( .A1(rnd_q[21]), .A2(cv_q[21]), .ZN(_add_98_5_n201 ) );
INV_X4 _add_98_5_U313  ( .A(_add_98_5_n201 ), .ZN(_add_98_5_n250 ) );
XNOR2_X2 _add_98_5_U312  ( .A(_add_98_5_n248 ), .B(_add_98_5_n249 ), .ZN(N178) );
INV_X4 _add_98_5_U311  ( .A(_add_98_5_n236 ), .ZN(_add_98_5_n245 ) );
INV_X4 _add_98_5_U310  ( .A(_add_98_5_n244 ), .ZN(_add_98_5_n243 ) );
NAND2_X2 _add_98_5_U309  ( .A1(_add_98_5_n202 ), .A2(_add_98_5_n201 ), .ZN(_add_98_5_n242 ) );
INV_X4 _add_98_5_U308  ( .A(rnd_q[22]), .ZN(_add_98_5_n239 ) );
INV_X4 _add_98_5_U307  ( .A(cv_q[22]), .ZN(_add_98_5_n240 ) );
NAND2_X2 _add_98_5_U306  ( .A1(_add_98_5_n239 ), .A2(_add_98_5_n240 ), .ZN(_add_98_5_n198 ) );
NAND2_X2 _add_98_5_U305  ( .A1(rnd_q[22]), .A2(cv_q[22]), .ZN(_add_98_5_n203 ) );
XNOR2_X2 _add_98_5_U304  ( .A(_add_98_5_n238 ), .B(_add_98_5_n28 ), .ZN(N179) );
NAND2_X2 _add_98_5_U303  ( .A1(_add_98_5_n202 ), .A2(_add_98_5_n201 ), .ZN(_add_98_5_n237 ) );
NAND2_X2 _add_98_5_U302  ( .A1(_add_98_5_n237 ), .A2(_add_98_5_n198 ), .ZN(_add_98_5_n234 ) );
NAND2_X2 _add_98_5_U301  ( .A1(_add_98_5_n236 ), .A2(_add_98_5_n198 ), .ZN(_add_98_5_n229 ) );
INV_X4 _add_98_5_U300  ( .A(rnd_q[23]), .ZN(_add_98_5_n232 ) );
INV_X4 _add_98_5_U299  ( .A(cv_q[23]), .ZN(_add_98_5_n233 ) );
NAND2_X2 _add_98_5_U298  ( .A1(_add_98_5_n232 ), .A2(_add_98_5_n233 ), .ZN(_add_98_5_n199 ) );
NAND2_X2 _add_98_5_U297  ( .A1(rnd_q[23]), .A2(cv_q[23]), .ZN(_add_98_5_n151 ) );
NAND2_X2 _add_98_5_U296  ( .A1(_add_98_5_n199 ), .A2(_add_98_5_n151 ), .ZN(_add_98_5_n231 ) );
XNOR2_X2 _add_98_5_U295  ( .A(_add_98_5_n230 ), .B(_add_98_5_n231 ), .ZN(N180) );
INV_X4 _add_98_5_U294  ( .A(_add_98_5_n229 ), .ZN(_add_98_5_n228 ) );
NAND2_X2 _add_98_5_U293  ( .A1(_add_98_5_n228 ), .A2(_add_98_5_n199 ), .ZN(_add_98_5_n146 ) );
NAND2_X2 _add_98_5_U292  ( .A1(rnd_q[5]), .A2(cv_q[5]), .ZN(_add_98_5_n227 ));
NAND2_X2 _add_98_5_U291  ( .A1(_add_98_5_n67 ), .A2(_add_98_5_n227 ), .ZN(_add_98_5_n226 ) );
NAND2_X2 _add_98_5_U290  ( .A1(_add_98_5_n225 ), .A2(_add_98_5_n226 ), .ZN(_add_98_5_n224 ) );
NAND2_X2 _add_98_5_U289  ( .A1(_add_98_5_n38 ), .A2(_add_98_5_n224 ), .ZN(_add_98_5_n222 ) );
INV_X4 _add_98_5_U288  ( .A(_add_98_5_n214 ), .ZN(_add_98_5_n223 ) );
NAND4_X2 _add_98_5_U287  ( .A1(_add_98_5_n222 ), .A2(_add_98_5_n3 ), .A3(_add_98_5_n314 ), .A4(_add_98_5_n223 ), .ZN(_add_98_5_n206 ) );
NAND2_X2 _add_98_5_U286  ( .A1(rnd_q[1]), .A2(cv_q[1]), .ZN(_add_98_5_n220 ));
NAND2_X2 _add_98_5_U285  ( .A1(_add_98_5_n220 ), .A2(_add_98_5_n221 ), .ZN(_add_98_5_n219 ) );
NAND2_X2 _add_98_5_U284  ( .A1(_add_98_5_n1 ), .A2(_add_98_5_n219 ), .ZN(_add_98_5_n216 ) );
INV_X4 _add_98_5_U283  ( .A(_add_98_5_n218 ), .ZN(_add_98_5_n217 ) );
NAND2_X2 _add_98_5_U282  ( .A1(_add_98_5_n204 ), .A2(_add_98_5_n205 ), .ZN(_add_98_5_n188 ) );
INV_X4 _add_98_5_U281  ( .A(_add_98_5_n145 ), .ZN(_add_98_5_n197 ) );
NAND2_X2 _add_98_5_U280  ( .A1(_add_98_5_n197 ), .A2(_add_98_5_n151 ), .ZN(_add_98_5_n190 ) );
INV_X4 _add_98_5_U279  ( .A(_add_98_5_n196 ), .ZN(_add_98_5_n193 ) );
INV_X4 _add_98_5_U278  ( .A(_add_98_5_n195 ), .ZN(_add_98_5_n194 ) );
NAND2_X2 _add_98_5_U277  ( .A1(_add_98_5_n188 ), .A2(_add_98_5_n189 ), .ZN(_add_98_5_n162 ) );
NAND2_X2 _add_98_5_U276  ( .A1(rnd_q[24]), .A2(cv_q[24]), .ZN(_add_98_5_n186 ) );
NAND2_X2 _add_98_5_U275  ( .A1(_add_98_5_n186 ), .A2(_add_98_5_n171 ), .ZN(_add_98_5_n187 ) );
XNOR2_X2 _add_98_5_U274  ( .A(_add_98_5_n162 ), .B(_add_98_5_n187 ), .ZN(N181) );
INV_X4 _add_98_5_U273  ( .A(_add_98_5_n180 ), .ZN(_add_98_5_n171 ) );
NAND2_X2 _add_98_5_U272  ( .A1(_add_98_5_n171 ), .A2(_add_98_5_n162 ), .ZN(_add_98_5_n185 ) );
NAND2_X2 _add_98_5_U271  ( .A1(_add_98_5_n185 ), .A2(_add_98_5_n186 ), .ZN(_add_98_5_n181 ) );
NAND2_X2 _add_98_5_U270  ( .A1(rnd_q[25]), .A2(cv_q[25]), .ZN(_add_98_5_n160 ) );
INV_X4 _add_98_5_U269  ( .A(rnd_q[25]), .ZN(_add_98_5_n183 ) );
INV_X4 _add_98_5_U268  ( .A(cv_q[25]), .ZN(_add_98_5_n184 ) );
NAND2_X2 _add_98_5_U267  ( .A1(_add_98_5_n183 ), .A2(_add_98_5_n184 ), .ZN(_add_98_5_n170 ) );
NAND2_X2 _add_98_5_U266  ( .A1(_add_98_5_n160 ), .A2(_add_98_5_n170 ), .ZN(_add_98_5_n182 ) );
XNOR2_X2 _add_98_5_U265  ( .A(_add_98_5_n181 ), .B(_add_98_5_n182 ), .ZN(N182) );
INV_X4 _add_98_5_U264  ( .A(_add_98_5_n162 ), .ZN(_add_98_5_n179 ) );
INV_X4 _add_98_5_U263  ( .A(_add_98_5_n170 ), .ZN(_add_98_5_n177 ) );
NAND2_X2 _add_98_5_U262  ( .A1(cv_q[24]), .A2(rnd_q[24]), .ZN(_add_98_5_n178 ) );
NAND2_X2 _add_98_5_U261  ( .A1(_add_98_5_n8 ), .A2(_add_98_5_n160 ), .ZN(_add_98_5_n176 ) );
INV_X4 _add_98_5_U260  ( .A(rnd_q[26]), .ZN(_add_98_5_n173 ) );
INV_X4 _add_98_5_U259  ( .A(cv_q[26]), .ZN(_add_98_5_n174 ) );
NAND2_X2 _add_98_5_U258  ( .A1(_add_98_5_n173 ), .A2(_add_98_5_n174 ), .ZN(_add_98_5_n158 ) );
NAND2_X2 _add_98_5_U257  ( .A1(rnd_q[26]), .A2(cv_q[26]), .ZN(_add_98_5_n161 ) );
XNOR2_X2 _add_98_5_U256  ( .A(_add_98_5_n172 ), .B(_add_98_5_n27 ), .ZN(N183) );
NAND2_X2 _add_98_5_U255  ( .A1(_add_98_5_n34 ), .A2(_add_98_5_n162 ), .ZN(_add_98_5_n167 ) );
NAND2_X2 _add_98_5_U254  ( .A1(_add_98_5_n169 ), .A2(_add_98_5_n158 ), .ZN(_add_98_5_n168 ) );
NAND2_X2 _add_98_5_U253  ( .A1(_add_98_5_n167 ), .A2(_add_98_5_n168 ), .ZN(_add_98_5_n163 ) );
INV_X4 _add_98_5_U252  ( .A(rnd_q[27]), .ZN(_add_98_5_n165 ) );
INV_X4 _add_98_5_U251  ( .A(cv_q[27]), .ZN(_add_98_5_n166 ) );
NAND2_X2 _add_98_5_U250  ( .A1(_add_98_5_n165 ), .A2(_add_98_5_n166 ), .ZN(_add_98_5_n149 ) );
NAND2_X2 _add_98_5_U249  ( .A1(rnd_q[27]), .A2(cv_q[27]), .ZN(_add_98_5_n157 ) );
NAND2_X2 _add_98_5_U248  ( .A1(_add_98_5_n149 ), .A2(_add_98_5_n157 ), .ZN(_add_98_5_n164 ) );
XNOR2_X2 _add_98_5_U247  ( .A(_add_98_5_n163 ), .B(_add_98_5_n164 ), .ZN(N184) );
NAND2_X2 _add_98_5_U246  ( .A1(_add_98_5_n156 ), .A2(_add_98_5_n157 ), .ZN(_add_98_5_n152 ) );
INV_X4 _add_98_5_U245  ( .A(rnd_q[28]), .ZN(_add_98_5_n154 ) );
INV_X4 _add_98_5_U244  ( .A(cv_q[28]), .ZN(_add_98_5_n155 ) );
NAND2_X2 _add_98_5_U243  ( .A1(_add_98_5_n154 ), .A2(_add_98_5_n155 ), .ZN(_add_98_5_n150 ) );
NAND2_X2 _add_98_5_U242  ( .A1(rnd_q[28]), .A2(cv_q[28]), .ZN(_add_98_5_n102 ) );
XNOR2_X2 _add_98_5_U241  ( .A(_add_98_5_n153 ), .B(_add_98_5_n29 ), .ZN(N185) );
INV_X4 _add_98_5_U240  ( .A(_add_98_5_n151 ), .ZN(_add_98_5_n148 ) );
INV_X4 _add_98_5_U239  ( .A(_add_98_5_n121 ), .ZN(_add_98_5_n105 ) );
INV_X4 _add_98_5_U238  ( .A(_add_98_5_n102 ), .ZN(_add_98_5_n147 ) );
INV_X4 _add_98_5_U237  ( .A(_add_98_5_n146 ), .ZN(_add_98_5_n104 ) );
INV_X4 _add_98_5_U236  ( .A(_add_98_5_n128 ), .ZN(_add_98_5_n88 ) );
NAND2_X2 _add_98_5_U235  ( .A1(_add_98_5_n125 ), .A2(_add_98_5_n126 ), .ZN(_add_98_5_n103 ) );
NAND2_X2 _add_98_5_U234  ( .A1(_add_98_5_n103 ), .A2(_add_98_5_n13 ), .ZN(_add_98_5_n144 ) );
NAND2_X2 _add_98_5_U233  ( .A1(_add_98_5_n145 ), .A2(_add_98_5_n105 ), .ZN(_add_98_5_n94 ) );
NAND4_X2 _add_98_5_U232  ( .A1(_add_98_5_n142 ), .A2(_add_98_5_n143 ), .A3(_add_98_5_n144 ), .A4(_add_98_5_n94 ), .ZN(_add_98_5_n138 ) );
NAND2_X2 _add_98_5_U231  ( .A1(rnd_q[29]), .A2(cv_q[29]), .ZN(_add_98_5_n92 ) );
INV_X4 _add_98_5_U230  ( .A(rnd_q[29]), .ZN(_add_98_5_n140 ) );
INV_X4 _add_98_5_U229  ( .A(cv_q[29]), .ZN(_add_98_5_n141 ) );
NAND2_X2 _add_98_5_U228  ( .A1(_add_98_5_n140 ), .A2(_add_98_5_n141 ), .ZN(_add_98_5_n118 ) );
NAND2_X2 _add_98_5_U227  ( .A1(_add_98_5_n92 ), .A2(_add_98_5_n118 ), .ZN(_add_98_5_n139 ) );
XNOR2_X2 _add_98_5_U226  ( .A(_add_98_5_n138 ), .B(_add_98_5_n139 ), .ZN(N186) );
XNOR2_X2 _add_98_5_U225  ( .A(_add_98_5_n81 ), .B(_add_98_5_n135 ), .ZN(N159) );
INV_X4 _add_98_5_U224  ( .A(_add_98_5_n133 ), .ZN(_add_98_5_n129 ) );
NAND2_X2 _add_98_5_U223  ( .A1(_add_98_5_n131 ), .A2(_add_98_5_n132 ), .ZN(_add_98_5_n130 ) );
NAND2_X2 _add_98_5_U222  ( .A1(_add_98_5_n125 ), .A2(_add_98_5_n126 ), .ZN(_add_98_5_n124 ) );
NAND2_X2 _add_98_5_U221  ( .A1(_add_98_5_n104 ), .A2(_add_98_5_n118 ), .ZN(_add_98_5_n122 ) );
NAND2_X2 _add_98_5_U220  ( .A1(_add_98_5_n21 ), .A2(_add_98_5_n118 ), .ZN(_add_98_5_n114 ) );
INV_X4 _add_98_5_U219  ( .A(_add_98_5_n94 ), .ZN(_add_98_5_n119 ) );
NAND2_X2 _add_98_5_U218  ( .A1(_add_98_5_n119 ), .A2(_add_98_5_n118 ), .ZN(_add_98_5_n115 ) );
INV_X4 _add_98_5_U217  ( .A(_add_98_5_n118 ), .ZN(_add_98_5_n106 ) );
NAND2_X2 _add_98_5_U216  ( .A1(_add_98_5_n11 ), .A2(_add_98_5_n118 ), .ZN(_add_98_5_n117 ) );
NAND4_X2 _add_98_5_U215  ( .A1(_add_98_5_n114 ), .A2(_add_98_5_n115 ), .A3(_add_98_5_n116 ), .A4(_add_98_5_n117 ), .ZN(_add_98_5_n113 ) );
INV_X4 _add_98_5_U214  ( .A(rnd_q[30]), .ZN(_add_98_5_n110 ) );
INV_X4 _add_98_5_U213  ( .A(cv_q[30]), .ZN(_add_98_5_n111 ) );
NAND2_X2 _add_98_5_U212  ( .A1(rnd_q[30]), .A2(cv_q[30]), .ZN(_add_98_5_n101 ) );
INV_X4 _add_98_5_U211  ( .A(_add_98_5_n101 ), .ZN(_add_98_5_n109 ) );
XNOR2_X2 _add_98_5_U210  ( .A(_add_98_5_n107 ), .B(_add_98_5_n108 ), .ZN(N187) );
NAND2_X2 _add_98_5_U209  ( .A1(_add_98_5_n12 ), .A2(_add_98_5_n103 ), .ZN(_add_98_5_n84 ) );
NAND2_X2 _add_98_5_U208  ( .A1(_add_98_5_n95 ), .A2(_add_98_5_n147 ), .ZN(_add_98_5_n100 ) );
NAND2_X2 _add_98_5_U207  ( .A1(_add_98_5_n100 ), .A2(_add_98_5_n101 ), .ZN(_add_98_5_n96 ) );
NAND2_X2 _add_98_5_U206  ( .A1(_add_98_5_n21 ), .A2(_add_98_5_n95 ), .ZN(_add_98_5_n98 ) );
NAND2_X2 _add_98_5_U205  ( .A1(_add_98_5_n11 ), .A2(_add_98_5_n95 ), .ZN(_add_98_5_n99 ) );
NAND2_X2 _add_98_5_U204  ( .A1(_add_98_5_n98 ), .A2(_add_98_5_n99 ), .ZN(_add_98_5_n97 ) );
INV_X4 _add_98_5_U203  ( .A(_add_98_5_n95 ), .ZN(_add_98_5_n93 ) );
NAND4_X2 _add_98_5_U202  ( .A1(_add_98_5_n84 ), .A2(_add_98_5_n85 ), .A3(_add_98_5_n86 ), .A4(_add_98_5_n87 ), .ZN(_add_98_5_n82 ) );
XNOR2_X2 _add_98_5_U201  ( .A(rnd_q[31]), .B(cv_q[31]), .ZN(_add_98_5_n83 ));
XNOR2_X2 _add_98_5_U200  ( .A(_add_98_5_n82 ), .B(_add_98_5_n83 ), .ZN(N188));
XNOR2_X2 _add_98_5_U199  ( .A(_add_98_5_n75 ), .B(_add_98_5_n76 ), .ZN(N160));
INV_X4 _add_98_5_U198  ( .A(_add_98_5_n67 ), .ZN(_add_98_5_n73 ) );
XNOR2_X2 _add_98_5_U197  ( .A(_add_98_5_n33 ), .B(_add_98_5_n74 ), .ZN(N161));
INV_X4 _add_98_5_U196  ( .A(_add_98_5_n64 ), .ZN(_add_98_5_n71 ) );
XNOR2_X2 _add_98_5_U195  ( .A(_add_98_5_n69 ), .B(_add_98_5_n70 ), .ZN(N162));
NAND2_X2 _add_98_5_U194  ( .A1(rnd_q[6]), .A2(cv_q[6]), .ZN(_add_98_5_n59 ));
NAND2_X2 _add_98_5_U193  ( .A1(_add_98_5_n59 ), .A2(_add_98_5_n5 ), .ZN(_add_98_5_n62 ) );
NAND2_X2 _add_98_5_U192  ( .A1(_add_98_5_n33 ), .A2(_add_98_5_n67 ), .ZN(_add_98_5_n66 ) );
NAND2_X2 _add_98_5_U191  ( .A1(_add_98_5_n65 ), .A2(_add_98_5_n66 ), .ZN(_add_98_5_n63 ) );
NAND2_X2 _add_98_5_U190  ( .A1(_add_98_5_n63 ), .A2(_add_98_5_n64 ), .ZN(_add_98_5_n60 ) );
XNOR2_X2 _add_98_5_U189  ( .A(_add_98_5_n62 ), .B(_add_98_5_n60 ), .ZN(N163));
NAND2_X2 _add_98_5_U188  ( .A1(_add_98_5_n60 ), .A2(_add_98_5_n5 ), .ZN(_add_98_5_n58 ) );
NAND2_X2 _add_98_5_U187  ( .A1(_add_98_5_n58 ), .A2(_add_98_5_n59 ), .ZN(_add_98_5_n55 ) );
NAND2_X2 _add_98_5_U186  ( .A1(_add_98_5_n57 ), .A2(_add_98_5_n3 ), .ZN(_add_98_5_n56 ) );
XNOR2_X2 _add_98_5_U185  ( .A(_add_98_5_n55 ), .B(_add_98_5_n56 ), .ZN(N164));
INV_X4 _add_98_5_U184  ( .A(_add_98_5_n53 ), .ZN(_add_98_5_n46 ) );
XNOR2_X2 _add_98_5_U183  ( .A(_add_98_5_n51 ), .B(_add_98_5_n52 ), .ZN(N165));
XNOR2_X2 _add_98_5_U182  ( .A(_add_98_5_n42 ), .B(_add_98_5_n43 ), .ZN(N166));
NAND2_X2 _add_98_5_U181  ( .A1(_add_98_5_n260 ), .A2(_add_98_5_n133 ), .ZN(_add_98_5_n259 ) );
NOR2_X2 _add_98_5_U180  ( .A1(_add_98_5_n20 ), .A2(_add_98_5_n109 ), .ZN(_add_98_5_n108 ) );
NOR2_X2 _add_98_5_U179  ( .A1(_add_98_5_n14 ), .A2(_add_98_5_n73 ), .ZN(_add_98_5_n74 ) );
NOR2_X2 _add_98_5_U178  ( .A1(_add_98_5_n262 ), .A2(_add_98_5_n136 ), .ZN(_add_98_5_n261 ) );
AND2_X2 _add_98_5_U177  ( .A1(cv_q[8]), .A2(rnd_q[8]), .ZN(_add_98_5_n354 ));
NOR2_X2 _add_98_5_U176  ( .A1(cv_q[9]), .A2(rnd_q[9]), .ZN(_add_98_5_n356 ));
NOR2_X2 _add_98_5_U175  ( .A1(cv_q[10]), .A2(rnd_q[10]), .ZN(_add_98_5_n357 ) );
NOR2_X2 _add_98_5_U174  ( .A1(_add_98_5_n356 ), .A2(_add_98_5_n357 ), .ZN(_add_98_5_n355 ) );
NOR2_X2 _add_98_5_U173  ( .A1(_add_98_5_n47 ), .A2(_add_98_5_n46 ), .ZN(_add_98_5_n52 ) );
NOR2_X2 _add_98_5_U172  ( .A1(_add_98_5_n77 ), .A2(_add_98_5_n78 ), .ZN(_add_98_5_n76 ) );
AND2_X2 _add_98_5_U171  ( .A1(rnd_q[2]), .A2(cv_q[2]), .ZN(_add_98_5_n41 ));
AND2_X2 _add_98_5_U170  ( .A1(rnd_q[9]), .A2(cv_q[9]), .ZN(_add_98_5_n40 ));
OR2_X2 _add_98_5_U169  ( .A1(cv_q[17]), .A2(rnd_q[17]), .ZN(_add_98_5_n39 ));
NOR2_X2 _add_98_5_U168  ( .A1(cv_q[17]), .A2(rnd_q[17]), .ZN(_add_98_5_n280 ) );
NOR2_X2 _add_98_5_U167  ( .A1(_add_98_5_n280 ), .A2(_add_98_5_n281 ), .ZN(_add_98_5_n273 ) );
NOR2_X2 _add_98_5_U166  ( .A1(cv_q[5]), .A2(rnd_q[5]), .ZN(_add_98_5_n297 ));
NOR2_X2 _add_98_5_U165  ( .A1(cv_q[6]), .A2(rnd_q[6]), .ZN(_add_98_5_n298 ));
NOR2_X2 _add_98_5_U164  ( .A1(_add_98_5_n297 ), .A2(_add_98_5_n298 ), .ZN(_add_98_5_n225 ) );
NOR2_X2 _add_98_5_U163  ( .A1(_add_98_5_n309 ), .A2(_add_98_5_n313 ), .ZN(_add_98_5_n311 ) );
NOR2_X2 _add_98_5_U162  ( .A1(_add_98_5_n22 ), .A2(_add_98_5_n252 ), .ZN(_add_98_5_n253 ) );
NOR2_X2 _add_98_5_U161  ( .A1(_add_98_5_n41 ), .A2(_add_98_5_n80 ), .ZN(_add_98_5_n135 ) );
NOR2_X2 _add_98_5_U160  ( .A1(_add_98_5_n344 ), .A2(_add_98_5_n319 ), .ZN(_add_98_5_n343 ) );
NOR2_X2 _add_98_5_U159  ( .A1(_add_98_5_n244 ), .A2(_add_98_5_n250 ), .ZN(_add_98_5_n249 ) );
NOR2_X2 _add_98_5_U158  ( .A1(_add_98_5_n40 ), .A2(_add_98_5_n44 ), .ZN(_add_98_5_n43 ) );
NOR2_X2 _add_98_5_U157  ( .A1(_add_98_5_n71 ), .A2(_add_98_5_n68 ), .ZN(_add_98_5_n70 ) );
NOR2_X2 _add_98_5_U156  ( .A1(_add_98_5_n318 ), .A2(_add_98_5_n15 ), .ZN(_add_98_5_n320 ) );
AND2_X2 _add_98_5_U155  ( .A1(_add_98_5_n57 ), .A2(_add_98_5_n377 ), .ZN(_add_98_5_n38 ) );
NOR2_X2 _add_98_5_U154  ( .A1(cv_q[5]), .A2(rnd_q[5]), .ZN(_add_98_5_n386 ));
NOR2_X2 _add_98_5_U153  ( .A1(cv_q[21]), .A2(rnd_q[21]), .ZN(_add_98_5_n244 ) );
NOR2_X2 _add_98_5_U152  ( .A1(cv_q[17]), .A2(rnd_q[17]), .ZN(_add_98_5_n283 ) );
NOR2_X2 _add_98_5_U151  ( .A1(cv_q[3]), .A2(rnd_q[3]), .ZN(_add_98_5_n77 ));
NOR2_X2 _add_98_5_U150  ( .A1(cv_q[2]), .A2(rnd_q[2]), .ZN(_add_98_5_n80 ));
NOR2_X2 _add_98_5_U149  ( .A1(cv_q[1]), .A2(rnd_q[1]), .ZN(_add_98_5_n136 ));
NOR2_X2 _add_98_5_U148  ( .A1(cv_q[20]), .A2(rnd_q[20]), .ZN(_add_98_5_n252 ) );
NAND3_X2 _add_98_5_U147  ( .A1(cv_q[20]), .A2(rnd_q[20]), .A3(_add_98_5_n243 ), .ZN(_add_98_5_n202 ) );
NOR2_X2 _add_98_5_U146  ( .A1(cv_q[16]), .A2(rnd_q[16]), .ZN(_add_98_5_n281 ) );
NOR2_X2 _add_98_5_U145  ( .A1(cv_q[6]), .A2(rnd_q[6]), .ZN(_add_98_5_n61 ));
NOR2_X2 _add_98_5_U144  ( .A1(cv_q[24]), .A2(rnd_q[24]), .ZN(_add_98_5_n180 ) );
NOR2_X2 _add_98_5_U143  ( .A1(cv_q[5]), .A2(rnd_q[5]), .ZN(_add_98_5_n68 ));
NOR2_X2 _add_98_5_U142  ( .A1(_add_98_5_n77 ), .A2(_add_98_5_n382 ), .ZN(_add_98_5_n218 ) );
NOR2_X2 _add_98_5_U141  ( .A1(cv_q[14]), .A2(rnd_q[14]), .ZN(_add_98_5_n309 ) );
NOR3_X2 _add_98_5_U140  ( .A1(_add_98_5_n308 ), .A2(_add_98_5_n309 ), .A3(_add_98_5_n310 ), .ZN(_add_98_5_n307 ) );
NOR2_X2 _add_98_5_U139  ( .A1(cv_q[20]), .A2(rnd_q[20]), .ZN(_add_98_5_n247 ) );
NOR2_X2 _add_98_5_U138  ( .A1(cv_q[21]), .A2(rnd_q[21]), .ZN(_add_98_5_n246 ) );
NOR2_X2 _add_98_5_U137  ( .A1(_add_98_5_n246 ), .A2(_add_98_5_n247 ), .ZN(_add_98_5_n236 ) );
NOR2_X2 _add_98_5_U136  ( .A1(cv_q[10]), .A2(rnd_q[10]), .ZN(_add_98_5_n352 ) );
NOR2_X2 _add_98_5_U135  ( .A1(cv_q[8]), .A2(rnd_q[8]), .ZN(_add_98_5_n47 ));
NOR2_X2 _add_98_5_U134  ( .A1(cv_q[9]), .A2(rnd_q[9]), .ZN(_add_98_5_n44 ));
NOR2_X2 _add_98_5_U133  ( .A1(cv_q[12]), .A2(rnd_q[12]), .ZN(_add_98_5_n319 ) );
NOR2_X2 _add_98_5_U132  ( .A1(cv_q[13]), .A2(rnd_q[13]), .ZN(_add_98_5_n310 ) );
NAND3_X2 _add_98_5_U131  ( .A1(_add_98_5_n201 ), .A2(_add_98_5_n202 ), .A3(_add_98_5_n203 ), .ZN(_add_98_5_n200 ) );
AND2_X4 _add_98_5_U130  ( .A1(_add_98_5_n198 ), .A2(_add_98_5_n199 ), .ZN(_add_98_5_n37 ) );
AND2_X2 _add_98_5_U129  ( .A1(_add_98_5_n200 ), .A2(_add_98_5_n37 ), .ZN(_add_98_5_n145 ) );
NOR2_X2 _add_98_5_U128  ( .A1(_add_98_5_n18 ), .A2(_add_98_5_n152 ), .ZN(_add_98_5_n153 ) );
NOR2_X2 _add_98_5_U127  ( .A1(_add_98_5_n263 ), .A2(_add_98_5_n218 ), .ZN(_add_98_5_n303 ) );
NOR2_X2 _add_98_5_U126  ( .A1(_add_98_5_n96 ), .A2(_add_98_5_n97 ), .ZN(_add_98_5_n85 ) );
OR2_X4 _add_98_5_U125  ( .A1(_add_98_5_n106 ), .A2(_add_98_5_n102 ), .ZN(_add_98_5_n36 ) );
AND2_X2 _add_98_5_U124  ( .A1(_add_98_5_n92 ), .A2(_add_98_5_n36 ), .ZN(_add_98_5_n116 ) );
NAND3_X2 _add_98_5_U123  ( .A1(_add_98_5_n378 ), .A2(_add_98_5_n372 ), .A3(_add_98_5_n379 ), .ZN(_add_98_5_n370 ) );
NOR2_X2 _add_98_5_U122  ( .A1(_add_98_5_n40 ), .A2(_add_98_5_n389 ), .ZN(_add_98_5_n369 ) );
NAND3_X2 _add_98_5_U121  ( .A1(_add_98_5_n369 ), .A2(_add_98_5_n370 ), .A3(_add_98_5_n371 ), .ZN(_add_98_5_n367 ) );
NAND3_X2 _add_98_5_U120  ( .A1(_add_98_5_n337 ), .A2(_add_98_5_n4 ), .A3(_add_98_5_n6 ), .ZN(_add_98_5_n336 ) );
NAND3_X2 _add_98_5_U119  ( .A1(_add_98_5_n26 ), .A2(_add_98_5_n330 ), .A3(_add_98_5_n336 ), .ZN(_add_98_5_n334 ) );
NOR2_X2 _add_98_5_U118  ( .A1(_add_98_5_n80 ), .A2(_add_98_5_n81 ), .ZN(_add_98_5_n79 ) );
NOR2_X2 _add_98_5_U117  ( .A1(_add_98_5_n79 ), .A2(_add_98_5_n41 ), .ZN(_add_98_5_n75 ) );
NOR2_X2 _add_98_5_U116  ( .A1(_add_98_5_n235 ), .A2(_add_98_5_n245 ), .ZN(_add_98_5_n241 ) );
NOR2_X2 _add_98_5_U115  ( .A1(_add_98_5_n241 ), .A2(_add_98_5_n242 ), .ZN(_add_98_5_n238 ) );
NOR2_X2 _add_98_5_U114  ( .A1(_add_98_5_n33 ), .A2(_add_98_5_n50 ), .ZN(_add_98_5_n49 ) );
NOR2_X2 _add_98_5_U113  ( .A1(_add_98_5_n49 ), .A2(_add_98_5_n19 ), .ZN(_add_98_5_n48 ) );
NOR2_X2 _add_98_5_U112  ( .A1(_add_98_5_n47 ), .A2(_add_98_5_n48 ), .ZN(_add_98_5_n45 ) );
NOR2_X2 _add_98_5_U111  ( .A1(_add_98_5_n45 ), .A2(_add_98_5_n46 ), .ZN(_add_98_5_n42 ) );
NOR2_X2 _add_98_5_U110  ( .A1(_add_98_5_n252 ), .A2(_add_98_5_n235 ), .ZN(_add_98_5_n251 ) );
NOR2_X2 _add_98_5_U109  ( .A1(_add_98_5_n251 ), .A2(_add_98_5_n22 ), .ZN(_add_98_5_n248 ) );
NOR2_X2 _add_98_5_U108  ( .A1(_add_98_5_n33 ), .A2(_add_98_5_n14 ), .ZN(_add_98_5_n72 ) );
NOR2_X2 _add_98_5_U107  ( .A1(_add_98_5_n72 ), .A2(_add_98_5_n73 ), .ZN(_add_98_5_n69 ) );
NOR2_X2 _add_98_5_U106  ( .A1(_add_98_5_n61 ), .A2(_add_98_5_n68 ), .ZN(_add_98_5_n375 ) );
NOR2_X2 _add_98_5_U105  ( .A1(_add_98_5_n348 ), .A2(_add_98_5_n349 ), .ZN(_add_98_5_n347 ) );
NAND3_X2 _add_98_5_U104  ( .A1(_add_98_5_n346 ), .A2(_add_98_5_n16 ), .A3(_add_98_5_n347 ), .ZN(_add_98_5_n316 ) );
NOR2_X2 _add_98_5_U103  ( .A1(_add_98_5_n14 ), .A2(_add_98_5_n68 ), .ZN(_add_98_5_n65 ) );
NAND3_X2 _add_98_5_U102  ( .A1(_add_98_5_n314 ), .A2(_add_98_5_n315 ), .A3(_add_98_5_n316 ), .ZN(_add_98_5_n132 ) );
NOR2_X2 _add_98_5_U101  ( .A1(_add_98_5_n20 ), .A2(_add_98_5_n92 ), .ZN(_add_98_5_n91 ) );
NOR2_X2 _add_98_5_U100  ( .A1(_add_98_5_n319 ), .A2(_add_98_5_n23 ), .ZN(_add_98_5_n325 ) );
NAND3_X2 _add_98_5_U99  ( .A1(_add_98_5_n160 ), .A2(_add_98_5_n8 ), .A3(_add_98_5_n161 ), .ZN(_add_98_5_n159 ) );
NAND3_X2 _add_98_5_U98  ( .A1(_add_98_5_n158 ), .A2(_add_98_5_n149 ), .A3(_add_98_5_n159 ), .ZN(_add_98_5_n156 ) );
NOR2_X2 _add_98_5_U97  ( .A1(_add_98_5_n44 ), .A2(_add_98_5_n53 ), .ZN(_add_98_5_n389 ) );
NAND3_X2 _add_98_5_U96  ( .A1(_add_98_5_n215 ), .A2(_add_98_5_n216 ), .A3(_add_98_5_n217 ), .ZN(_add_98_5_n211 ) );
NOR3_X2 _add_98_5_U95  ( .A1(_add_98_5_n134 ), .A2(_add_98_5_n129 ), .A3(_add_98_5_n130 ), .ZN(_add_98_5_n127 ) );
NOR2_X2 _add_98_5_U94  ( .A1(_add_98_5_n127 ), .A2(_add_98_5_n128 ), .ZN(_add_98_5_n123 ) );
NOR2_X2 _add_98_5_U93  ( .A1(_add_98_5_n123 ), .A2(_add_98_5_n124 ), .ZN(_add_98_5_n120 ) );
NOR3_X2 _add_98_5_U92  ( .A1(_add_98_5_n179 ), .A2(_add_98_5_n177 ), .A3(_add_98_5_n180 ), .ZN(_add_98_5_n175 ) );
NOR2_X2 _add_98_5_U91  ( .A1(_add_98_5_n175 ), .A2(_add_98_5_n176 ), .ZN(_add_98_5_n172 ) );
OR2_X4 _add_98_5_U90  ( .A1(_add_98_5_n136 ), .A2(_add_98_5_n221 ), .ZN(_add_98_5_n35 ) );
AND2_X2 _add_98_5_U89  ( .A1(_add_98_5_n137 ), .A2(_add_98_5_n35 ), .ZN(_add_98_5_n81 ) );
AND3_X2 _add_98_5_U88  ( .A1(_add_98_5_n170 ), .A2(_add_98_5_n158 ), .A3(_add_98_5_n171 ), .ZN(_add_98_5_n34 ) );
NAND3_X2 _add_98_5_U87  ( .A1(_add_98_5_n149 ), .A2(_add_98_5_n150 ), .A3(_add_98_5_n34 ), .ZN(_add_98_5_n121 ) );
NOR2_X2 _add_98_5_U86  ( .A1(_add_98_5_n319 ), .A2(_add_98_5_n23 ), .ZN(_add_98_5_n337 ) );
NOR2_X2 _add_98_5_U85  ( .A1(_add_98_5_n47 ), .A2(_add_98_5_n44 ), .ZN(_add_98_5_n372 ) );
AND3_X2 _add_98_5_U84  ( .A1(_add_98_5_n217 ), .A2(_add_98_5_n215 ), .A3(_add_98_5_n380 ), .ZN(_add_98_5_n33 ) );
NOR2_X2 _add_98_5_U83  ( .A1(_add_98_5_n14 ), .A2(_add_98_5_n386 ), .ZN(_add_98_5_n385 ) );
NAND3_X2 _add_98_5_U82  ( .A1(_add_98_5_n3 ), .A2(_add_98_5_n5 ), .A3(_add_98_5_n385 ), .ZN(_add_98_5_n50 ) );
NOR3_X2 _add_98_5_U81  ( .A1(_add_98_5_n120 ), .A2(_add_98_5_n121 ), .A3(_add_98_5_n122 ), .ZN(_add_98_5_n112 ) );
NOR2_X2 _add_98_5_U80  ( .A1(_add_98_5_n112 ), .A2(_add_98_5_n113 ), .ZN(_add_98_5_n107 ) );
NOR2_X2 _add_98_5_U79  ( .A1(_add_98_5_n20 ), .A2(_add_98_5_n106 ), .ZN(_add_98_5_n95 ) );
NAND3_X2 _add_98_5_U78  ( .A1(_add_98_5_n234 ), .A2(_add_98_5_n203 ), .A3(_add_98_5_n17 ), .ZN(_add_98_5_n230 ) );
NOR2_X2 _add_98_5_U77  ( .A1(_add_98_5_n213 ), .A2(_add_98_5_n214 ), .ZN(_add_98_5_n293 ) );
NAND3_X2 _add_98_5_U76  ( .A1(_add_98_5_n161 ), .A2(_add_98_5_n8 ), .A3(_add_98_5_n160 ), .ZN(_add_98_5_n169 ) );
NOR2_X2 _add_98_5_U75  ( .A1(_add_98_5_n146 ), .A2(_add_98_5_n126 ), .ZN(_add_98_5_n192 ) );
NOR2_X2 _add_98_5_U74  ( .A1(_add_98_5_n209 ), .A2(_add_98_5_n210 ), .ZN(_add_98_5_n208 ) );
NAND3_X2 _add_98_5_U73  ( .A1(_add_98_5_n211 ), .A2(_add_98_5_n212 ), .A3(_add_98_5_n378 ), .ZN(_add_98_5_n207 ) );
NAND3_X2 _add_98_5_U72  ( .A1(_add_98_5_n207 ), .A2(_add_98_5_n208 ), .A3(_add_98_5_n206 ), .ZN(_add_98_5_n205 ) );
NOR3_X2 _add_98_5_U71  ( .A1(_add_98_5_n259 ), .A2(_add_98_5_n210 ), .A3(_add_98_5_n209 ), .ZN(_add_98_5_n256 ) );
NOR2_X2 _add_98_5_U70  ( .A1(_add_98_5_n256 ), .A2(_add_98_5_n128 ), .ZN(_add_98_5_n254 ) );
NOR2_X2 _add_98_5_U69  ( .A1(_add_98_5_n254 ), .A2(_add_98_5_n255 ), .ZN(_add_98_5_n235 ) );
NOR3_X2 _add_98_5_U68  ( .A1(_add_98_5_n218 ), .A2(_add_98_5_n78 ), .A3(_add_98_5_n1 ), .ZN(_add_98_5_n302 ) );
NOR2_X2 _add_98_5_U67  ( .A1(_add_98_5_n318 ), .A2(_add_98_5_n319 ), .ZN(_add_98_5_n317 ) );
NAND3_X2 _add_98_5_U66  ( .A1(_add_98_5_n4 ), .A2(_add_98_5_n9 ), .A3(_add_98_5_n317 ), .ZN(_add_98_5_n213 ) );
NOR3_X2 _add_98_5_U65  ( .A1(_add_98_5_n193 ), .A2(_add_98_5_n146 ), .A3(_add_98_5_n194 ), .ZN(_add_98_5_n191 ) );
OR3_X4 _add_98_5_U64  ( .A1(_add_98_5_n311 ), .A2(_add_98_5_n312 ), .A3(_add_98_5_n15 ), .ZN(_add_98_5_n32 ) );
OR2_X2 _add_98_5_U63  ( .A1(_add_98_5_n32 ), .A2(_add_98_5_n307 ), .ZN(_add_98_5_n305 ) );
NOR2_X2 _add_98_5_U62  ( .A1(_add_98_5_n352 ), .A2(_add_98_5_n362 ), .ZN(_add_98_5_n361 ) );
NAND3_X2 _add_98_5_U61  ( .A1(_add_98_5_n359 ), .A2(_add_98_5_n360 ), .A3(_add_98_5_n361 ), .ZN(_add_98_5_n214 ) );
NOR2_X2 _add_98_5_U60  ( .A1(_add_98_5_n262 ), .A2(_add_98_5_n78 ), .ZN(_add_98_5_n304 ) );
NOR2_X2 _add_98_5_U59  ( .A1(_add_98_5_n325 ), .A2(_add_98_5_n326 ), .ZN(_add_98_5_n324 ) );
NOR3_X2 _add_98_5_U58  ( .A1(_add_98_5_n323 ), .A2(_add_98_5_n324 ), .A3(_add_98_5_n24 ), .ZN(_add_98_5_n322 ) );
NOR2_X2 _add_98_5_U57  ( .A1(_add_98_5_n312 ), .A2(_add_98_5_n322 ), .ZN(_add_98_5_n321 ) );
NOR2_X2 _add_98_5_U56  ( .A1(_add_98_5_n33 ), .A2(_add_98_5_n50 ), .ZN(_add_98_5_n54 ) );
NOR2_X2 _add_98_5_U55  ( .A1(_add_98_5_n54 ), .A2(_add_98_5_n19 ), .ZN(_add_98_5_n51 ) );
NOR2_X2 _add_98_5_U54  ( .A1(_add_98_5_n272 ), .A2(_add_98_5_n258 ), .ZN(_add_98_5_n267 ) );
NOR2_X2 _add_98_5_U53  ( .A1(_add_98_5_n267 ), .A2(_add_98_5_n196 ), .ZN(_add_98_5_n264 ) );
NOR2_X2 _add_98_5_U52  ( .A1(_add_98_5_n33 ), .A2(_add_98_5_n50 ), .ZN(_add_98_5_n363 ) );
NOR2_X2 _add_98_5_U51  ( .A1(_add_98_5_n363 ), .A2(_add_98_5_n19 ), .ZN(_add_98_5_n358 ) );
NOR2_X2 _add_98_5_U50  ( .A1(_add_98_5_n358 ), .A2(_add_98_5_n214 ), .ZN(_add_98_5_n345 ) );
NOR2_X2 _add_98_5_U49  ( .A1(_add_98_5_n345 ), .A2(_add_98_5_n328 ), .ZN(_add_98_5_n342 ) );
NOR2_X2 _add_98_5_U48  ( .A1(_add_98_5_n93 ), .A2(_add_98_5_n94 ), .ZN(_add_98_5_n90 ) );
NOR2_X2 _add_98_5_U47  ( .A1(_add_98_5_n213 ), .A2(_add_98_5_n214 ), .ZN(_add_98_5_n212 ) );
NOR2_X2 _add_98_5_U46  ( .A1(_add_98_5_n33 ), .A2(_add_98_5_n50 ), .ZN(_add_98_5_n327 ) );
NAND3_X2 _add_98_5_U45  ( .A1(_add_98_5_n89 ), .A2(_add_98_5_n13 ), .A3(_add_98_5_n88 ), .ZN(_add_98_5_n143 ) );
NOR3_X2 _add_98_5_U44  ( .A1(_add_98_5_n11 ), .A2(_add_98_5_n21 ), .A3(_add_98_5_n147 ), .ZN(_add_98_5_n142 ) );
NAND3_X2 _add_98_5_U43  ( .A1(_add_98_5_n88 ), .A2(_add_98_5_n89 ), .A3(_add_98_5_n12 ), .ZN(_add_98_5_n87 ) );
NOR2_X2 _add_98_5_U42  ( .A1(_add_98_5_n90 ), .A2(_add_98_5_n91 ), .ZN(_add_98_5_n86 ) );
NOR4_X2 _add_98_5_U41  ( .A1(_add_98_5_n327 ), .A2(_add_98_5_n328 ), .A3(_add_98_5_n19 ), .A4(_add_98_5_n326 ), .ZN(_add_98_5_n323 ) );
NOR2_X2 _add_98_5_U40  ( .A1(_add_98_5_n50 ), .A2(_add_98_5_n302 ), .ZN(_add_98_5_n301 ) );
NOR2_X2 _add_98_5_U39  ( .A1(_add_98_5_n213 ), .A2(_add_98_5_n214 ), .ZN(_add_98_5_n299 ) );
NAND3_X2 _add_98_5_U38  ( .A1(_add_98_5_n299 ), .A2(_add_98_5_n300 ), .A3(_add_98_5_n301 ), .ZN(_add_98_5_n133 ) );
NOR2_X2 _add_98_5_U37  ( .A1(_add_98_5_n128 ), .A2(_add_98_5_n146 ), .ZN(_add_98_5_n204 ) );
NOR3_X2 _add_98_5_U36  ( .A1(_add_98_5_n190 ), .A2(_add_98_5_n191 ), .A3(_add_98_5_n192 ), .ZN(_add_98_5_n189 ) );
NOR2_X2 _add_98_5_U35  ( .A1(_add_98_5_n210 ), .A2(_add_98_5_n209 ), .ZN(_add_98_5_n291 ) );
NAND3_X2 _add_98_5_U34  ( .A1(_add_98_5_n291 ), .A2(_add_98_5_n133 ), .A3(_add_98_5_n260 ), .ZN(_add_98_5_n89 ) );
OR2_X4 _add_98_5_U33  ( .A1(rnd_q[11]), .A2(cv_q[11]), .ZN(_add_98_5_n315 ));
OR2_X4 _add_98_5_U32  ( .A1(_add_98_5_n283 ), .A2(_add_98_5_n284 ), .ZN(_add_98_5_n31 ) );
AND2_X4 _add_98_5_U31  ( .A1(_add_98_5_n381 ), .A2(_add_98_5_n221 ), .ZN(N157) );
AND2_X4 _add_98_5_U30  ( .A1(_add_98_5_n150 ), .A2(_add_98_5_n102 ), .ZN(_add_98_5_n29 ) );
AND2_X4 _add_98_5_U29  ( .A1(_add_98_5_n198 ), .A2(_add_98_5_n203 ), .ZN(_add_98_5_n28 ) );
AND2_X4 _add_98_5_U28  ( .A1(_add_98_5_n158 ), .A2(_add_98_5_n161 ), .ZN(_add_98_5_n27 ) );
OR2_X4 _add_98_5_U27  ( .A1(_add_98_5_n310 ), .A2(_add_98_5_n329 ), .ZN(_add_98_5_n26 ) );
AND2_X4 _add_98_5_U26  ( .A1(_add_98_5_n126 ), .A2(_add_98_5_n195 ), .ZN(_add_98_5_n25 ) );
OR2_X4 _add_98_5_U25  ( .A1(_add_98_5_n309 ), .A2(_add_98_5_n310 ), .ZN(_add_98_5_n24 ) );
AND2_X4 _add_98_5_U24  ( .A1(_add_98_5_n214 ), .A2(_add_98_5_n341 ), .ZN(_add_98_5_n23 ) );
AND2_X4 _add_98_5_U23  ( .A1(rnd_q[20]), .A2(cv_q[20]), .ZN(_add_98_5_n22 ));
AND2_X4 _add_98_5_U22  ( .A1(_add_98_5_n148 ), .A2(_add_98_5_n105 ), .ZN(_add_98_5_n21 ) );
AND2_X4 _add_98_5_U21  ( .A1(_add_98_5_n110 ), .A2(_add_98_5_n111 ), .ZN(_add_98_5_n20 ) );
AND2_X4 _add_98_5_U20  ( .A1(_add_98_5_n373 ), .A2(_add_98_5_n3 ), .ZN(_add_98_5_n19 ) );
AND3_X4 _add_98_5_U19  ( .A1(_add_98_5_n34 ), .A2(_add_98_5_n149 ), .A3(_add_98_5_n162 ), .ZN(_add_98_5_n18 ) );
OR2_X4 _add_98_5_U18  ( .A1(_add_98_5_n235 ), .A2(_add_98_5_n229 ), .ZN(_add_98_5_n17 ) );
OR2_X4 _add_98_5_U17  ( .A1(_add_98_5_n352 ), .A2(_add_98_5_n353 ), .ZN(_add_98_5_n16 ) );
AND2_X4 _add_98_5_U16  ( .A1(rnd_q[15]), .A2(cv_q[15]), .ZN(_add_98_5_n15 ));
AND2_X4 _add_98_5_U15  ( .A1(_add_98_5_n387 ), .A2(_add_98_5_n388 ), .ZN(_add_98_5_n14 ) );
AND2_X4 _add_98_5_U14  ( .A1(_add_98_5_n104 ), .A2(_add_98_5_n105 ), .ZN(_add_98_5_n13 ) );
AND3_X4 _add_98_5_U13  ( .A1(_add_98_5_n104 ), .A2(_add_98_5_n95 ), .A3(_add_98_5_n105 ), .ZN(_add_98_5_n12 ) );
AND2_X4 _add_98_5_U12  ( .A1(_add_98_5_n152 ), .A2(_add_98_5_n150 ), .ZN(_add_98_5_n11 ) );
OR2_X4 _add_98_5_U11  ( .A1(cv_q[3]), .A2(rnd_q[3]), .ZN(_add_98_5_n10 ) );
OR2_X4 _add_98_5_U10  ( .A1(cv_q[14]), .A2(rnd_q[14]), .ZN(_add_98_5_n9 ) );
OR2_X4 _add_98_5_U9  ( .A1(_add_98_5_n177 ), .A2(_add_98_5_n178 ), .ZN(_add_98_5_n8 ) );
OR2_X4 _add_98_5_U8  ( .A1(cv_q[2]), .A2(rnd_q[2]), .ZN(_add_98_5_n7 ) );
OR3_X4 _add_98_5_U7  ( .A1(_add_98_5_n327 ), .A2(_add_98_5_n19 ), .A3(_add_98_5_n328 ), .ZN(_add_98_5_n6 ) );
OR2_X4 _add_98_5_U6  ( .A1(cv_q[6]), .A2(rnd_q[6]), .ZN(_add_98_5_n5 ) );
OR2_X4 _add_98_5_U5  ( .A1(cv_q[13]), .A2(rnd_q[13]), .ZN(_add_98_5_n4 ) );
OR2_X4 _add_98_5_U4  ( .A1(cv_q[7]), .A2(rnd_q[7]), .ZN(_add_98_5_n3 ) );
OR2_X4 _add_98_5_U3  ( .A1(cv_q[1]), .A2(rnd_q[1]), .ZN(_add_98_5_n2 ) );
AND3_X4 _add_98_5_U2  ( .A1(_add_98_5_n7 ), .A2(_add_98_5_n10 ), .A3(_add_98_5_n2 ), .ZN(_add_98_5_n1 ) );
INV_X4 _add_98_U426  ( .A(rnd_q[128]), .ZN(_add_98_n393 ) );
INV_X4 _add_98_U425  ( .A(cv_q[128]), .ZN(_add_98_n394 ) );
NAND2_X2 _add_98_U424  ( .A1(_add_98_n393 ), .A2(_add_98_n394 ), .ZN(_add_98_n383 ) );
NAND2_X2 _add_98_U423  ( .A1(rnd_q[128]), .A2(cv_q[128]), .ZN(_add_98_n220 ));
INV_X4 _add_98_U422  ( .A(_add_98_n351 ), .ZN(_add_98_n392 ) );
NAND2_X2 _add_98_U421  ( .A1(rnd_q[138]), .A2(cv_q[138]), .ZN(_add_98_n350 ));
NAND2_X2 _add_98_U420  ( .A1(_add_98_n392 ), .A2(_add_98_n350 ), .ZN(_add_98_n369 ) );
NAND2_X2 _add_98_U419  ( .A1(rnd_q[136]), .A2(cv_q[136]), .ZN(_add_98_n53 ));
INV_X4 _add_98_U418  ( .A(rnd_q[132]), .ZN(_add_98_n389 ) );
INV_X4 _add_98_U417  ( .A(cv_q[132]), .ZN(_add_98_n390 ) );
INV_X4 _add_98_U416  ( .A(_add_98_n50 ), .ZN(_add_98_n379 ) );
NAND2_X2 _add_98_U415  ( .A1(rnd_q[129]), .A2(cv_q[129]), .ZN(_add_98_n386 ));
NAND2_X2 _add_98_U414  ( .A1(_add_98_n386 ), .A2(_add_98_n220 ), .ZN(_add_98_n385 ) );
NAND2_X2 _add_98_U413  ( .A1(_add_98_n1 ), .A2(_add_98_n385 ), .ZN(_add_98_n381 ) );
NAND2_X2 _add_98_U412  ( .A1(cv_q[130]), .A2(rnd_q[130]), .ZN(_add_98_n384 ));
INV_X4 _add_98_U411  ( .A(_add_98_n217 ), .ZN(_add_98_n382 ) );
NAND2_X2 _add_98_U410  ( .A1(rnd_q[131]), .A2(cv_q[131]), .ZN(_add_98_n215 ));
INV_X4 _add_98_U409  ( .A(_add_98_n35 ), .ZN(_add_98_n380 ) );
NAND2_X2 _add_98_U408  ( .A1(rnd_q[135]), .A2(cv_q[135]), .ZN(_add_98_n57 ));
NAND2_X2 _add_98_U407  ( .A1(rnd_q[134]), .A2(cv_q[134]), .ZN(_add_98_n378 ));
NAND2_X2 _add_98_U406  ( .A1(rnd_q[132]), .A2(cv_q[132]), .ZN(_add_98_n67 ));
NAND2_X2 _add_98_U405  ( .A1(rnd_q[133]), .A2(cv_q[133]), .ZN(_add_98_n64 ));
NAND2_X2 _add_98_U404  ( .A1(_add_98_n67 ), .A2(_add_98_n64 ), .ZN(_add_98_n377 ) );
NAND2_X2 _add_98_U403  ( .A1(_add_98_n376 ), .A2(_add_98_n377 ), .ZN(_add_98_n375 ) );
NAND2_X2 _add_98_U402  ( .A1(_add_98_n22 ), .A2(_add_98_n375 ), .ZN(_add_98_n374 ) );
NAND2_X2 _add_98_U401  ( .A1(_add_98_n19 ), .A2(_add_98_n373 ), .ZN(_add_98_n372 ) );
XNOR2_X2 _add_98_U400  ( .A(_add_98_n369 ), .B(_add_98_n368 ), .ZN(N39) );
NAND2_X2 _add_98_U399  ( .A1(_add_98_n368 ), .A2(_add_98_n392 ), .ZN(_add_98_n367 ) );
NAND2_X2 _add_98_U398  ( .A1(_add_98_n367 ), .A2(_add_98_n350 ), .ZN(_add_98_n363 ) );
NAND2_X2 _add_98_U397  ( .A1(rnd_q[139]), .A2(cv_q[139]), .ZN(_add_98_n349 ));
INV_X4 _add_98_U396  ( .A(rnd_q[139]), .ZN(_add_98_n365 ) );
INV_X4 _add_98_U395  ( .A(cv_q[139]), .ZN(_add_98_n366 ) );
NAND2_X2 _add_98_U394  ( .A1(_add_98_n365 ), .A2(_add_98_n366 ), .ZN(_add_98_n314 ) );
NAND2_X2 _add_98_U393  ( .A1(_add_98_n349 ), .A2(_add_98_n314 ), .ZN(_add_98_n364 ) );
XNOR2_X2 _add_98_U392  ( .A(_add_98_n363 ), .B(_add_98_n364 ), .ZN(N40) );
INV_X4 _add_98_U391  ( .A(_add_98_n44 ), .ZN(_add_98_n358 ) );
INV_X4 _add_98_U390  ( .A(_add_98_n47 ), .ZN(_add_98_n359 ) );
INV_X4 _add_98_U389  ( .A(_add_98_n314 ), .ZN(_add_98_n361 ) );
NAND2_X2 _add_98_U388  ( .A1(_add_98_n353 ), .A2(_add_98_n354 ), .ZN(_add_98_n345 ) );
NAND2_X2 _add_98_U387  ( .A1(cv_q[137]), .A2(rnd_q[137]), .ZN(_add_98_n352 ));
INV_X4 _add_98_U386  ( .A(_add_98_n350 ), .ZN(_add_98_n347 ) );
INV_X4 _add_98_U385  ( .A(_add_98_n349 ), .ZN(_add_98_n348 ) );
NAND2_X2 _add_98_U384  ( .A1(_add_98_n315 ), .A2(_add_98_n314 ), .ZN(_add_98_n340 ) );
INV_X4 _add_98_U383  ( .A(_add_98_n340 ), .ZN(_add_98_n327 ) );
NAND2_X2 _add_98_U382  ( .A1(rnd_q[140]), .A2(cv_q[140]), .ZN(_add_98_n328 ));
INV_X4 _add_98_U381  ( .A(_add_98_n328 ), .ZN(_add_98_n343 ) );
XNOR2_X2 _add_98_U380  ( .A(_add_98_n341 ), .B(_add_98_n342 ), .ZN(N41) );
NAND2_X2 _add_98_U379  ( .A1(_add_98_n336 ), .A2(_add_98_n6 ), .ZN(_add_98_n339 ) );
NAND2_X2 _add_98_U378  ( .A1(_add_98_n339 ), .A2(_add_98_n328 ), .ZN(_add_98_n337 ) );
NAND2_X2 _add_98_U377  ( .A1(rnd_q[141]), .A2(cv_q[141]), .ZN(_add_98_n329 ));
NAND2_X2 _add_98_U376  ( .A1(_add_98_n329 ), .A2(_add_98_n4 ), .ZN(_add_98_n338 ) );
XNOR2_X2 _add_98_U375  ( .A(_add_98_n337 ), .B(_add_98_n338 ), .ZN(N42) );
NAND2_X2 _add_98_U374  ( .A1(rnd_q[142]), .A2(cv_q[142]), .ZN(_add_98_n330 ));
NAND2_X2 _add_98_U373  ( .A1(_add_98_n9 ), .A2(_add_98_n330 ), .ZN(_add_98_n334 ) );
XNOR2_X2 _add_98_U372  ( .A(_add_98_n333 ), .B(_add_98_n334 ), .ZN(N43) );
INV_X4 _add_98_U371  ( .A(rnd_q[143]), .ZN(_add_98_n331 ) );
INV_X4 _add_98_U370  ( .A(cv_q[143]), .ZN(_add_98_n332 ) );
NAND2_X2 _add_98_U369  ( .A1(_add_98_n331 ), .A2(_add_98_n332 ), .ZN(_add_98_n305 ) );
INV_X4 _add_98_U368  ( .A(_add_98_n305 ), .ZN(_add_98_n317 ) );
INV_X4 _add_98_U367  ( .A(_add_98_n330 ), .ZN(_add_98_n311 ) );
NAND2_X2 _add_98_U366  ( .A1(_add_98_n328 ), .A2(_add_98_n329 ), .ZN(_add_98_n325 ) );
XNOR2_X2 _add_98_U365  ( .A(_add_98_n319 ), .B(_add_98_n320 ), .ZN(N44) );
NAND2_X2 _add_98_U364  ( .A1(rnd_q[144]), .A2(cv_q[144]), .ZN(_add_98_n285 ));
NAND2_X2 _add_98_U363  ( .A1(_add_98_n285 ), .A2(_add_98_n287 ), .ZN(_add_98_n288 ) );
INV_X4 _add_98_U362  ( .A(_add_98_n213 ), .ZN(_add_98_n313 ) );
INV_X4 _add_98_U361  ( .A(_add_98_n132 ), .ZN(_add_98_n210 ) );
NAND2_X2 _add_98_U360  ( .A1(cv_q[141]), .A2(rnd_q[141]), .ZN(_add_98_n312 ));
NAND2_X2 _add_98_U359  ( .A1(rnd_q[140]), .A2(cv_q[140]), .ZN(_add_98_n307 ));
NAND2_X2 _add_98_U358  ( .A1(_add_98_n304 ), .A2(_add_98_n305 ), .ZN(_add_98_n131 ) );
INV_X4 _add_98_U357  ( .A(_add_98_n131 ), .ZN(_add_98_n209 ) );
INV_X4 _add_98_U356  ( .A(_add_98_n220 ), .ZN(_add_98_n303 ) );
NAND2_X2 _add_98_U355  ( .A1(rnd_q[129]), .A2(cv_q[129]), .ZN(_add_98_n137 ));
INV_X4 _add_98_U354  ( .A(_add_98_n137 ), .ZN(_add_98_n261 ) );
INV_X4 _add_98_U353  ( .A(_add_98_n215 ), .ZN(_add_98_n78 ) );
NAND2_X2 _add_98_U352  ( .A1(_add_98_n301 ), .A2(_add_98_n302 ), .ZN(_add_98_n298 ) );
NAND2_X2 _add_98_U351  ( .A1(rnd_q[133]), .A2(cv_q[133]), .ZN(_add_98_n294 ));
NAND2_X2 _add_98_U350  ( .A1(_add_98_n67 ), .A2(_add_98_n294 ), .ZN(_add_98_n293 ) );
NAND2_X2 _add_98_U349  ( .A1(_add_98_n224 ), .A2(_add_98_n293 ), .ZN(_add_98_n292 ) );
NAND2_X2 _add_98_U348  ( .A1(_add_98_n22 ), .A2(_add_98_n292 ), .ZN(_add_98_n290 ) );
NAND3_X2 _add_98_U347  ( .A1(_add_98_n290 ), .A2(_add_98_n3 ), .A3(_add_98_n291 ), .ZN(_add_98_n259 ) );
INV_X4 _add_98_U346  ( .A(_add_98_n259 ), .ZN(_add_98_n134 ) );
XNOR2_X2 _add_98_U345  ( .A(_add_98_n288 ), .B(_add_98_n89 ), .ZN(N45) );
INV_X4 _add_98_U344  ( .A(_add_98_n279 ), .ZN(_add_98_n287 ) );
NAND2_X2 _add_98_U343  ( .A1(_add_98_n89 ), .A2(_add_98_n287 ), .ZN(_add_98_n286 ) );
NAND2_X2 _add_98_U342  ( .A1(_add_98_n285 ), .A2(_add_98_n286 ), .ZN(_add_98_n283 ) );
NAND2_X2 _add_98_U341  ( .A1(rnd_q[145]), .A2(cv_q[145]), .ZN(_add_98_n280 ));
NAND2_X2 _add_98_U340  ( .A1(_add_98_n41 ), .A2(_add_98_n280 ), .ZN(_add_98_n284 ) );
XNOR2_X2 _add_98_U339  ( .A(_add_98_n283 ), .B(_add_98_n284 ), .ZN(N46) );
NAND2_X2 _add_98_U338  ( .A1(cv_q[144]), .A2(rnd_q[144]), .ZN(_add_98_n282 ));
NAND2_X2 _add_98_U337  ( .A1(_add_98_n40 ), .A2(_add_98_n280 ), .ZN(_add_98_n268 ) );
INV_X4 _add_98_U336  ( .A(_add_98_n268 ), .ZN(_add_98_n276 ) );
NAND2_X2 _add_98_U335  ( .A1(_add_98_n271 ), .A2(_add_98_n89 ), .ZN(_add_98_n277 ) );
NAND2_X2 _add_98_U334  ( .A1(_add_98_n276 ), .A2(_add_98_n277 ), .ZN(_add_98_n272 ) );
NAND2_X2 _add_98_U333  ( .A1(rnd_q[146]), .A2(cv_q[146]), .ZN(_add_98_n267 ));
INV_X4 _add_98_U332  ( .A(rnd_q[146]), .ZN(_add_98_n274 ) );
INV_X4 _add_98_U331  ( .A(cv_q[146]), .ZN(_add_98_n275 ) );
NAND2_X2 _add_98_U330  ( .A1(_add_98_n274 ), .A2(_add_98_n275 ), .ZN(_add_98_n269 ) );
NAND2_X2 _add_98_U329  ( .A1(_add_98_n267 ), .A2(_add_98_n269 ), .ZN(_add_98_n273 ) );
XNOR2_X2 _add_98_U328  ( .A(_add_98_n272 ), .B(_add_98_n273 ), .ZN(N47) );
INV_X4 _add_98_U327  ( .A(_add_98_n89 ), .ZN(_add_98_n270 ) );
NAND2_X2 _add_98_U326  ( .A1(_add_98_n271 ), .A2(_add_98_n269 ), .ZN(_add_98_n257 ) );
NAND2_X2 _add_98_U325  ( .A1(_add_98_n268 ), .A2(_add_98_n269 ), .ZN(_add_98_n266 ) );
NAND2_X2 _add_98_U324  ( .A1(_add_98_n266 ), .A2(_add_98_n267 ), .ZN(_add_98_n196 ) );
NAND2_X2 _add_98_U323  ( .A1(rnd_q[147]), .A2(cv_q[147]), .ZN(_add_98_n126 ));
INV_X4 _add_98_U322  ( .A(rnd_q[147]), .ZN(_add_98_n263 ) );
INV_X4 _add_98_U321  ( .A(cv_q[147]), .ZN(_add_98_n264 ) );
NAND2_X2 _add_98_U320  ( .A1(_add_98_n263 ), .A2(_add_98_n264 ), .ZN(_add_98_n195 ) );
XNOR2_X2 _add_98_U319  ( .A(_add_98_n262 ), .B(_add_98_n28 ), .ZN(N48) );
XNOR2_X2 _add_98_U318  ( .A(_add_98_n220 ), .B(_add_98_n260 ), .ZN(N30) );
INV_X4 _add_98_U317  ( .A(_add_98_n257 ), .ZN(_add_98_n256 ) );
NAND2_X2 _add_98_U316  ( .A1(_add_98_n256 ), .A2(_add_98_n195 ), .ZN(_add_98_n128 ) );
NAND2_X2 _add_98_U315  ( .A1(_add_98_n196 ), .A2(_add_98_n195 ), .ZN(_add_98_n125 ) );
NAND2_X2 _add_98_U314  ( .A1(_add_98_n125 ), .A2(_add_98_n126 ), .ZN(_add_98_n254 ) );
XNOR2_X2 _add_98_U313  ( .A(_add_98_n234 ), .B(_add_98_n252 ), .ZN(N49) );
NAND2_X2 _add_98_U312  ( .A1(rnd_q[149]), .A2(cv_q[149]), .ZN(_add_98_n201 ));
INV_X4 _add_98_U311  ( .A(_add_98_n201 ), .ZN(_add_98_n249 ) );
XNOR2_X2 _add_98_U310  ( .A(_add_98_n247 ), .B(_add_98_n248 ), .ZN(N50) );
INV_X4 _add_98_U309  ( .A(_add_98_n235 ), .ZN(_add_98_n244 ) );
INV_X4 _add_98_U308  ( .A(_add_98_n243 ), .ZN(_add_98_n242 ) );
NAND2_X2 _add_98_U307  ( .A1(_add_98_n202 ), .A2(_add_98_n201 ), .ZN(_add_98_n241 ) );
INV_X4 _add_98_U306  ( .A(rnd_q[150]), .ZN(_add_98_n238 ) );
INV_X4 _add_98_U305  ( .A(cv_q[150]), .ZN(_add_98_n239 ) );
NAND2_X2 _add_98_U304  ( .A1(_add_98_n238 ), .A2(_add_98_n239 ), .ZN(_add_98_n198 ) );
NAND2_X2 _add_98_U303  ( .A1(rnd_q[150]), .A2(cv_q[150]), .ZN(_add_98_n203 ));
XNOR2_X2 _add_98_U302  ( .A(_add_98_n237 ), .B(_add_98_n31 ), .ZN(N51) );
NAND2_X2 _add_98_U301  ( .A1(_add_98_n202 ), .A2(_add_98_n201 ), .ZN(_add_98_n236 ) );
NAND2_X2 _add_98_U300  ( .A1(_add_98_n236 ), .A2(_add_98_n198 ), .ZN(_add_98_n233 ) );
NAND2_X2 _add_98_U299  ( .A1(_add_98_n235 ), .A2(_add_98_n198 ), .ZN(_add_98_n228 ) );
INV_X4 _add_98_U298  ( .A(rnd_q[151]), .ZN(_add_98_n231 ) );
INV_X4 _add_98_U297  ( .A(cv_q[151]), .ZN(_add_98_n232 ) );
NAND2_X2 _add_98_U296  ( .A1(_add_98_n231 ), .A2(_add_98_n232 ), .ZN(_add_98_n199 ) );
NAND2_X2 _add_98_U295  ( .A1(rnd_q[151]), .A2(cv_q[151]), .ZN(_add_98_n151 ));
NAND2_X2 _add_98_U294  ( .A1(_add_98_n199 ), .A2(_add_98_n151 ), .ZN(_add_98_n230 ) );
XNOR2_X2 _add_98_U293  ( .A(_add_98_n229 ), .B(_add_98_n230 ), .ZN(N52) );
INV_X4 _add_98_U292  ( .A(_add_98_n228 ), .ZN(_add_98_n227 ) );
NAND2_X2 _add_98_U291  ( .A1(_add_98_n227 ), .A2(_add_98_n199 ), .ZN(_add_98_n146 ) );
NAND2_X2 _add_98_U290  ( .A1(rnd_q[133]), .A2(cv_q[133]), .ZN(_add_98_n226 ));
NAND2_X2 _add_98_U289  ( .A1(_add_98_n67 ), .A2(_add_98_n226 ), .ZN(_add_98_n225 ) );
NAND2_X2 _add_98_U288  ( .A1(_add_98_n224 ), .A2(_add_98_n225 ), .ZN(_add_98_n223 ) );
NAND2_X2 _add_98_U287  ( .A1(_add_98_n22 ), .A2(_add_98_n223 ), .ZN(_add_98_n221 ) );
INV_X4 _add_98_U286  ( .A(_add_98_n214 ), .ZN(_add_98_n222 ) );
NAND4_X2 _add_98_U285  ( .A1(_add_98_n221 ), .A2(_add_98_n3 ), .A3(_add_98_n313 ), .A4(_add_98_n222 ), .ZN(_add_98_n206 ) );
NAND2_X2 _add_98_U284  ( .A1(rnd_q[129]), .A2(cv_q[129]), .ZN(_add_98_n219 ));
NAND2_X2 _add_98_U283  ( .A1(_add_98_n219 ), .A2(_add_98_n220 ), .ZN(_add_98_n218 ) );
NAND2_X2 _add_98_U282  ( .A1(_add_98_n1 ), .A2(_add_98_n218 ), .ZN(_add_98_n216 ) );
NAND2_X2 _add_98_U281  ( .A1(_add_98_n204 ), .A2(_add_98_n205 ), .ZN(_add_98_n188 ) );
INV_X4 _add_98_U280  ( .A(_add_98_n145 ), .ZN(_add_98_n197 ) );
NAND2_X2 _add_98_U279  ( .A1(_add_98_n197 ), .A2(_add_98_n151 ), .ZN(_add_98_n190 ) );
INV_X4 _add_98_U278  ( .A(_add_98_n196 ), .ZN(_add_98_n193 ) );
INV_X4 _add_98_U277  ( .A(_add_98_n195 ), .ZN(_add_98_n194 ) );
NAND2_X2 _add_98_U276  ( .A1(_add_98_n188 ), .A2(_add_98_n189 ), .ZN(_add_98_n162 ) );
NAND2_X2 _add_98_U275  ( .A1(rnd_q[152]), .A2(cv_q[152]), .ZN(_add_98_n186 ));
NAND2_X2 _add_98_U274  ( .A1(_add_98_n186 ), .A2(_add_98_n171 ), .ZN(_add_98_n187 ) );
XNOR2_X2 _add_98_U273  ( .A(_add_98_n162 ), .B(_add_98_n187 ), .ZN(N53) );
INV_X4 _add_98_U272  ( .A(_add_98_n180 ), .ZN(_add_98_n171 ) );
NAND2_X2 _add_98_U271  ( .A1(_add_98_n171 ), .A2(_add_98_n162 ), .ZN(_add_98_n185 ) );
NAND2_X2 _add_98_U270  ( .A1(_add_98_n185 ), .A2(_add_98_n186 ), .ZN(_add_98_n181 ) );
NAND2_X2 _add_98_U269  ( .A1(rnd_q[153]), .A2(cv_q[153]), .ZN(_add_98_n160 ));
INV_X4 _add_98_U268  ( .A(rnd_q[153]), .ZN(_add_98_n183 ) );
INV_X4 _add_98_U267  ( .A(cv_q[153]), .ZN(_add_98_n184 ) );
NAND2_X2 _add_98_U266  ( .A1(_add_98_n183 ), .A2(_add_98_n184 ), .ZN(_add_98_n170 ) );
NAND2_X2 _add_98_U265  ( .A1(_add_98_n160 ), .A2(_add_98_n170 ), .ZN(_add_98_n182 ) );
XNOR2_X2 _add_98_U264  ( .A(_add_98_n181 ), .B(_add_98_n182 ), .ZN(N54) );
INV_X4 _add_98_U263  ( .A(_add_98_n162 ), .ZN(_add_98_n179 ) );
INV_X4 _add_98_U262  ( .A(_add_98_n170 ), .ZN(_add_98_n177 ) );
NAND2_X2 _add_98_U261  ( .A1(cv_q[152]), .A2(rnd_q[152]), .ZN(_add_98_n178 ));
NAND2_X2 _add_98_U260  ( .A1(_add_98_n8 ), .A2(_add_98_n160 ), .ZN(_add_98_n176 ) );
INV_X4 _add_98_U259  ( .A(rnd_q[154]), .ZN(_add_98_n173 ) );
INV_X4 _add_98_U258  ( .A(cv_q[154]), .ZN(_add_98_n174 ) );
NAND2_X2 _add_98_U257  ( .A1(_add_98_n173 ), .A2(_add_98_n174 ), .ZN(_add_98_n158 ) );
NAND2_X2 _add_98_U256  ( .A1(rnd_q[154]), .A2(cv_q[154]), .ZN(_add_98_n161 ));
XNOR2_X2 _add_98_U255  ( .A(_add_98_n172 ), .B(_add_98_n30 ), .ZN(N55) );
NAND2_X2 _add_98_U254  ( .A1(_add_98_n36 ), .A2(_add_98_n162 ), .ZN(_add_98_n167 ) );
NAND2_X2 _add_98_U253  ( .A1(_add_98_n169 ), .A2(_add_98_n158 ), .ZN(_add_98_n168 ) );
NAND2_X2 _add_98_U252  ( .A1(_add_98_n167 ), .A2(_add_98_n168 ), .ZN(_add_98_n163 ) );
INV_X4 _add_98_U251  ( .A(rnd_q[155]), .ZN(_add_98_n165 ) );
INV_X4 _add_98_U250  ( .A(cv_q[155]), .ZN(_add_98_n166 ) );
NAND2_X2 _add_98_U249  ( .A1(_add_98_n165 ), .A2(_add_98_n166 ), .ZN(_add_98_n149 ) );
NAND2_X2 _add_98_U248  ( .A1(rnd_q[155]), .A2(cv_q[155]), .ZN(_add_98_n157 ));
NAND2_X2 _add_98_U247  ( .A1(_add_98_n149 ), .A2(_add_98_n157 ), .ZN(_add_98_n164 ) );
XNOR2_X2 _add_98_U246  ( .A(_add_98_n163 ), .B(_add_98_n164 ), .ZN(N56) );
NAND2_X2 _add_98_U245  ( .A1(_add_98_n156 ), .A2(_add_98_n157 ), .ZN(_add_98_n152 ) );
INV_X4 _add_98_U244  ( .A(rnd_q[156]), .ZN(_add_98_n154 ) );
INV_X4 _add_98_U243  ( .A(cv_q[156]), .ZN(_add_98_n155 ) );
NAND2_X2 _add_98_U242  ( .A1(_add_98_n154 ), .A2(_add_98_n155 ), .ZN(_add_98_n150 ) );
NAND2_X2 _add_98_U241  ( .A1(rnd_q[156]), .A2(cv_q[156]), .ZN(_add_98_n102 ));
XNOR2_X2 _add_98_U240  ( .A(_add_98_n153 ), .B(_add_98_n32 ), .ZN(N57) );
INV_X4 _add_98_U239  ( .A(_add_98_n151 ), .ZN(_add_98_n148 ) );
INV_X4 _add_98_U238  ( .A(_add_98_n121 ), .ZN(_add_98_n105 ) );
INV_X4 _add_98_U237  ( .A(_add_98_n102 ), .ZN(_add_98_n147 ) );
INV_X4 _add_98_U236  ( .A(_add_98_n146 ), .ZN(_add_98_n104 ) );
INV_X4 _add_98_U235  ( .A(_add_98_n128 ), .ZN(_add_98_n88 ) );
NAND2_X2 _add_98_U234  ( .A1(_add_98_n125 ), .A2(_add_98_n126 ), .ZN(_add_98_n103 ) );
NAND2_X2 _add_98_U233  ( .A1(_add_98_n103 ), .A2(_add_98_n13 ), .ZN(_add_98_n144 ) );
NAND2_X2 _add_98_U232  ( .A1(_add_98_n145 ), .A2(_add_98_n105 ), .ZN(_add_98_n94 ) );
NAND4_X2 _add_98_U231  ( .A1(_add_98_n142 ), .A2(_add_98_n143 ), .A3(_add_98_n144 ), .A4(_add_98_n94 ), .ZN(_add_98_n138 ) );
NAND2_X2 _add_98_U230  ( .A1(rnd_q[157]), .A2(cv_q[157]), .ZN(_add_98_n92 ));
INV_X4 _add_98_U229  ( .A(rnd_q[157]), .ZN(_add_98_n140 ) );
INV_X4 _add_98_U228  ( .A(cv_q[157]), .ZN(_add_98_n141 ) );
NAND2_X2 _add_98_U227  ( .A1(_add_98_n140 ), .A2(_add_98_n141 ), .ZN(_add_98_n118 ) );
NAND2_X2 _add_98_U226  ( .A1(_add_98_n92 ), .A2(_add_98_n118 ), .ZN(_add_98_n139 ) );
XNOR2_X2 _add_98_U225  ( .A(_add_98_n138 ), .B(_add_98_n139 ), .ZN(N58) );
XNOR2_X2 _add_98_U224  ( .A(_add_98_n81 ), .B(_add_98_n135 ), .ZN(N31) );
INV_X4 _add_98_U223  ( .A(_add_98_n133 ), .ZN(_add_98_n129 ) );
NAND2_X2 _add_98_U222  ( .A1(_add_98_n131 ), .A2(_add_98_n132 ), .ZN(_add_98_n130 ) );
NAND2_X2 _add_98_U221  ( .A1(_add_98_n125 ), .A2(_add_98_n126 ), .ZN(_add_98_n124 ) );
NAND2_X2 _add_98_U220  ( .A1(_add_98_n104 ), .A2(_add_98_n118 ), .ZN(_add_98_n122 ) );
NAND2_X2 _add_98_U219  ( .A1(_add_98_n21 ), .A2(_add_98_n118 ), .ZN(_add_98_n114 ) );
INV_X4 _add_98_U218  ( .A(_add_98_n94 ), .ZN(_add_98_n119 ) );
NAND2_X2 _add_98_U217  ( .A1(_add_98_n119 ), .A2(_add_98_n118 ), .ZN(_add_98_n115 ) );
INV_X4 _add_98_U216  ( .A(_add_98_n118 ), .ZN(_add_98_n106 ) );
NAND2_X2 _add_98_U215  ( .A1(_add_98_n11 ), .A2(_add_98_n118 ), .ZN(_add_98_n117 ) );
NAND4_X2 _add_98_U214  ( .A1(_add_98_n114 ), .A2(_add_98_n115 ), .A3(_add_98_n116 ), .A4(_add_98_n117 ), .ZN(_add_98_n113 ) );
INV_X4 _add_98_U213  ( .A(rnd_q[158]), .ZN(_add_98_n110 ) );
INV_X4 _add_98_U212  ( .A(cv_q[158]), .ZN(_add_98_n111 ) );
NAND2_X2 _add_98_U211  ( .A1(rnd_q[158]), .A2(cv_q[158]), .ZN(_add_98_n101 ));
INV_X4 _add_98_U210  ( .A(_add_98_n101 ), .ZN(_add_98_n109 ) );
XNOR2_X2 _add_98_U209  ( .A(_add_98_n107 ), .B(_add_98_n108 ), .ZN(N59) );
NAND2_X2 _add_98_U208  ( .A1(_add_98_n12 ), .A2(_add_98_n103 ), .ZN(_add_98_n84 ) );
NAND2_X2 _add_98_U207  ( .A1(_add_98_n95 ), .A2(_add_98_n147 ), .ZN(_add_98_n100 ) );
NAND2_X2 _add_98_U206  ( .A1(_add_98_n100 ), .A2(_add_98_n101 ), .ZN(_add_98_n96 ) );
NAND2_X2 _add_98_U205  ( .A1(_add_98_n21 ), .A2(_add_98_n95 ), .ZN(_add_98_n98 ) );
NAND2_X2 _add_98_U204  ( .A1(_add_98_n11 ), .A2(_add_98_n95 ), .ZN(_add_98_n99 ) );
NAND2_X2 _add_98_U203  ( .A1(_add_98_n98 ), .A2(_add_98_n99 ), .ZN(_add_98_n97 ) );
INV_X4 _add_98_U202  ( .A(_add_98_n95 ), .ZN(_add_98_n93 ) );
NAND4_X2 _add_98_U201  ( .A1(_add_98_n84 ), .A2(_add_98_n85 ), .A3(_add_98_n86 ), .A4(_add_98_n87 ), .ZN(_add_98_n82 ) );
XNOR2_X2 _add_98_U200  ( .A(rnd_q[159]), .B(cv_q[159]), .ZN(_add_98_n83 ) );
XNOR2_X2 _add_98_U199  ( .A(_add_98_n82 ), .B(_add_98_n83 ), .ZN(N60) );
XNOR2_X2 _add_98_U198  ( .A(_add_98_n75 ), .B(_add_98_n76 ), .ZN(N32) );
INV_X4 _add_98_U197  ( .A(_add_98_n67 ), .ZN(_add_98_n73 ) );
XNOR2_X2 _add_98_U196  ( .A(_add_98_n35 ), .B(_add_98_n74 ), .ZN(N33) );
INV_X4 _add_98_U195  ( .A(_add_98_n64 ), .ZN(_add_98_n71 ) );
XNOR2_X2 _add_98_U194  ( .A(_add_98_n69 ), .B(_add_98_n70 ), .ZN(N34) );
NAND2_X2 _add_98_U193  ( .A1(rnd_q[134]), .A2(cv_q[134]), .ZN(_add_98_n59 ));
NAND2_X2 _add_98_U192  ( .A1(_add_98_n59 ), .A2(_add_98_n5 ), .ZN(_add_98_n62 ) );
NAND2_X2 _add_98_U191  ( .A1(_add_98_n35 ), .A2(_add_98_n67 ), .ZN(_add_98_n66 ) );
NAND2_X2 _add_98_U190  ( .A1(_add_98_n65 ), .A2(_add_98_n66 ), .ZN(_add_98_n63 ) );
NAND2_X2 _add_98_U189  ( .A1(_add_98_n63 ), .A2(_add_98_n64 ), .ZN(_add_98_n60 ) );
XNOR2_X2 _add_98_U188  ( .A(_add_98_n62 ), .B(_add_98_n60 ), .ZN(N35) );
NAND2_X2 _add_98_U187  ( .A1(_add_98_n60 ), .A2(_add_98_n5 ), .ZN(_add_98_n58 ) );
NAND2_X2 _add_98_U186  ( .A1(_add_98_n58 ), .A2(_add_98_n59 ), .ZN(_add_98_n55 ) );
NAND2_X2 _add_98_U185  ( .A1(_add_98_n57 ), .A2(_add_98_n3 ), .ZN(_add_98_n56 ) );
XNOR2_X2 _add_98_U184  ( .A(_add_98_n55 ), .B(_add_98_n56 ), .ZN(N36) );
INV_X4 _add_98_U183  ( .A(_add_98_n53 ), .ZN(_add_98_n46 ) );
XNOR2_X2 _add_98_U182  ( .A(_add_98_n51 ), .B(_add_98_n52 ), .ZN(N37) );
XNOR2_X2 _add_98_U181  ( .A(_add_98_n42 ), .B(_add_98_n43 ), .ZN(N38) );
NAND2_X2 _add_98_U180  ( .A1(_add_98_n259 ), .A2(_add_98_n133 ), .ZN(_add_98_n258 ) );
OR2_X2 _add_98_U179  ( .A1(cv_q[145]), .A2(rnd_q[145]), .ZN(_add_98_n41 ) );
NOR2_X2 _add_98_U178  ( .A1(_add_98_n20 ), .A2(_add_98_n109 ), .ZN(_add_98_n108 ) );
NOR2_X2 _add_98_U177  ( .A1(_add_98_n243 ), .A2(_add_98_n249 ), .ZN(_add_98_n248 ) );
NOR2_X2 _add_98_U176  ( .A1(_add_98_n317 ), .A2(_add_98_n15 ), .ZN(_add_98_n319 ) );
NOR2_X2 _add_98_U175  ( .A1(_add_98_n23 ), .A2(_add_98_n44 ), .ZN(_add_98_n43 ) );
NOR2_X2 _add_98_U174  ( .A1(_add_98_n71 ), .A2(_add_98_n68 ), .ZN(_add_98_n70 ) );
NOR2_X2 _add_98_U173  ( .A1(_add_98_n14 ), .A2(_add_98_n73 ), .ZN(_add_98_n74 ) );
NOR2_X2 _add_98_U172  ( .A1(_add_98_n77 ), .A2(_add_98_n78 ), .ZN(_add_98_n76 ) );
AND2_X2 _add_98_U171  ( .A1(cv_q[136]), .A2(rnd_q[136]), .ZN(_add_98_n353 ));
NOR2_X2 _add_98_U170  ( .A1(_add_98_n24 ), .A2(_add_98_n251 ), .ZN(_add_98_n252 ) );
NOR2_X2 _add_98_U169  ( .A1(_add_98_n47 ), .A2(_add_98_n46 ), .ZN(_add_98_n52 ) );
NOR2_X2 _add_98_U168  ( .A1(_add_98_n26 ), .A2(_add_98_n80 ), .ZN(_add_98_n135 ) );
NOR2_X2 _add_98_U167  ( .A1(_add_98_n261 ), .A2(_add_98_n136 ), .ZN(_add_98_n260 ) );
NOR2_X2 _add_98_U166  ( .A1(cv_q[145]), .A2(rnd_q[145]), .ZN(_add_98_n278 ));
NOR2_X2 _add_98_U165  ( .A1(_add_98_n278 ), .A2(_add_98_n279 ), .ZN(_add_98_n271 ) );
NOR2_X2 _add_98_U164  ( .A1(cv_q[137]), .A2(rnd_q[137]), .ZN(_add_98_n355 ));
NOR2_X2 _add_98_U163  ( .A1(cv_q[138]), .A2(rnd_q[138]), .ZN(_add_98_n356 ));
NOR2_X2 _add_98_U162  ( .A1(_add_98_n355 ), .A2(_add_98_n356 ), .ZN(_add_98_n354 ) );
NOR2_X2 _add_98_U161  ( .A1(cv_q[145]), .A2(rnd_q[145]), .ZN(_add_98_n281 ));
NOR2_X2 _add_98_U160  ( .A1(_add_98_n308 ), .A2(_add_98_n312 ), .ZN(_add_98_n310 ) );
NOR2_X2 _add_98_U159  ( .A1(cv_q[148]), .A2(rnd_q[148]), .ZN(_add_98_n246 ));
NOR2_X2 _add_98_U158  ( .A1(cv_q[149]), .A2(rnd_q[149]), .ZN(_add_98_n245 ));
NOR2_X2 _add_98_U157  ( .A1(_add_98_n245 ), .A2(_add_98_n246 ), .ZN(_add_98_n235 ) );
NOR2_X2 _add_98_U156  ( .A1(cv_q[133]), .A2(rnd_q[133]), .ZN(_add_98_n295 ));
NOR2_X2 _add_98_U155  ( .A1(cv_q[134]), .A2(rnd_q[134]), .ZN(_add_98_n296 ));
NOR2_X2 _add_98_U154  ( .A1(_add_98_n295 ), .A2(_add_98_n296 ), .ZN(_add_98_n224 ) );
NOR2_X2 _add_98_U153  ( .A1(cv_q[133]), .A2(rnd_q[133]), .ZN(_add_98_n388 ));
NOR2_X2 _add_98_U152  ( .A1(_add_98_n343 ), .A2(_add_98_n318 ), .ZN(_add_98_n342 ) );
NOR2_X2 _add_98_U151  ( .A1(cv_q[149]), .A2(rnd_q[149]), .ZN(_add_98_n243 ));
OR2_X2 _add_98_U150  ( .A1(_add_98_n281 ), .A2(_add_98_n282 ), .ZN(_add_98_n40 ) );
NAND3_X2 _add_98_U149  ( .A1(cv_q[148]), .A2(rnd_q[148]), .A3(_add_98_n242 ),.ZN(_add_98_n202 ) );
NOR2_X2 _add_98_U148  ( .A1(cv_q[130]), .A2(rnd_q[130]), .ZN(_add_98_n80 ));
NOR2_X2 _add_98_U147  ( .A1(cv_q[131]), .A2(rnd_q[131]), .ZN(_add_98_n77 ));
NOR2_X2 _add_98_U146  ( .A1(cv_q[129]), .A2(rnd_q[129]), .ZN(_add_98_n136 ));
NOR2_X2 _add_98_U145  ( .A1(cv_q[148]), .A2(rnd_q[148]), .ZN(_add_98_n251 ));
NOR2_X2 _add_98_U144  ( .A1(cv_q[144]), .A2(rnd_q[144]), .ZN(_add_98_n279 ));
NOR2_X2 _add_98_U143  ( .A1(cv_q[134]), .A2(rnd_q[134]), .ZN(_add_98_n61 ));
NOR2_X2 _add_98_U142  ( .A1(cv_q[152]), .A2(rnd_q[152]), .ZN(_add_98_n180 ));
NOR2_X2 _add_98_U141  ( .A1(cv_q[133]), .A2(rnd_q[133]), .ZN(_add_98_n68 ));
NOR2_X2 _add_98_U140  ( .A1(_add_98_n77 ), .A2(_add_98_n384 ), .ZN(_add_98_n217 ) );
NOR2_X2 _add_98_U139  ( .A1(cv_q[142]), .A2(rnd_q[142]), .ZN(_add_98_n308 ));
NOR3_X2 _add_98_U138  ( .A1(_add_98_n307 ), .A2(_add_98_n308 ), .A3(_add_98_n309 ), .ZN(_add_98_n306 ) );
NOR2_X2 _add_98_U137  ( .A1(cv_q[138]), .A2(rnd_q[138]), .ZN(_add_98_n351 ));
NOR2_X2 _add_98_U136  ( .A1(cv_q[136]), .A2(rnd_q[136]), .ZN(_add_98_n47 ));
NOR2_X2 _add_98_U135  ( .A1(cv_q[137]), .A2(rnd_q[137]), .ZN(_add_98_n44 ));
NOR2_X2 _add_98_U134  ( .A1(cv_q[140]), .A2(rnd_q[140]), .ZN(_add_98_n318 ));
NOR2_X2 _add_98_U133  ( .A1(cv_q[141]), .A2(rnd_q[141]), .ZN(_add_98_n309 ));
NOR2_X2 _add_98_U132  ( .A1(_add_98_n18 ), .A2(_add_98_n152 ), .ZN(_add_98_n153 ) );
NOR2_X2 _add_98_U131  ( .A1(_add_98_n347 ), .A2(_add_98_n348 ), .ZN(_add_98_n346 ) );
NAND3_X2 _add_98_U130  ( .A1(_add_98_n345 ), .A2(_add_98_n16 ), .A3(_add_98_n346 ), .ZN(_add_98_n315 ) );
NOR2_X2 _add_98_U129  ( .A1(_add_98_n303 ), .A2(_add_98_n217 ), .ZN(_add_98_n301 ) );
NAND3_X2 _add_98_U128  ( .A1(_add_98_n379 ), .A2(_add_98_n373 ), .A3(_add_98_n380 ), .ZN(_add_98_n371 ) );
NOR2_X2 _add_98_U127  ( .A1(_add_98_n23 ), .A2(_add_98_n391 ), .ZN(_add_98_n370 ) );
NAND3_X2 _add_98_U126  ( .A1(_add_98_n370 ), .A2(_add_98_n371 ), .A3(_add_98_n372 ), .ZN(_add_98_n368 ) );
NOR2_X2 _add_98_U125  ( .A1(_add_98_n96 ), .A2(_add_98_n97 ), .ZN(_add_98_n85 ) );
OR2_X4 _add_98_U124  ( .A1(_add_98_n106 ), .A2(_add_98_n102 ), .ZN(_add_98_n39 ) );
AND2_X2 _add_98_U123  ( .A1(_add_98_n92 ), .A2(_add_98_n39 ), .ZN(_add_98_n116 ) );
NAND3_X2 _add_98_U122  ( .A1(_add_98_n336 ), .A2(_add_98_n4 ), .A3(_add_98_n6 ), .ZN(_add_98_n335 ) );
NAND3_X2 _add_98_U121  ( .A1(_add_98_n29 ), .A2(_add_98_n329 ), .A3(_add_98_n335 ), .ZN(_add_98_n333 ) );
NOR2_X2 _add_98_U120  ( .A1(_add_98_n80 ), .A2(_add_98_n81 ), .ZN(_add_98_n79 ) );
NOR2_X2 _add_98_U119  ( .A1(_add_98_n79 ), .A2(_add_98_n26 ), .ZN(_add_98_n75 ) );
NOR2_X2 _add_98_U118  ( .A1(_add_98_n35 ), .A2(_add_98_n50 ), .ZN(_add_98_n49 ) );
NOR2_X2 _add_98_U117  ( .A1(_add_98_n49 ), .A2(_add_98_n19 ), .ZN(_add_98_n48 ) );
NOR2_X2 _add_98_U116  ( .A1(_add_98_n47 ), .A2(_add_98_n48 ), .ZN(_add_98_n45 ) );
NOR2_X2 _add_98_U115  ( .A1(_add_98_n45 ), .A2(_add_98_n46 ), .ZN(_add_98_n42 ) );
NOR2_X2 _add_98_U114  ( .A1(_add_98_n251 ), .A2(_add_98_n234 ), .ZN(_add_98_n250 ) );
NOR2_X2 _add_98_U113  ( .A1(_add_98_n250 ), .A2(_add_98_n24 ), .ZN(_add_98_n247 ) );
NOR2_X2 _add_98_U112  ( .A1(_add_98_n35 ), .A2(_add_98_n14 ), .ZN(_add_98_n72 ) );
NOR2_X2 _add_98_U111  ( .A1(_add_98_n72 ), .A2(_add_98_n73 ), .ZN(_add_98_n69 ) );
NOR3_X2 _add_98_U110  ( .A1(_add_98_n179 ), .A2(_add_98_n177 ), .A3(_add_98_n180 ), .ZN(_add_98_n175 ) );
NOR2_X2 _add_98_U109  ( .A1(_add_98_n175 ), .A2(_add_98_n176 ), .ZN(_add_98_n172 ) );
NOR2_X2 _add_98_U108  ( .A1(_add_98_n61 ), .A2(_add_98_n68 ), .ZN(_add_98_n376 ) );
NAND3_X2 _add_98_U107  ( .A1(_add_98_n313 ), .A2(_add_98_n314 ), .A3(_add_98_n315 ), .ZN(_add_98_n132 ) );
NOR2_X2 _add_98_U106  ( .A1(_add_98_n234 ), .A2(_add_98_n244 ), .ZN(_add_98_n240 ) );
NOR2_X2 _add_98_U105  ( .A1(_add_98_n240 ), .A2(_add_98_n241 ), .ZN(_add_98_n237 ) );
NOR3_X2 _add_98_U104  ( .A1(_add_98_n134 ), .A2(_add_98_n129 ), .A3(_add_98_n130 ), .ZN(_add_98_n127 ) );
NOR2_X2 _add_98_U103  ( .A1(_add_98_n127 ), .A2(_add_98_n128 ), .ZN(_add_98_n123 ) );
NOR2_X2 _add_98_U102  ( .A1(_add_98_n123 ), .A2(_add_98_n124 ), .ZN(_add_98_n120 ) );
NAND3_X2 _add_98_U101  ( .A1(_add_98_n201 ), .A2(_add_98_n202 ), .A3(_add_98_n203 ), .ZN(_add_98_n200 ) );
AND2_X4 _add_98_U100  ( .A1(_add_98_n198 ), .A2(_add_98_n199 ), .ZN(_add_98_n38 ) );
AND2_X2 _add_98_U99  ( .A1(_add_98_n200 ), .A2(_add_98_n38 ), .ZN(_add_98_n145 ) );
NOR2_X2 _add_98_U98  ( .A1(_add_98_n318 ), .A2(_add_98_n25 ), .ZN(_add_98_n324 ) );
NOR2_X2 _add_98_U97  ( .A1(_add_98_n44 ), .A2(_add_98_n53 ), .ZN(_add_98_n391 ) );
NOR2_X2 _add_98_U96  ( .A1(_add_98_n20 ), .A2(_add_98_n92 ), .ZN(_add_98_n91 ) );
NOR2_X2 _add_98_U95  ( .A1(_add_98_n146 ), .A2(_add_98_n126 ), .ZN(_add_98_n192 ) );
OR2_X4 _add_98_U94  ( .A1(_add_98_n136 ), .A2(_add_98_n220 ), .ZN(_add_98_n37 ) );
AND2_X2 _add_98_U93  ( .A1(_add_98_n137 ), .A2(_add_98_n37 ), .ZN(_add_98_n81 ) );
AND3_X2 _add_98_U92  ( .A1(_add_98_n170 ), .A2(_add_98_n158 ), .A3(_add_98_n171 ), .ZN(_add_98_n36 ) );
NAND3_X2 _add_98_U91  ( .A1(_add_98_n149 ), .A2(_add_98_n150 ), .A3(_add_98_n36 ), .ZN(_add_98_n121 ) );
NOR3_X2 _add_98_U90  ( .A1(_add_98_n193 ), .A2(_add_98_n146 ), .A3(_add_98_n194 ), .ZN(_add_98_n191 ) );
NOR2_X2 _add_98_U89  ( .A1(_add_98_n318 ), .A2(_add_98_n25 ), .ZN(_add_98_n336 ) );
NOR2_X2 _add_98_U88  ( .A1(_add_98_n47 ), .A2(_add_98_n44 ), .ZN(_add_98_n373 ) );
NOR2_X2 _add_98_U87  ( .A1(_add_98_n14 ), .A2(_add_98_n68 ), .ZN(_add_98_n65 ) );
NAND3_X2 _add_98_U86  ( .A1(_add_98_n215 ), .A2(_add_98_n216 ), .A3(_add_98_n382 ), .ZN(_add_98_n211 ) );
AND3_X2 _add_98_U85  ( .A1(_add_98_n382 ), .A2(_add_98_n215 ), .A3(_add_98_n381 ), .ZN(_add_98_n35 ) );
NAND3_X2 _add_98_U84  ( .A1(_add_98_n160 ), .A2(_add_98_n8 ), .A3(_add_98_n161 ), .ZN(_add_98_n159 ) );
NAND3_X2 _add_98_U83  ( .A1(_add_98_n158 ), .A2(_add_98_n149 ), .A3(_add_98_n159 ), .ZN(_add_98_n156 ) );
NOR2_X2 _add_98_U82  ( .A1(_add_98_n14 ), .A2(_add_98_n388 ), .ZN(_add_98_n387 ) );
NAND3_X2 _add_98_U81  ( .A1(_add_98_n3 ), .A2(_add_98_n5 ), .A3(_add_98_n387 ), .ZN(_add_98_n50 ) );
NOR3_X2 _add_98_U80  ( .A1(_add_98_n120 ), .A2(_add_98_n121 ), .A3(_add_98_n122 ), .ZN(_add_98_n112 ) );
NOR2_X2 _add_98_U79  ( .A1(_add_98_n112 ), .A2(_add_98_n113 ), .ZN(_add_98_n107 ) );
NOR2_X2 _add_98_U78  ( .A1(_add_98_n20 ), .A2(_add_98_n106 ), .ZN(_add_98_n95 ) );
NOR2_X2 _add_98_U77  ( .A1(_add_98_n209 ), .A2(_add_98_n210 ), .ZN(_add_98_n208 ) );
NAND3_X2 _add_98_U76  ( .A1(_add_98_n211 ), .A2(_add_98_n212 ), .A3(_add_98_n379 ), .ZN(_add_98_n207 ) );
NAND3_X2 _add_98_U75  ( .A1(_add_98_n207 ), .A2(_add_98_n208 ), .A3(_add_98_n206 ), .ZN(_add_98_n205 ) );
NAND3_X2 _add_98_U74  ( .A1(_add_98_n233 ), .A2(_add_98_n203 ), .A3(_add_98_n17 ), .ZN(_add_98_n229 ) );
NOR2_X2 _add_98_U73  ( .A1(_add_98_n213 ), .A2(_add_98_n214 ), .ZN(_add_98_n291 ) );
NAND3_X2 _add_98_U72  ( .A1(_add_98_n161 ), .A2(_add_98_n8 ), .A3(_add_98_n160 ), .ZN(_add_98_n169 ) );
NOR3_X2 _add_98_U71  ( .A1(_add_98_n258 ), .A2(_add_98_n210 ), .A3(_add_98_n209 ), .ZN(_add_98_n255 ) );
NOR2_X2 _add_98_U70  ( .A1(_add_98_n255 ), .A2(_add_98_n128 ), .ZN(_add_98_n253 ) );
NOR2_X2 _add_98_U69  ( .A1(_add_98_n253 ), .A2(_add_98_n254 ), .ZN(_add_98_n234 ) );
NOR3_X2 _add_98_U68  ( .A1(_add_98_n217 ), .A2(_add_98_n78 ), .A3(_add_98_n1 ), .ZN(_add_98_n300 ) );
NOR2_X2 _add_98_U67  ( .A1(_add_98_n317 ), .A2(_add_98_n318 ), .ZN(_add_98_n316 ) );
NAND3_X2 _add_98_U66  ( .A1(_add_98_n4 ), .A2(_add_98_n9 ), .A3(_add_98_n316 ), .ZN(_add_98_n213 ) );
OR3_X4 _add_98_U65  ( .A1(_add_98_n310 ), .A2(_add_98_n311 ), .A3(_add_98_n15 ), .ZN(_add_98_n34 ) );
OR2_X2 _add_98_U64  ( .A1(_add_98_n34 ), .A2(_add_98_n306 ), .ZN(_add_98_n304 ) );
NOR2_X2 _add_98_U63  ( .A1(_add_98_n351 ), .A2(_add_98_n361 ), .ZN(_add_98_n360 ) );
NAND3_X2 _add_98_U62  ( .A1(_add_98_n358 ), .A2(_add_98_n359 ), .A3(_add_98_n360 ), .ZN(_add_98_n214 ) );
NOR3_X2 _add_98_U61  ( .A1(_add_98_n190 ), .A2(_add_98_n191 ), .A3(_add_98_n192 ), .ZN(_add_98_n189 ) );
NOR2_X2 _add_98_U60  ( .A1(_add_98_n270 ), .A2(_add_98_n257 ), .ZN(_add_98_n265 ) );
NOR2_X2 _add_98_U59  ( .A1(_add_98_n265 ), .A2(_add_98_n196 ), .ZN(_add_98_n262 ) );
NOR2_X2 _add_98_U58  ( .A1(_add_98_n35 ), .A2(_add_98_n50 ), .ZN(_add_98_n54 ) );
NOR2_X2 _add_98_U57  ( .A1(_add_98_n54 ), .A2(_add_98_n19 ), .ZN(_add_98_n51 ) );
NOR2_X2 _add_98_U56  ( .A1(_add_98_n128 ), .A2(_add_98_n146 ), .ZN(_add_98_n204 ) );
NOR2_X2 _add_98_U55  ( .A1(_add_98_n35 ), .A2(_add_98_n50 ), .ZN(_add_98_n362 ) );
NOR2_X2 _add_98_U54  ( .A1(_add_98_n362 ), .A2(_add_98_n19 ), .ZN(_add_98_n357 ) );
NOR2_X2 _add_98_U53  ( .A1(_add_98_n357 ), .A2(_add_98_n214 ), .ZN(_add_98_n344 ) );
NOR2_X2 _add_98_U52  ( .A1(_add_98_n344 ), .A2(_add_98_n327 ), .ZN(_add_98_n341 ) );
NOR2_X2 _add_98_U51  ( .A1(_add_98_n93 ), .A2(_add_98_n94 ), .ZN(_add_98_n90 ) );
NOR2_X2 _add_98_U50  ( .A1(_add_98_n213 ), .A2(_add_98_n214 ), .ZN(_add_98_n212 ) );
NOR2_X2 _add_98_U49  ( .A1(_add_98_n324 ), .A2(_add_98_n325 ), .ZN(_add_98_n323 ) );
NOR3_X2 _add_98_U48  ( .A1(_add_98_n322 ), .A2(_add_98_n323 ), .A3(_add_98_n27 ), .ZN(_add_98_n321 ) );
NOR2_X2 _add_98_U47  ( .A1(_add_98_n311 ), .A2(_add_98_n321 ), .ZN(_add_98_n320 ) );
NOR2_X2 _add_98_U46  ( .A1(_add_98_n35 ), .A2(_add_98_n50 ), .ZN(_add_98_n326 ) );
NAND3_X2 _add_98_U45  ( .A1(_add_98_n89 ), .A2(_add_98_n13 ), .A3(_add_98_n88 ), .ZN(_add_98_n143 ) );
NOR3_X2 _add_98_U44  ( .A1(_add_98_n11 ), .A2(_add_98_n21 ), .A3(_add_98_n147 ), .ZN(_add_98_n142 ) );
NAND3_X2 _add_98_U43  ( .A1(_add_98_n88 ), .A2(_add_98_n89 ), .A3(_add_98_n12 ), .ZN(_add_98_n87 ) );
NOR2_X2 _add_98_U42  ( .A1(_add_98_n90 ), .A2(_add_98_n91 ), .ZN(_add_98_n86 ) );
NOR4_X2 _add_98_U41  ( .A1(_add_98_n326 ), .A2(_add_98_n327 ), .A3(_add_98_n19 ), .A4(_add_98_n325 ), .ZN(_add_98_n322 ) );
NOR2_X2 _add_98_U40  ( .A1(_add_98_n261 ), .A2(_add_98_n78 ), .ZN(_add_98_n302 ) );
NOR2_X2 _add_98_U39  ( .A1(_add_98_n50 ), .A2(_add_98_n300 ), .ZN(_add_98_n299 ) );
NOR2_X2 _add_98_U38  ( .A1(_add_98_n213 ), .A2(_add_98_n214 ), .ZN(_add_98_n297 ) );
NAND3_X2 _add_98_U37  ( .A1(_add_98_n297 ), .A2(_add_98_n298 ), .A3(_add_98_n299 ), .ZN(_add_98_n133 ) );
NOR2_X2 _add_98_U36  ( .A1(_add_98_n210 ), .A2(_add_98_n209 ), .ZN(_add_98_n289 ) );
NAND3_X2 _add_98_U35  ( .A1(_add_98_n289 ), .A2(_add_98_n133 ), .A3(_add_98_n259 ), .ZN(_add_98_n89 ) );
AND2_X4 _add_98_U34  ( .A1(_add_98_n383 ), .A2(_add_98_n220 ), .ZN(N29) );
AND2_X4 _add_98_U33  ( .A1(_add_98_n150 ), .A2(_add_98_n102 ), .ZN(_add_98_n32 ) );
AND2_X4 _add_98_U32  ( .A1(_add_98_n198 ), .A2(_add_98_n203 ), .ZN(_add_98_n31 ) );
AND2_X4 _add_98_U31  ( .A1(_add_98_n158 ), .A2(_add_98_n161 ), .ZN(_add_98_n30 ) );
OR2_X4 _add_98_U30  ( .A1(_add_98_n309 ), .A2(_add_98_n328 ), .ZN(_add_98_n29 ) );
AND2_X4 _add_98_U29  ( .A1(_add_98_n126 ), .A2(_add_98_n195 ), .ZN(_add_98_n28 ) );
OR2_X4 _add_98_U28  ( .A1(_add_98_n308 ), .A2(_add_98_n309 ), .ZN(_add_98_n27 ) );
AND2_X4 _add_98_U27  ( .A1(rnd_q[130]), .A2(cv_q[130]), .ZN(_add_98_n26 ) );
AND2_X4 _add_98_U26  ( .A1(_add_98_n214 ), .A2(_add_98_n340 ), .ZN(_add_98_n25 ) );
AND2_X4 _add_98_U25  ( .A1(rnd_q[148]), .A2(cv_q[148]), .ZN(_add_98_n24 ) );
AND2_X4 _add_98_U24  ( .A1(rnd_q[137]), .A2(cv_q[137]), .ZN(_add_98_n23 ) );
AND2_X4 _add_98_U23  ( .A1(_add_98_n57 ), .A2(_add_98_n378 ), .ZN(_add_98_n22 ) );
AND2_X4 _add_98_U22  ( .A1(_add_98_n148 ), .A2(_add_98_n105 ), .ZN(_add_98_n21 ) );
AND2_X4 _add_98_U21  ( .A1(_add_98_n110 ), .A2(_add_98_n111 ), .ZN(_add_98_n20 ) );
AND2_X4 _add_98_U20  ( .A1(_add_98_n374 ), .A2(_add_98_n3 ), .ZN(_add_98_n19 ) );
AND3_X4 _add_98_U19  ( .A1(_add_98_n36 ), .A2(_add_98_n149 ), .A3(_add_98_n162 ), .ZN(_add_98_n18 ) );
OR2_X4 _add_98_U18  ( .A1(_add_98_n234 ), .A2(_add_98_n228 ), .ZN(_add_98_n17 ) );
OR2_X4 _add_98_U17  ( .A1(_add_98_n351 ), .A2(_add_98_n352 ), .ZN(_add_98_n16 ) );
AND2_X4 _add_98_U16  ( .A1(rnd_q[143]), .A2(cv_q[143]), .ZN(_add_98_n15 ) );
AND2_X4 _add_98_U15  ( .A1(_add_98_n389 ), .A2(_add_98_n390 ), .ZN(_add_98_n14 ) );
AND2_X4 _add_98_U14  ( .A1(_add_98_n104 ), .A2(_add_98_n105 ), .ZN(_add_98_n13 ) );
AND3_X4 _add_98_U13  ( .A1(_add_98_n104 ), .A2(_add_98_n95 ), .A3(_add_98_n105 ), .ZN(_add_98_n12 ) );
AND2_X4 _add_98_U12  ( .A1(_add_98_n152 ), .A2(_add_98_n150 ), .ZN(_add_98_n11 ) );
OR2_X4 _add_98_U11  ( .A1(cv_q[130]), .A2(rnd_q[130]), .ZN(_add_98_n10 ) );
OR2_X4 _add_98_U10  ( .A1(cv_q[142]), .A2(rnd_q[142]), .ZN(_add_98_n9 ) );
OR2_X4 _add_98_U9  ( .A1(_add_98_n177 ), .A2(_add_98_n178 ), .ZN(_add_98_n8 ) );
OR2_X4 _add_98_U8  ( .A1(cv_q[131]), .A2(rnd_q[131]), .ZN(_add_98_n7 ) );
OR3_X4 _add_98_U7  ( .A1(_add_98_n326 ), .A2(_add_98_n19 ), .A3(_add_98_n327 ), .ZN(_add_98_n6 ) );
OR2_X4 _add_98_U6  ( .A1(cv_q[134]), .A2(rnd_q[134]), .ZN(_add_98_n5 ) );
OR2_X4 _add_98_U5  ( .A1(cv_q[141]), .A2(rnd_q[141]), .ZN(_add_98_n4 ) );
OR2_X4 _add_98_U4  ( .A1(cv_q[135]), .A2(rnd_q[135]), .ZN(_add_98_n3 ) );
OR2_X4 _add_98_U3  ( .A1(cv_q[129]), .A2(rnd_q[129]), .ZN(_add_98_n2 ) );
AND3_X4 _add_98_U2  ( .A1(_add_98_n10 ), .A2(_add_98_n7 ), .A3(_add_98_n2 ),.ZN(_add_98_n1 ) );
NAND2_X2 _add_98_4_U421  ( .A1(rnd_q[32]), .A2(cv_q[32]), .ZN(_add_98_4_n221 ) );
INV_X4 _add_98_4_U420  ( .A(_add_98_4_n352 ), .ZN(_add_98_4_n389 ) );
NAND2_X2 _add_98_4_U419  ( .A1(rnd_q[42]), .A2(cv_q[42]), .ZN(_add_98_4_n351 ) );
NAND2_X2 _add_98_4_U418  ( .A1(_add_98_4_n389 ), .A2(_add_98_4_n351 ), .ZN(_add_98_4_n368 ) );
NAND2_X2 _add_98_4_U417  ( .A1(rnd_q[40]), .A2(cv_q[40]), .ZN(_add_98_4_n52 ) );
INV_X4 _add_98_4_U416  ( .A(_add_98_4_n49 ), .ZN(_add_98_4_n378 ) );
NAND2_X2 _add_98_4_U415  ( .A1(rnd_q[33]), .A2(cv_q[33]), .ZN(_add_98_4_n385 ) );
NAND2_X2 _add_98_4_U414  ( .A1(_add_98_4_n385 ), .A2(_add_98_4_n221 ), .ZN(_add_98_4_n384 ) );
NAND2_X2 _add_98_4_U413  ( .A1(_add_98_4_n1 ), .A2(_add_98_4_n384 ), .ZN(_add_98_4_n380 ) );
NAND2_X2 _add_98_4_U412  ( .A1(cv_q[34]), .A2(rnd_q[34]), .ZN(_add_98_4_n383 ) );
INV_X4 _add_98_4_U411  ( .A(_add_98_4_n218 ), .ZN(_add_98_4_n381 ) );
NAND2_X2 _add_98_4_U410  ( .A1(rnd_q[35]), .A2(cv_q[35]), .ZN(_add_98_4_n216 ) );
INV_X4 _add_98_4_U409  ( .A(_add_98_4_n30 ), .ZN(_add_98_4_n379 ) );
NAND2_X2 _add_98_4_U408  ( .A1(rnd_q[39]), .A2(cv_q[39]), .ZN(_add_98_4_n56 ) );
NAND2_X2 _add_98_4_U407  ( .A1(rnd_q[38]), .A2(cv_q[38]), .ZN(_add_98_4_n377 ) );
NAND2_X2 _add_98_4_U406  ( .A1(rnd_q[36]), .A2(cv_q[36]), .ZN(_add_98_4_n66 ) );
NAND2_X2 _add_98_4_U405  ( .A1(rnd_q[37]), .A2(cv_q[37]), .ZN(_add_98_4_n63 ) );
NAND2_X2 _add_98_4_U404  ( .A1(_add_98_4_n66 ), .A2(_add_98_4_n63 ), .ZN(_add_98_4_n376 ) );
NAND2_X2 _add_98_4_U403  ( .A1(_add_98_4_n375 ), .A2(_add_98_4_n376 ), .ZN(_add_98_4_n374 ) );
NAND2_X2 _add_98_4_U402  ( .A1(_add_98_4_n35 ), .A2(_add_98_4_n374 ), .ZN(_add_98_4_n373 ) );
NAND2_X2 _add_98_4_U401  ( .A1(_add_98_4_n19 ), .A2(_add_98_4_n372 ), .ZN(_add_98_4_n371 ) );
XNOR2_X2 _add_98_4_U400  ( .A(_add_98_4_n368 ), .B(_add_98_4_n367 ), .ZN(N135) );
NAND2_X2 _add_98_4_U399  ( .A1(_add_98_4_n367 ), .A2(_add_98_4_n389 ), .ZN(_add_98_4_n366 ) );
NAND2_X2 _add_98_4_U398  ( .A1(_add_98_4_n366 ), .A2(_add_98_4_n351 ), .ZN(_add_98_4_n364 ) );
NAND2_X2 _add_98_4_U397  ( .A1(rnd_q[43]), .A2(cv_q[43]), .ZN(_add_98_4_n350 ) );
NAND2_X2 _add_98_4_U396  ( .A1(_add_98_4_n350 ), .A2(_add_98_4_n315 ), .ZN(_add_98_4_n365 ) );
XNOR2_X2 _add_98_4_U395  ( .A(_add_98_4_n364 ), .B(_add_98_4_n365 ), .ZN(N136) );
INV_X4 _add_98_4_U394  ( .A(_add_98_4_n43 ), .ZN(_add_98_4_n359 ) );
INV_X4 _add_98_4_U393  ( .A(_add_98_4_n46 ), .ZN(_add_98_4_n360 ) );
INV_X4 _add_98_4_U392  ( .A(_add_98_4_n315 ), .ZN(_add_98_4_n362 ) );
NAND2_X2 _add_98_4_U391  ( .A1(_add_98_4_n354 ), .A2(_add_98_4_n355 ), .ZN(_add_98_4_n346 ) );
NAND2_X2 _add_98_4_U390  ( .A1(cv_q[41]), .A2(rnd_q[41]), .ZN(_add_98_4_n353 ) );
INV_X4 _add_98_4_U389  ( .A(_add_98_4_n351 ), .ZN(_add_98_4_n348 ) );
INV_X4 _add_98_4_U388  ( .A(_add_98_4_n350 ), .ZN(_add_98_4_n349 ) );
NAND2_X2 _add_98_4_U387  ( .A1(_add_98_4_n316 ), .A2(_add_98_4_n315 ), .ZN(_add_98_4_n341 ) );
INV_X4 _add_98_4_U386  ( .A(_add_98_4_n341 ), .ZN(_add_98_4_n328 ) );
NAND2_X2 _add_98_4_U385  ( .A1(rnd_q[44]), .A2(cv_q[44]), .ZN(_add_98_4_n329 ) );
INV_X4 _add_98_4_U384  ( .A(_add_98_4_n329 ), .ZN(_add_98_4_n344 ) );
XNOR2_X2 _add_98_4_U383  ( .A(_add_98_4_n342 ), .B(_add_98_4_n343 ), .ZN(N137) );
NAND2_X2 _add_98_4_U382  ( .A1(_add_98_4_n337 ), .A2(_add_98_4_n7 ), .ZN(_add_98_4_n340 ) );
NAND2_X2 _add_98_4_U381  ( .A1(_add_98_4_n340 ), .A2(_add_98_4_n329 ), .ZN(_add_98_4_n338 ) );
NAND2_X2 _add_98_4_U380  ( .A1(rnd_q[45]), .A2(cv_q[45]), .ZN(_add_98_4_n330 ) );
NAND2_X2 _add_98_4_U379  ( .A1(_add_98_4_n330 ), .A2(_add_98_4_n4 ), .ZN(_add_98_4_n339 ) );
XNOR2_X2 _add_98_4_U378  ( .A(_add_98_4_n338 ), .B(_add_98_4_n339 ), .ZN(N138) );
NAND2_X2 _add_98_4_U377  ( .A1(rnd_q[46]), .A2(cv_q[46]), .ZN(_add_98_4_n331 ) );
NAND2_X2 _add_98_4_U376  ( .A1(_add_98_4_n10 ), .A2(_add_98_4_n331 ), .ZN(_add_98_4_n335 ) );
XNOR2_X2 _add_98_4_U375  ( .A(_add_98_4_n334 ), .B(_add_98_4_n335 ), .ZN(N139) );
INV_X4 _add_98_4_U374  ( .A(rnd_q[47]), .ZN(_add_98_4_n332 ) );
INV_X4 _add_98_4_U373  ( .A(cv_q[47]), .ZN(_add_98_4_n333 ) );
NAND2_X2 _add_98_4_U372  ( .A1(_add_98_4_n332 ), .A2(_add_98_4_n333 ), .ZN(_add_98_4_n306 ) );
INV_X4 _add_98_4_U371  ( .A(_add_98_4_n306 ), .ZN(_add_98_4_n318 ) );
INV_X4 _add_98_4_U370  ( .A(_add_98_4_n331 ), .ZN(_add_98_4_n312 ) );
NAND2_X2 _add_98_4_U369  ( .A1(_add_98_4_n329 ), .A2(_add_98_4_n330 ), .ZN(_add_98_4_n326 ) );
XNOR2_X2 _add_98_4_U368  ( .A(_add_98_4_n320 ), .B(_add_98_4_n321 ), .ZN(N140) );
NAND2_X2 _add_98_4_U367  ( .A1(rnd_q[48]), .A2(cv_q[48]), .ZN(_add_98_4_n287 ) );
NAND2_X2 _add_98_4_U366  ( .A1(_add_98_4_n287 ), .A2(_add_98_4_n289 ), .ZN(_add_98_4_n290 ) );
INV_X4 _add_98_4_U365  ( .A(_add_98_4_n214 ), .ZN(_add_98_4_n314 ) );
INV_X4 _add_98_4_U364  ( .A(_add_98_4_n133 ), .ZN(_add_98_4_n211 ) );
NAND2_X2 _add_98_4_U363  ( .A1(cv_q[45]), .A2(rnd_q[45]), .ZN(_add_98_4_n313 ) );
NAND2_X2 _add_98_4_U362  ( .A1(rnd_q[44]), .A2(cv_q[44]), .ZN(_add_98_4_n308 ) );
NAND2_X2 _add_98_4_U361  ( .A1(_add_98_4_n305 ), .A2(_add_98_4_n306 ), .ZN(_add_98_4_n132 ) );
INV_X4 _add_98_4_U360  ( .A(_add_98_4_n132 ), .ZN(_add_98_4_n210 ) );
NAND2_X2 _add_98_4_U359  ( .A1(rnd_q[33]), .A2(cv_q[33]), .ZN(_add_98_4_n138 ) );
INV_X4 _add_98_4_U358  ( .A(_add_98_4_n138 ), .ZN(_add_98_4_n262 ) );
INV_X4 _add_98_4_U357  ( .A(_add_98_4_n216 ), .ZN(_add_98_4_n77 ) );
NAND2_X2 _add_98_4_U356  ( .A1(_add_98_4_n303 ), .A2(_add_98_4_n304 ), .ZN(_add_98_4_n300 ) );
NAND2_X2 _add_98_4_U355  ( .A1(rnd_q[37]), .A2(cv_q[37]), .ZN(_add_98_4_n296 ) );
NAND2_X2 _add_98_4_U354  ( .A1(_add_98_4_n66 ), .A2(_add_98_4_n296 ), .ZN(_add_98_4_n295 ) );
NAND2_X2 _add_98_4_U353  ( .A1(_add_98_4_n225 ), .A2(_add_98_4_n295 ), .ZN(_add_98_4_n294 ) );
NAND2_X2 _add_98_4_U352  ( .A1(_add_98_4_n35 ), .A2(_add_98_4_n294 ), .ZN(_add_98_4_n292 ) );
NAND3_X2 _add_98_4_U351  ( .A1(_add_98_4_n292 ), .A2(_add_98_4_n3 ), .A3(_add_98_4_n293 ), .ZN(_add_98_4_n260 ) );
INV_X4 _add_98_4_U350  ( .A(_add_98_4_n260 ), .ZN(_add_98_4_n135 ) );
XNOR2_X2 _add_98_4_U349  ( .A(_add_98_4_n290 ), .B(_add_98_4_n88 ), .ZN(N141) );
INV_X4 _add_98_4_U348  ( .A(_add_98_4_n281 ), .ZN(_add_98_4_n289 ) );
NAND2_X2 _add_98_4_U347  ( .A1(_add_98_4_n88 ), .A2(_add_98_4_n289 ), .ZN(_add_98_4_n288 ) );
NAND2_X2 _add_98_4_U346  ( .A1(_add_98_4_n287 ), .A2(_add_98_4_n288 ), .ZN(_add_98_4_n285 ) );
NAND2_X2 _add_98_4_U345  ( .A1(rnd_q[49]), .A2(cv_q[49]), .ZN(_add_98_4_n282 ) );
NAND2_X2 _add_98_4_U344  ( .A1(_add_98_4_n37 ), .A2(_add_98_4_n282 ), .ZN(_add_98_4_n286 ) );
XNOR2_X2 _add_98_4_U343  ( .A(_add_98_4_n285 ), .B(_add_98_4_n286 ), .ZN(N142) );
NAND2_X2 _add_98_4_U342  ( .A1(cv_q[48]), .A2(rnd_q[48]), .ZN(_add_98_4_n284 ) );
NAND2_X2 _add_98_4_U341  ( .A1(_add_98_4_n34 ), .A2(_add_98_4_n282 ), .ZN(_add_98_4_n270 ) );
INV_X4 _add_98_4_U340  ( .A(_add_98_4_n270 ), .ZN(_add_98_4_n278 ) );
NAND2_X2 _add_98_4_U339  ( .A1(_add_98_4_n273 ), .A2(_add_98_4_n88 ), .ZN(_add_98_4_n279 ) );
NAND2_X2 _add_98_4_U338  ( .A1(_add_98_4_n278 ), .A2(_add_98_4_n279 ), .ZN(_add_98_4_n274 ) );
NAND2_X2 _add_98_4_U337  ( .A1(rnd_q[50]), .A2(cv_q[50]), .ZN(_add_98_4_n269 ) );
INV_X4 _add_98_4_U336  ( .A(rnd_q[50]), .ZN(_add_98_4_n276 ) );
INV_X4 _add_98_4_U335  ( .A(cv_q[50]), .ZN(_add_98_4_n277 ) );
NAND2_X2 _add_98_4_U334  ( .A1(_add_98_4_n276 ), .A2(_add_98_4_n277 ), .ZN(_add_98_4_n271 ) );
NAND2_X2 _add_98_4_U333  ( .A1(_add_98_4_n269 ), .A2(_add_98_4_n271 ), .ZN(_add_98_4_n275 ) );
XNOR2_X2 _add_98_4_U332  ( .A(_add_98_4_n274 ), .B(_add_98_4_n275 ), .ZN(N143) );
INV_X4 _add_98_4_U331  ( .A(_add_98_4_n88 ), .ZN(_add_98_4_n272 ) );
NAND2_X2 _add_98_4_U330  ( .A1(_add_98_4_n273 ), .A2(_add_98_4_n271 ), .ZN(_add_98_4_n258 ) );
NAND2_X2 _add_98_4_U329  ( .A1(_add_98_4_n270 ), .A2(_add_98_4_n271 ), .ZN(_add_98_4_n268 ) );
NAND2_X2 _add_98_4_U328  ( .A1(_add_98_4_n268 ), .A2(_add_98_4_n269 ), .ZN(_add_98_4_n197 ) );
NAND2_X2 _add_98_4_U327  ( .A1(rnd_q[51]), .A2(cv_q[51]), .ZN(_add_98_4_n127 ) );
INV_X4 _add_98_4_U326  ( .A(rnd_q[51]), .ZN(_add_98_4_n265 ) );
INV_X4 _add_98_4_U325  ( .A(cv_q[51]), .ZN(_add_98_4_n266 ) );
NAND2_X2 _add_98_4_U324  ( .A1(_add_98_4_n265 ), .A2(_add_98_4_n266 ), .ZN(_add_98_4_n196 ) );
XNOR2_X2 _add_98_4_U323  ( .A(_add_98_4_n264 ), .B(_add_98_4_n23 ), .ZN(N144) );
INV_X4 _add_98_4_U322  ( .A(_add_98_4_n221 ), .ZN(_add_98_4_n263 ) );
XNOR2_X2 _add_98_4_U321  ( .A(_add_98_4_n221 ), .B(_add_98_4_n261 ), .ZN(N126) );
INV_X4 _add_98_4_U320  ( .A(_add_98_4_n258 ), .ZN(_add_98_4_n257 ) );
NAND2_X2 _add_98_4_U319  ( .A1(_add_98_4_n257 ), .A2(_add_98_4_n196 ), .ZN(_add_98_4_n129 ) );
NAND2_X2 _add_98_4_U318  ( .A1(_add_98_4_n197 ), .A2(_add_98_4_n196 ), .ZN(_add_98_4_n126 ) );
NAND2_X2 _add_98_4_U317  ( .A1(_add_98_4_n126 ), .A2(_add_98_4_n127 ), .ZN(_add_98_4_n255 ) );
XNOR2_X2 _add_98_4_U316  ( .A(_add_98_4_n235 ), .B(_add_98_4_n253 ), .ZN(N145) );
NAND2_X2 _add_98_4_U315  ( .A1(rnd_q[53]), .A2(cv_q[53]), .ZN(_add_98_4_n202 ) );
INV_X4 _add_98_4_U314  ( .A(_add_98_4_n202 ), .ZN(_add_98_4_n250 ) );
XNOR2_X2 _add_98_4_U313  ( .A(_add_98_4_n248 ), .B(_add_98_4_n249 ), .ZN(N146) );
INV_X4 _add_98_4_U312  ( .A(_add_98_4_n236 ), .ZN(_add_98_4_n245 ) );
INV_X4 _add_98_4_U311  ( .A(_add_98_4_n244 ), .ZN(_add_98_4_n243 ) );
NAND2_X2 _add_98_4_U310  ( .A1(_add_98_4_n203 ), .A2(_add_98_4_n202 ), .ZN(_add_98_4_n242 ) );
INV_X4 _add_98_4_U309  ( .A(rnd_q[54]), .ZN(_add_98_4_n239 ) );
INV_X4 _add_98_4_U308  ( .A(cv_q[54]), .ZN(_add_98_4_n240 ) );
NAND2_X2 _add_98_4_U307  ( .A1(_add_98_4_n239 ), .A2(_add_98_4_n240 ), .ZN(_add_98_4_n199 ) );
NAND2_X2 _add_98_4_U306  ( .A1(rnd_q[54]), .A2(cv_q[54]), .ZN(_add_98_4_n204 ) );
XNOR2_X2 _add_98_4_U305  ( .A(_add_98_4_n238 ), .B(_add_98_4_n26 ), .ZN(N147) );
NAND2_X2 _add_98_4_U304  ( .A1(_add_98_4_n203 ), .A2(_add_98_4_n202 ), .ZN(_add_98_4_n237 ) );
NAND2_X2 _add_98_4_U303  ( .A1(_add_98_4_n237 ), .A2(_add_98_4_n199 ), .ZN(_add_98_4_n234 ) );
NAND2_X2 _add_98_4_U302  ( .A1(_add_98_4_n236 ), .A2(_add_98_4_n199 ), .ZN(_add_98_4_n229 ) );
INV_X4 _add_98_4_U301  ( .A(rnd_q[55]), .ZN(_add_98_4_n232 ) );
INV_X4 _add_98_4_U300  ( .A(cv_q[55]), .ZN(_add_98_4_n233 ) );
NAND2_X2 _add_98_4_U299  ( .A1(_add_98_4_n232 ), .A2(_add_98_4_n233 ), .ZN(_add_98_4_n200 ) );
NAND2_X2 _add_98_4_U298  ( .A1(rnd_q[55]), .A2(cv_q[55]), .ZN(_add_98_4_n152 ) );
NAND2_X2 _add_98_4_U297  ( .A1(_add_98_4_n200 ), .A2(_add_98_4_n152 ), .ZN(_add_98_4_n231 ) );
XNOR2_X2 _add_98_4_U296  ( .A(_add_98_4_n230 ), .B(_add_98_4_n231 ), .ZN(N148) );
INV_X4 _add_98_4_U295  ( .A(_add_98_4_n229 ), .ZN(_add_98_4_n228 ) );
NAND2_X2 _add_98_4_U294  ( .A1(_add_98_4_n228 ), .A2(_add_98_4_n200 ), .ZN(_add_98_4_n147 ) );
NAND2_X2 _add_98_4_U293  ( .A1(rnd_q[37]), .A2(cv_q[37]), .ZN(_add_98_4_n227 ) );
NAND2_X2 _add_98_4_U292  ( .A1(_add_98_4_n66 ), .A2(_add_98_4_n227 ), .ZN(_add_98_4_n226 ) );
NAND2_X2 _add_98_4_U291  ( .A1(_add_98_4_n225 ), .A2(_add_98_4_n226 ), .ZN(_add_98_4_n224 ) );
NAND2_X2 _add_98_4_U290  ( .A1(_add_98_4_n35 ), .A2(_add_98_4_n224 ), .ZN(_add_98_4_n222 ) );
INV_X4 _add_98_4_U289  ( .A(_add_98_4_n215 ), .ZN(_add_98_4_n223 ) );
NAND4_X2 _add_98_4_U288  ( .A1(_add_98_4_n222 ), .A2(_add_98_4_n3 ), .A3(_add_98_4_n314 ), .A4(_add_98_4_n223 ), .ZN(_add_98_4_n207 ) );
NAND2_X2 _add_98_4_U287  ( .A1(rnd_q[33]), .A2(cv_q[33]), .ZN(_add_98_4_n220 ) );
NAND2_X2 _add_98_4_U286  ( .A1(_add_98_4_n220 ), .A2(_add_98_4_n221 ), .ZN(_add_98_4_n219 ) );
NAND2_X2 _add_98_4_U285  ( .A1(_add_98_4_n1 ), .A2(_add_98_4_n219 ), .ZN(_add_98_4_n217 ) );
NAND2_X2 _add_98_4_U284  ( .A1(_add_98_4_n205 ), .A2(_add_98_4_n206 ), .ZN(_add_98_4_n189 ) );
INV_X4 _add_98_4_U283  ( .A(_add_98_4_n146 ), .ZN(_add_98_4_n198 ) );
NAND2_X2 _add_98_4_U282  ( .A1(_add_98_4_n198 ), .A2(_add_98_4_n152 ), .ZN(_add_98_4_n191 ) );
INV_X4 _add_98_4_U281  ( .A(_add_98_4_n197 ), .ZN(_add_98_4_n194 ) );
INV_X4 _add_98_4_U280  ( .A(_add_98_4_n196 ), .ZN(_add_98_4_n195 ) );
NAND2_X2 _add_98_4_U279  ( .A1(_add_98_4_n189 ), .A2(_add_98_4_n190 ), .ZN(_add_98_4_n163 ) );
NAND2_X2 _add_98_4_U278  ( .A1(rnd_q[56]), .A2(cv_q[56]), .ZN(_add_98_4_n187 ) );
NAND2_X2 _add_98_4_U277  ( .A1(_add_98_4_n187 ), .A2(_add_98_4_n172 ), .ZN(_add_98_4_n188 ) );
XNOR2_X2 _add_98_4_U276  ( .A(_add_98_4_n163 ), .B(_add_98_4_n188 ), .ZN(N149) );
INV_X4 _add_98_4_U275  ( .A(_add_98_4_n181 ), .ZN(_add_98_4_n172 ) );
NAND2_X2 _add_98_4_U274  ( .A1(_add_98_4_n172 ), .A2(_add_98_4_n163 ), .ZN(_add_98_4_n186 ) );
NAND2_X2 _add_98_4_U273  ( .A1(_add_98_4_n186 ), .A2(_add_98_4_n187 ), .ZN(_add_98_4_n182 ) );
NAND2_X2 _add_98_4_U272  ( .A1(rnd_q[57]), .A2(cv_q[57]), .ZN(_add_98_4_n161 ) );
INV_X4 _add_98_4_U271  ( .A(rnd_q[57]), .ZN(_add_98_4_n184 ) );
INV_X4 _add_98_4_U270  ( .A(cv_q[57]), .ZN(_add_98_4_n185 ) );
NAND2_X2 _add_98_4_U269  ( .A1(_add_98_4_n184 ), .A2(_add_98_4_n185 ), .ZN(_add_98_4_n171 ) );
NAND2_X2 _add_98_4_U268  ( .A1(_add_98_4_n161 ), .A2(_add_98_4_n171 ), .ZN(_add_98_4_n183 ) );
XNOR2_X2 _add_98_4_U267  ( .A(_add_98_4_n182 ), .B(_add_98_4_n183 ), .ZN(N150) );
INV_X4 _add_98_4_U266  ( .A(_add_98_4_n163 ), .ZN(_add_98_4_n180 ) );
INV_X4 _add_98_4_U265  ( .A(_add_98_4_n171 ), .ZN(_add_98_4_n178 ) );
NAND2_X2 _add_98_4_U264  ( .A1(cv_q[56]), .A2(rnd_q[56]), .ZN(_add_98_4_n179 ) );
NAND2_X2 _add_98_4_U263  ( .A1(_add_98_4_n9 ), .A2(_add_98_4_n161 ), .ZN(_add_98_4_n177 ) );
INV_X4 _add_98_4_U262  ( .A(rnd_q[58]), .ZN(_add_98_4_n174 ) );
INV_X4 _add_98_4_U261  ( .A(cv_q[58]), .ZN(_add_98_4_n175 ) );
NAND2_X2 _add_98_4_U260  ( .A1(_add_98_4_n174 ), .A2(_add_98_4_n175 ), .ZN(_add_98_4_n159 ) );
NAND2_X2 _add_98_4_U259  ( .A1(rnd_q[58]), .A2(cv_q[58]), .ZN(_add_98_4_n162 ) );
XNOR2_X2 _add_98_4_U258  ( .A(_add_98_4_n173 ), .B(_add_98_4_n25 ), .ZN(N151) );
NAND2_X2 _add_98_4_U257  ( .A1(_add_98_4_n31 ), .A2(_add_98_4_n163 ), .ZN(_add_98_4_n168 ) );
NAND2_X2 _add_98_4_U256  ( .A1(_add_98_4_n170 ), .A2(_add_98_4_n159 ), .ZN(_add_98_4_n169 ) );
NAND2_X2 _add_98_4_U255  ( .A1(_add_98_4_n168 ), .A2(_add_98_4_n169 ), .ZN(_add_98_4_n164 ) );
INV_X4 _add_98_4_U254  ( .A(rnd_q[59]), .ZN(_add_98_4_n166 ) );
INV_X4 _add_98_4_U253  ( .A(cv_q[59]), .ZN(_add_98_4_n167 ) );
NAND2_X2 _add_98_4_U252  ( .A1(_add_98_4_n166 ), .A2(_add_98_4_n167 ), .ZN(_add_98_4_n150 ) );
NAND2_X2 _add_98_4_U251  ( .A1(rnd_q[59]), .A2(cv_q[59]), .ZN(_add_98_4_n158 ) );
NAND2_X2 _add_98_4_U250  ( .A1(_add_98_4_n150 ), .A2(_add_98_4_n158 ), .ZN(_add_98_4_n165 ) );
XNOR2_X2 _add_98_4_U249  ( .A(_add_98_4_n164 ), .B(_add_98_4_n165 ), .ZN(N152) );
NAND2_X2 _add_98_4_U248  ( .A1(_add_98_4_n157 ), .A2(_add_98_4_n158 ), .ZN(_add_98_4_n153 ) );
INV_X4 _add_98_4_U247  ( .A(rnd_q[60]), .ZN(_add_98_4_n155 ) );
INV_X4 _add_98_4_U246  ( .A(cv_q[60]), .ZN(_add_98_4_n156 ) );
NAND2_X2 _add_98_4_U245  ( .A1(_add_98_4_n155 ), .A2(_add_98_4_n156 ), .ZN(_add_98_4_n151 ) );
NAND2_X2 _add_98_4_U244  ( .A1(rnd_q[60]), .A2(cv_q[60]), .ZN(_add_98_4_n101 ) );
XNOR2_X2 _add_98_4_U243  ( .A(_add_98_4_n154 ), .B(_add_98_4_n27 ), .ZN(N153) );
INV_X4 _add_98_4_U242  ( .A(_add_98_4_n152 ), .ZN(_add_98_4_n149 ) );
INV_X4 _add_98_4_U241  ( .A(_add_98_4_n122 ), .ZN(_add_98_4_n104 ) );
INV_X4 _add_98_4_U240  ( .A(_add_98_4_n101 ), .ZN(_add_98_4_n148 ) );
INV_X4 _add_98_4_U239  ( .A(_add_98_4_n147 ), .ZN(_add_98_4_n103 ) );
INV_X4 _add_98_4_U238  ( .A(_add_98_4_n129 ), .ZN(_add_98_4_n87 ) );
NAND2_X2 _add_98_4_U237  ( .A1(_add_98_4_n126 ), .A2(_add_98_4_n127 ), .ZN(_add_98_4_n102 ) );
NAND2_X2 _add_98_4_U236  ( .A1(_add_98_4_n102 ), .A2(_add_98_4_n13 ), .ZN(_add_98_4_n145 ) );
NAND2_X2 _add_98_4_U235  ( .A1(_add_98_4_n146 ), .A2(_add_98_4_n104 ), .ZN(_add_98_4_n93 ) );
NAND4_X2 _add_98_4_U234  ( .A1(_add_98_4_n143 ), .A2(_add_98_4_n144 ), .A3(_add_98_4_n145 ), .A4(_add_98_4_n93 ), .ZN(_add_98_4_n139 ) );
NAND2_X2 _add_98_4_U233  ( .A1(rnd_q[61]), .A2(cv_q[61]), .ZN(_add_98_4_n91 ) );
INV_X4 _add_98_4_U232  ( .A(rnd_q[61]), .ZN(_add_98_4_n141 ) );
INV_X4 _add_98_4_U231  ( .A(cv_q[61]), .ZN(_add_98_4_n142 ) );
NAND2_X2 _add_98_4_U230  ( .A1(_add_98_4_n141 ), .A2(_add_98_4_n142 ), .ZN(_add_98_4_n117 ) );
NAND2_X2 _add_98_4_U229  ( .A1(_add_98_4_n91 ), .A2(_add_98_4_n117 ), .ZN(_add_98_4_n140 ) );
XNOR2_X2 _add_98_4_U228  ( .A(_add_98_4_n139 ), .B(_add_98_4_n140 ), .ZN(N154) );
XNOR2_X2 _add_98_4_U227  ( .A(_add_98_4_n80 ), .B(_add_98_4_n136 ), .ZN(N127) );
INV_X4 _add_98_4_U226  ( .A(_add_98_4_n134 ), .ZN(_add_98_4_n130 ) );
NAND2_X2 _add_98_4_U225  ( .A1(_add_98_4_n132 ), .A2(_add_98_4_n133 ), .ZN(_add_98_4_n131 ) );
NAND2_X2 _add_98_4_U224  ( .A1(_add_98_4_n126 ), .A2(_add_98_4_n127 ), .ZN(_add_98_4_n125 ) );
NAND2_X2 _add_98_4_U223  ( .A1(_add_98_4_n103 ), .A2(_add_98_4_n117 ), .ZN(_add_98_4_n123 ) );
NAND2_X2 _add_98_4_U222  ( .A1(_add_98_4_n21 ), .A2(_add_98_4_n117 ), .ZN(_add_98_4_n113 ) );
INV_X4 _add_98_4_U221  ( .A(_add_98_4_n93 ), .ZN(_add_98_4_n120 ) );
NAND2_X2 _add_98_4_U220  ( .A1(_add_98_4_n120 ), .A2(_add_98_4_n117 ), .ZN(_add_98_4_n114 ) );
INV_X4 _add_98_4_U219  ( .A(_add_98_4_n91 ), .ZN(_add_98_4_n118 ) );
INV_X4 _add_98_4_U218  ( .A(_add_98_4_n117 ), .ZN(_add_98_4_n105 ) );
NAND2_X2 _add_98_4_U217  ( .A1(_add_98_4_n11 ), .A2(_add_98_4_n117 ), .ZN(_add_98_4_n116 ) );
NAND4_X2 _add_98_4_U216  ( .A1(_add_98_4_n113 ), .A2(_add_98_4_n114 ), .A3(_add_98_4_n115 ), .A4(_add_98_4_n116 ), .ZN(_add_98_4_n112 ) );
INV_X4 _add_98_4_U215  ( .A(rnd_q[62]), .ZN(_add_98_4_n109 ) );
INV_X4 _add_98_4_U214  ( .A(cv_q[62]), .ZN(_add_98_4_n110 ) );
NAND2_X2 _add_98_4_U213  ( .A1(rnd_q[62]), .A2(cv_q[62]), .ZN(_add_98_4_n100 ) );
INV_X4 _add_98_4_U212  ( .A(_add_98_4_n100 ), .ZN(_add_98_4_n108 ) );
XNOR2_X2 _add_98_4_U211  ( .A(_add_98_4_n106 ), .B(_add_98_4_n107 ), .ZN(N155) );
NAND2_X2 _add_98_4_U210  ( .A1(_add_98_4_n12 ), .A2(_add_98_4_n102 ), .ZN(_add_98_4_n83 ) );
NAND2_X2 _add_98_4_U209  ( .A1(_add_98_4_n94 ), .A2(_add_98_4_n148 ), .ZN(_add_98_4_n99 ) );
NAND2_X2 _add_98_4_U208  ( .A1(_add_98_4_n99 ), .A2(_add_98_4_n100 ), .ZN(_add_98_4_n95 ) );
NAND2_X2 _add_98_4_U207  ( .A1(_add_98_4_n21 ), .A2(_add_98_4_n94 ), .ZN(_add_98_4_n97 ) );
NAND2_X2 _add_98_4_U206  ( .A1(_add_98_4_n11 ), .A2(_add_98_4_n94 ), .ZN(_add_98_4_n98 ) );
NAND2_X2 _add_98_4_U205  ( .A1(_add_98_4_n97 ), .A2(_add_98_4_n98 ), .ZN(_add_98_4_n96 ) );
INV_X4 _add_98_4_U204  ( .A(_add_98_4_n94 ), .ZN(_add_98_4_n92 ) );
NAND4_X2 _add_98_4_U203  ( .A1(_add_98_4_n83 ), .A2(_add_98_4_n84 ), .A3(_add_98_4_n85 ), .A4(_add_98_4_n86 ), .ZN(_add_98_4_n81 ) );
XNOR2_X2 _add_98_4_U202  ( .A(rnd_q[63]), .B(cv_q[63]), .ZN(_add_98_4_n82 ));
XNOR2_X2 _add_98_4_U201  ( .A(_add_98_4_n81 ), .B(_add_98_4_n82 ), .ZN(N156));
XNOR2_X2 _add_98_4_U200  ( .A(_add_98_4_n74 ), .B(_add_98_4_n75 ), .ZN(N128));
INV_X4 _add_98_4_U199  ( .A(_add_98_4_n66 ), .ZN(_add_98_4_n72 ) );
XNOR2_X2 _add_98_4_U198  ( .A(_add_98_4_n30 ), .B(_add_98_4_n73 ), .ZN(N129));
INV_X4 _add_98_4_U197  ( .A(_add_98_4_n63 ), .ZN(_add_98_4_n70 ) );
XNOR2_X2 _add_98_4_U196  ( .A(_add_98_4_n68 ), .B(_add_98_4_n69 ), .ZN(N130));
NAND2_X2 _add_98_4_U195  ( .A1(rnd_q[38]), .A2(cv_q[38]), .ZN(_add_98_4_n58 ) );
NAND2_X2 _add_98_4_U194  ( .A1(_add_98_4_n58 ), .A2(_add_98_4_n6 ), .ZN(_add_98_4_n61 ) );
NAND2_X2 _add_98_4_U193  ( .A1(_add_98_4_n30 ), .A2(_add_98_4_n66 ), .ZN(_add_98_4_n65 ) );
NAND2_X2 _add_98_4_U192  ( .A1(_add_98_4_n64 ), .A2(_add_98_4_n65 ), .ZN(_add_98_4_n62 ) );
NAND2_X2 _add_98_4_U191  ( .A1(_add_98_4_n62 ), .A2(_add_98_4_n63 ), .ZN(_add_98_4_n59 ) );
XNOR2_X2 _add_98_4_U190  ( .A(_add_98_4_n61 ), .B(_add_98_4_n59 ), .ZN(N131));
NAND2_X2 _add_98_4_U189  ( .A1(_add_98_4_n59 ), .A2(_add_98_4_n6 ), .ZN(_add_98_4_n57 ) );
NAND2_X2 _add_98_4_U188  ( .A1(_add_98_4_n57 ), .A2(_add_98_4_n58 ), .ZN(_add_98_4_n54 ) );
NAND2_X2 _add_98_4_U187  ( .A1(_add_98_4_n56 ), .A2(_add_98_4_n3 ), .ZN(_add_98_4_n55 ) );
XNOR2_X2 _add_98_4_U186  ( .A(_add_98_4_n54 ), .B(_add_98_4_n55 ), .ZN(N132));
INV_X4 _add_98_4_U185  ( .A(_add_98_4_n52 ), .ZN(_add_98_4_n45 ) );
XNOR2_X2 _add_98_4_U184  ( .A(_add_98_4_n50 ), .B(_add_98_4_n51 ), .ZN(N133));
XNOR2_X2 _add_98_4_U183  ( .A(_add_98_4_n41 ), .B(_add_98_4_n42 ), .ZN(N134));
NAND2_X2 _add_98_4_U182  ( .A1(_add_98_4_n260 ), .A2(_add_98_4_n134 ), .ZN(_add_98_4_n259 ) );
NOR2_X2 _add_98_4_U181  ( .A1(_add_98_4_n20 ), .A2(_add_98_4_n108 ), .ZN(_add_98_4_n107 ) );
NOR2_X2 _add_98_4_U180  ( .A1(_add_98_4_n244 ), .A2(_add_98_4_n250 ), .ZN(_add_98_4_n249 ) );
AND2_X2 _add_98_4_U179  ( .A1(cv_q[40]), .A2(rnd_q[40]), .ZN(_add_98_4_n354 ) );
NOR2_X2 _add_98_4_U178  ( .A1(_add_98_4_n39 ), .A2(_add_98_4_n252 ), .ZN(_add_98_4_n253 ) );
NOR2_X2 _add_98_4_U177  ( .A1(_add_98_4_n40 ), .A2(_add_98_4_n43 ), .ZN(_add_98_4_n42 ) );
NOR2_X2 _add_98_4_U176  ( .A1(_add_98_4_n76 ), .A2(_add_98_4_n77 ), .ZN(_add_98_4_n75 ) );
NOR2_X2 _add_98_4_U175  ( .A1(_add_98_4_n262 ), .A2(_add_98_4_n137 ), .ZN(_add_98_4_n261 ) );
AND2_X2 _add_98_4_U174  ( .A1(rnd_q[41]), .A2(cv_q[41]), .ZN(_add_98_4_n40 ));
AND2_X2 _add_98_4_U173  ( .A1(rnd_q[52]), .A2(cv_q[52]), .ZN(_add_98_4_n39 ));
AND2_X2 _add_98_4_U172  ( .A1(rnd_q[34]), .A2(cv_q[34]), .ZN(_add_98_4_n38 ));
OR2_X2 _add_98_4_U171  ( .A1(cv_q[49]), .A2(rnd_q[49]), .ZN(_add_98_4_n37 ));
NOR2_X2 _add_98_4_U170  ( .A1(cv_q[49]), .A2(rnd_q[49]), .ZN(_add_98_4_n280 ) );
NOR2_X2 _add_98_4_U169  ( .A1(_add_98_4_n280 ), .A2(_add_98_4_n281 ), .ZN(_add_98_4_n273 ) );
NOR2_X2 _add_98_4_U168  ( .A1(cv_q[37]), .A2(rnd_q[37]), .ZN(_add_98_4_n297 ) );
NOR2_X2 _add_98_4_U167  ( .A1(cv_q[38]), .A2(rnd_q[38]), .ZN(_add_98_4_n298 ) );
NOR2_X2 _add_98_4_U166  ( .A1(_add_98_4_n297 ), .A2(_add_98_4_n298 ), .ZN(_add_98_4_n225 ) );
NOR2_X2 _add_98_4_U165  ( .A1(rnd_q[36]), .A2(cv_q[36]), .ZN(_add_98_4_n36 ));
NOR2_X2 _add_98_4_U164  ( .A1(cv_q[41]), .A2(rnd_q[41]), .ZN(_add_98_4_n356 ) );
NOR2_X2 _add_98_4_U163  ( .A1(_add_98_4_n356 ), .A2(_add_98_4_n357 ), .ZN(_add_98_4_n355 ) );
AND2_X2 _add_98_4_U162  ( .A1(_add_98_4_n56 ), .A2(_add_98_4_n377 ), .ZN(_add_98_4_n35 ) );
NOR2_X2 _add_98_4_U161  ( .A1(cv_q[49]), .A2(rnd_q[49]), .ZN(_add_98_4_n283 ) );
NOR2_X2 _add_98_4_U160  ( .A1(_add_98_4_n309 ), .A2(_add_98_4_n313 ), .ZN(_add_98_4_n311 ) );
NOR2_X2 _add_98_4_U159  ( .A1(cv_q[52]), .A2(rnd_q[52]), .ZN(_add_98_4_n247 ) );
NOR2_X2 _add_98_4_U158  ( .A1(cv_q[53]), .A2(rnd_q[53]), .ZN(_add_98_4_n246 ) );
NOR2_X2 _add_98_4_U157  ( .A1(_add_98_4_n246 ), .A2(_add_98_4_n247 ), .ZN(_add_98_4_n236 ) );
NOR2_X2 _add_98_4_U156  ( .A1(cv_q[37]), .A2(rnd_q[37]), .ZN(_add_98_4_n387 ) );
NOR2_X2 _add_98_4_U155  ( .A1(_add_98_4_n46 ), .A2(_add_98_4_n45 ), .ZN(_add_98_4_n51 ) );
NOR2_X2 _add_98_4_U154  ( .A1(_add_98_4_n38 ), .A2(_add_98_4_n79 ), .ZN(_add_98_4_n136 ) );
NOR2_X2 _add_98_4_U153  ( .A1(_add_98_4_n344 ), .A2(_add_98_4_n319 ), .ZN(_add_98_4_n343 ) );
NOR2_X2 _add_98_4_U152  ( .A1(_add_98_4_n70 ), .A2(_add_98_4_n67 ), .ZN(_add_98_4_n69 ) );
NOR2_X2 _add_98_4_U151  ( .A1(_add_98_4_n318 ), .A2(_add_98_4_n16 ), .ZN(_add_98_4_n320 ) );
NOR2_X2 _add_98_4_U150  ( .A1(_add_98_4_n36 ), .A2(_add_98_4_n72 ), .ZN(_add_98_4_n73 ) );
NOR2_X2 _add_98_4_U149  ( .A1(cv_q[53]), .A2(rnd_q[53]), .ZN(_add_98_4_n244 ) );
OR2_X2 _add_98_4_U148  ( .A1(_add_98_4_n283 ), .A2(_add_98_4_n284 ), .ZN(_add_98_4_n34 ) );
NAND3_X2 _add_98_4_U147  ( .A1(cv_q[52]), .A2(rnd_q[52]), .A3(_add_98_4_n243 ), .ZN(_add_98_4_n203 ) );
NOR2_X2 _add_98_4_U146  ( .A1(cv_q[52]), .A2(rnd_q[52]), .ZN(_add_98_4_n252 ) );
NOR2_X2 _add_98_4_U145  ( .A1(cv_q[33]), .A2(rnd_q[33]), .ZN(_add_98_4_n137 ) );
NOR2_X2 _add_98_4_U144  ( .A1(cv_q[48]), .A2(rnd_q[48]), .ZN(_add_98_4_n281 ) );
NOR2_X2 _add_98_4_U143  ( .A1(cv_q[38]), .A2(rnd_q[38]), .ZN(_add_98_4_n60 ));
NOR2_X2 _add_98_4_U142  ( .A1(cv_q[56]), .A2(rnd_q[56]), .ZN(_add_98_4_n181 ) );
NOR2_X2 _add_98_4_U141  ( .A1(cv_q[37]), .A2(rnd_q[37]), .ZN(_add_98_4_n67 ));
NOR2_X2 _add_98_4_U140  ( .A1(_add_98_4_n76 ), .A2(_add_98_4_n383 ), .ZN(_add_98_4_n218 ) );
NOR2_X2 _add_98_4_U139  ( .A1(cv_q[40]), .A2(rnd_q[40]), .ZN(_add_98_4_n46 ));
NOR2_X2 _add_98_4_U138  ( .A1(cv_q[41]), .A2(rnd_q[41]), .ZN(_add_98_4_n43 ));
NOR2_X2 _add_98_4_U137  ( .A1(cv_q[46]), .A2(rnd_q[46]), .ZN(_add_98_4_n309 ) );
NOR2_X2 _add_98_4_U136  ( .A1(cv_q[44]), .A2(rnd_q[44]), .ZN(_add_98_4_n319 ) );
NOR3_X2 _add_98_4_U135  ( .A1(_add_98_4_n308 ), .A2(_add_98_4_n309 ), .A3(_add_98_4_n310 ), .ZN(_add_98_4_n307 ) );
NOR2_X2 _add_98_4_U134  ( .A1(cv_q[45]), .A2(rnd_q[45]), .ZN(_add_98_4_n310 ) );
NAND3_X2 _add_98_4_U133  ( .A1(_add_98_4_n202 ), .A2(_add_98_4_n203 ), .A3(_add_98_4_n204 ), .ZN(_add_98_4_n201 ) );
AND2_X4 _add_98_4_U132  ( .A1(_add_98_4_n199 ), .A2(_add_98_4_n200 ), .ZN(_add_98_4_n33 ) );
AND2_X2 _add_98_4_U131  ( .A1(_add_98_4_n201 ), .A2(_add_98_4_n33 ), .ZN(_add_98_4_n146 ) );
NOR2_X2 _add_98_4_U130  ( .A1(_add_98_4_n348 ), .A2(_add_98_4_n349 ), .ZN(_add_98_4_n347 ) );
NAND3_X2 _add_98_4_U129  ( .A1(_add_98_4_n346 ), .A2(_add_98_4_n15 ), .A3(_add_98_4_n347 ), .ZN(_add_98_4_n316 ) );
NOR2_X2 _add_98_4_U128  ( .A1(_add_98_4_n263 ), .A2(_add_98_4_n218 ), .ZN(_add_98_4_n303 ) );
NAND3_X2 _add_98_4_U127  ( .A1(_add_98_4_n378 ), .A2(_add_98_4_n372 ), .A3(_add_98_4_n379 ), .ZN(_add_98_4_n370 ) );
NOR2_X2 _add_98_4_U126  ( .A1(_add_98_4_n40 ), .A2(_add_98_4_n388 ), .ZN(_add_98_4_n369 ) );
NAND3_X2 _add_98_4_U125  ( .A1(_add_98_4_n369 ), .A2(_add_98_4_n370 ), .A3(_add_98_4_n371 ), .ZN(_add_98_4_n367 ) );
NAND3_X2 _add_98_4_U124  ( .A1(_add_98_4_n337 ), .A2(_add_98_4_n4 ), .A3(_add_98_4_n7 ), .ZN(_add_98_4_n336 ) );
NAND3_X2 _add_98_4_U123  ( .A1(_add_98_4_n24 ), .A2(_add_98_4_n330 ), .A3(_add_98_4_n336 ), .ZN(_add_98_4_n334 ) );
NOR2_X2 _add_98_4_U122  ( .A1(_add_98_4_n79 ), .A2(_add_98_4_n80 ), .ZN(_add_98_4_n78 ) );
NOR2_X2 _add_98_4_U121  ( .A1(_add_98_4_n78 ), .A2(_add_98_4_n38 ), .ZN(_add_98_4_n74 ) );
NOR2_X2 _add_98_4_U120  ( .A1(_add_98_4_n18 ), .A2(_add_98_4_n153 ), .ZN(_add_98_4_n154 ) );
NOR2_X2 _add_98_4_U119  ( .A1(_add_98_4_n60 ), .A2(_add_98_4_n67 ), .ZN(_add_98_4_n375 ) );
NOR2_X2 _add_98_4_U118  ( .A1(_add_98_4_n235 ), .A2(_add_98_4_n245 ), .ZN(_add_98_4_n241 ) );
NOR2_X2 _add_98_4_U117  ( .A1(_add_98_4_n241 ), .A2(_add_98_4_n242 ), .ZN(_add_98_4_n238 ) );
NOR2_X2 _add_98_4_U116  ( .A1(_add_98_4_n30 ), .A2(_add_98_4_n49 ), .ZN(_add_98_4_n48 ) );
NOR2_X2 _add_98_4_U115  ( .A1(_add_98_4_n48 ), .A2(_add_98_4_n19 ), .ZN(_add_98_4_n47 ) );
NOR2_X2 _add_98_4_U114  ( .A1(_add_98_4_n46 ), .A2(_add_98_4_n47 ), .ZN(_add_98_4_n44 ) );
NOR2_X2 _add_98_4_U113  ( .A1(_add_98_4_n44 ), .A2(_add_98_4_n45 ), .ZN(_add_98_4_n41 ) );
NOR2_X2 _add_98_4_U112  ( .A1(_add_98_4_n252 ), .A2(_add_98_4_n235 ), .ZN(_add_98_4_n251 ) );
NOR2_X2 _add_98_4_U111  ( .A1(_add_98_4_n251 ), .A2(_add_98_4_n39 ), .ZN(_add_98_4_n248 ) );
NOR2_X2 _add_98_4_U110  ( .A1(_add_98_4_n30 ), .A2(_add_98_4_n36 ), .ZN(_add_98_4_n71 ) );
NOR2_X2 _add_98_4_U109  ( .A1(_add_98_4_n71 ), .A2(_add_98_4_n72 ), .ZN(_add_98_4_n68 ) );
NOR3_X2 _add_98_4_U108  ( .A1(_add_98_4_n180 ), .A2(_add_98_4_n178 ), .A3(_add_98_4_n181 ), .ZN(_add_98_4_n176 ) );
NOR2_X2 _add_98_4_U107  ( .A1(_add_98_4_n176 ), .A2(_add_98_4_n177 ), .ZN(_add_98_4_n173 ) );
NOR2_X2 _add_98_4_U106  ( .A1(_add_98_4_n36 ), .A2(_add_98_4_n67 ), .ZN(_add_98_4_n64 ) );
NAND3_X2 _add_98_4_U105  ( .A1(_add_98_4_n314 ), .A2(_add_98_4_n315 ), .A3(_add_98_4_n316 ), .ZN(_add_98_4_n133 ) );
NOR2_X2 _add_98_4_U104  ( .A1(_add_98_4_n20 ), .A2(_add_98_4_n91 ), .ZN(_add_98_4_n90 ) );
NOR2_X2 _add_98_4_U103  ( .A1(_add_98_4_n105 ), .A2(_add_98_4_n101 ), .ZN(_add_98_4_n119 ) );
NOR2_X2 _add_98_4_U102  ( .A1(_add_98_4_n319 ), .A2(_add_98_4_n14 ), .ZN(_add_98_4_n325 ) );
OR2_X4 _add_98_4_U101  ( .A1(_add_98_4_n137 ), .A2(_add_98_4_n221 ), .ZN(_add_98_4_n32 ) );
AND2_X2 _add_98_4_U100  ( .A1(_add_98_4_n138 ), .A2(_add_98_4_n32 ), .ZN(_add_98_4_n80 ) );
NOR2_X2 _add_98_4_U99  ( .A1(_add_98_4_n43 ), .A2(_add_98_4_n52 ), .ZN(_add_98_4_n388 ) );
NAND3_X2 _add_98_4_U98  ( .A1(_add_98_4_n161 ), .A2(_add_98_4_n9 ), .A3(_add_98_4_n162 ), .ZN(_add_98_4_n160 ) );
NAND3_X2 _add_98_4_U97  ( .A1(_add_98_4_n159 ), .A2(_add_98_4_n150 ), .A3(_add_98_4_n160 ), .ZN(_add_98_4_n157 ) );
NOR2_X2 _add_98_4_U96  ( .A1(_add_98_4_n147 ), .A2(_add_98_4_n127 ), .ZN(_add_98_4_n193 ) );
NOR3_X2 _add_98_4_U95  ( .A1(_add_98_4_n135 ), .A2(_add_98_4_n130 ), .A3(_add_98_4_n131 ), .ZN(_add_98_4_n128 ) );
NOR2_X2 _add_98_4_U94  ( .A1(_add_98_4_n128 ), .A2(_add_98_4_n129 ), .ZN(_add_98_4_n124 ) );
NOR2_X2 _add_98_4_U93  ( .A1(_add_98_4_n124 ), .A2(_add_98_4_n125 ), .ZN(_add_98_4_n121 ) );
NOR2_X2 _add_98_4_U92  ( .A1(_add_98_4_n318 ), .A2(_add_98_4_n319 ), .ZN(_add_98_4_n317 ) );
NAND3_X2 _add_98_4_U91  ( .A1(_add_98_4_n4 ), .A2(_add_98_4_n10 ), .A3(_add_98_4_n317 ), .ZN(_add_98_4_n214 ) );
AND3_X2 _add_98_4_U90  ( .A1(_add_98_4_n171 ), .A2(_add_98_4_n159 ), .A3(_add_98_4_n172 ), .ZN(_add_98_4_n31 ) );
NAND3_X2 _add_98_4_U89  ( .A1(_add_98_4_n150 ), .A2(_add_98_4_n151 ), .A3(_add_98_4_n31 ), .ZN(_add_98_4_n122 ) );
NOR3_X2 _add_98_4_U88  ( .A1(_add_98_4_n194 ), .A2(_add_98_4_n147 ), .A3(_add_98_4_n195 ), .ZN(_add_98_4_n192 ) );
NOR2_X2 _add_98_4_U87  ( .A1(_add_98_4_n319 ), .A2(_add_98_4_n14 ), .ZN(_add_98_4_n337 ) );
NOR2_X2 _add_98_4_U86  ( .A1(_add_98_4_n46 ), .A2(_add_98_4_n43 ), .ZN(_add_98_4_n372 ) );
NAND3_X2 _add_98_4_U85  ( .A1(_add_98_4_n216 ), .A2(_add_98_4_n217 ), .A3(_add_98_4_n381 ), .ZN(_add_98_4_n212 ) );
NOR2_X2 _add_98_4_U84  ( .A1(_add_98_4_n36 ), .A2(_add_98_4_n387 ), .ZN(_add_98_4_n386 ) );
NAND3_X2 _add_98_4_U83  ( .A1(_add_98_4_n3 ), .A2(_add_98_4_n6 ), .A3(_add_98_4_n386 ), .ZN(_add_98_4_n49 ) );
NOR2_X2 _add_98_4_U82  ( .A1(_add_98_4_n20 ), .A2(_add_98_4_n105 ), .ZN(_add_98_4_n94 ) );
AND3_X2 _add_98_4_U81  ( .A1(_add_98_4_n381 ), .A2(_add_98_4_n216 ), .A3(_add_98_4_n380 ), .ZN(_add_98_4_n30 ) );
OR3_X4 _add_98_4_U80  ( .A1(_add_98_4_n311 ), .A2(_add_98_4_n312 ), .A3(_add_98_4_n16 ), .ZN(_add_98_4_n29 ) );
OR2_X2 _add_98_4_U79  ( .A1(_add_98_4_n29 ), .A2(_add_98_4_n307 ), .ZN(_add_98_4_n305 ) );
NOR2_X2 _add_98_4_U78  ( .A1(_add_98_4_n210 ), .A2(_add_98_4_n211 ), .ZN(_add_98_4_n209 ) );
NAND3_X2 _add_98_4_U77  ( .A1(_add_98_4_n212 ), .A2(_add_98_4_n213 ), .A3(_add_98_4_n378 ), .ZN(_add_98_4_n208 ) );
NAND3_X2 _add_98_4_U76  ( .A1(_add_98_4_n208 ), .A2(_add_98_4_n209 ), .A3(_add_98_4_n207 ), .ZN(_add_98_4_n206 ) );
NAND3_X2 _add_98_4_U75  ( .A1(_add_98_4_n234 ), .A2(_add_98_4_n204 ), .A3(_add_98_4_n17 ), .ZN(_add_98_4_n230 ) );
NAND3_X2 _add_98_4_U74  ( .A1(_add_98_4_n162 ), .A2(_add_98_4_n9 ), .A3(_add_98_4_n161 ), .ZN(_add_98_4_n170 ) );
NOR3_X2 _add_98_4_U73  ( .A1(_add_98_4_n259 ), .A2(_add_98_4_n211 ), .A3(_add_98_4_n210 ), .ZN(_add_98_4_n256 ) );
NOR2_X2 _add_98_4_U72  ( .A1(_add_98_4_n256 ), .A2(_add_98_4_n129 ), .ZN(_add_98_4_n254 ) );
NOR2_X2 _add_98_4_U71  ( .A1(_add_98_4_n254 ), .A2(_add_98_4_n255 ), .ZN(_add_98_4_n235 ) );
NOR3_X2 _add_98_4_U70  ( .A1(_add_98_4_n218 ), .A2(_add_98_4_n77 ), .A3(_add_98_4_n1 ), .ZN(_add_98_4_n302 ) );
NOR2_X2 _add_98_4_U69  ( .A1(_add_98_4_n352 ), .A2(_add_98_4_n362 ), .ZN(_add_98_4_n361 ) );
NAND3_X2 _add_98_4_U68  ( .A1(_add_98_4_n359 ), .A2(_add_98_4_n360 ), .A3(_add_98_4_n361 ), .ZN(_add_98_4_n215 ) );
NOR2_X2 _add_98_4_U67  ( .A1(_add_98_4_n214 ), .A2(_add_98_4_n215 ), .ZN(_add_98_4_n293 ) );
NOR3_X2 _add_98_4_U66  ( .A1(_add_98_4_n191 ), .A2(_add_98_4_n192 ), .A3(_add_98_4_n193 ), .ZN(_add_98_4_n190 ) );
NOR2_X2 _add_98_4_U65  ( .A1(_add_98_4_n30 ), .A2(_add_98_4_n49 ), .ZN(_add_98_4_n363 ) );
NOR2_X2 _add_98_4_U64  ( .A1(_add_98_4_n363 ), .A2(_add_98_4_n19 ), .ZN(_add_98_4_n358 ) );
NOR2_X2 _add_98_4_U63  ( .A1(_add_98_4_n358 ), .A2(_add_98_4_n215 ), .ZN(_add_98_4_n345 ) );
NOR2_X2 _add_98_4_U62  ( .A1(_add_98_4_n345 ), .A2(_add_98_4_n328 ), .ZN(_add_98_4_n342 ) );
NOR2_X2 _add_98_4_U61  ( .A1(_add_98_4_n118 ), .A2(_add_98_4_n119 ), .ZN(_add_98_4_n115 ) );
NOR3_X2 _add_98_4_U60  ( .A1(_add_98_4_n121 ), .A2(_add_98_4_n122 ), .A3(_add_98_4_n123 ), .ZN(_add_98_4_n111 ) );
NOR2_X2 _add_98_4_U59  ( .A1(_add_98_4_n111 ), .A2(_add_98_4_n112 ), .ZN(_add_98_4_n106 ) );
NOR2_X2 _add_98_4_U58  ( .A1(_add_98_4_n30 ), .A2(_add_98_4_n49 ), .ZN(_add_98_4_n53 ) );
NOR2_X2 _add_98_4_U57  ( .A1(_add_98_4_n53 ), .A2(_add_98_4_n19 ), .ZN(_add_98_4_n50 ) );
NOR2_X2 _add_98_4_U56  ( .A1(_add_98_4_n272 ), .A2(_add_98_4_n258 ), .ZN(_add_98_4_n267 ) );
NOR2_X2 _add_98_4_U55  ( .A1(_add_98_4_n267 ), .A2(_add_98_4_n197 ), .ZN(_add_98_4_n264 ) );
NOR2_X2 _add_98_4_U54  ( .A1(_add_98_4_n129 ), .A2(_add_98_4_n147 ), .ZN(_add_98_4_n205 ) );
NOR2_X2 _add_98_4_U53  ( .A1(_add_98_4_n92 ), .A2(_add_98_4_n93 ), .ZN(_add_98_4_n89 ) );
NOR2_X2 _add_98_4_U52  ( .A1(_add_98_4_n214 ), .A2(_add_98_4_n215 ), .ZN(_add_98_4_n213 ) );
NOR2_X2 _add_98_4_U51  ( .A1(_add_98_4_n325 ), .A2(_add_98_4_n326 ), .ZN(_add_98_4_n324 ) );
NOR3_X2 _add_98_4_U50  ( .A1(_add_98_4_n323 ), .A2(_add_98_4_n324 ), .A3(_add_98_4_n22 ), .ZN(_add_98_4_n322 ) );
NOR2_X2 _add_98_4_U49  ( .A1(_add_98_4_n312 ), .A2(_add_98_4_n322 ), .ZN(_add_98_4_n321 ) );
NOR2_X2 _add_98_4_U48  ( .A1(_add_98_4_n30 ), .A2(_add_98_4_n49 ), .ZN(_add_98_4_n327 ) );
NAND3_X2 _add_98_4_U47  ( .A1(_add_98_4_n88 ), .A2(_add_98_4_n13 ), .A3(_add_98_4_n87 ), .ZN(_add_98_4_n144 ) );
NOR3_X2 _add_98_4_U46  ( .A1(_add_98_4_n11 ), .A2(_add_98_4_n21 ), .A3(_add_98_4_n148 ), .ZN(_add_98_4_n143 ) );
NOR2_X2 _add_98_4_U45  ( .A1(_add_98_4_n95 ), .A2(_add_98_4_n96 ), .ZN(_add_98_4_n84 ) );
NOR2_X2 _add_98_4_U44  ( .A1(_add_98_4_n89 ), .A2(_add_98_4_n90 ), .ZN(_add_98_4_n85 ) );
NOR4_X2 _add_98_4_U43  ( .A1(_add_98_4_n327 ), .A2(_add_98_4_n328 ), .A3(_add_98_4_n19 ), .A4(_add_98_4_n326 ), .ZN(_add_98_4_n323 ) );
NOR2_X2 _add_98_4_U42  ( .A1(_add_98_4_n262 ), .A2(_add_98_4_n77 ), .ZN(_add_98_4_n304 ) );
NOR2_X2 _add_98_4_U41  ( .A1(_add_98_4_n49 ), .A2(_add_98_4_n302 ), .ZN(_add_98_4_n301 ) );
NOR2_X2 _add_98_4_U40  ( .A1(_add_98_4_n214 ), .A2(_add_98_4_n215 ), .ZN(_add_98_4_n299 ) );
NAND3_X2 _add_98_4_U39  ( .A1(_add_98_4_n299 ), .A2(_add_98_4_n300 ), .A3(_add_98_4_n301 ), .ZN(_add_98_4_n134 ) );
NAND3_X2 _add_98_4_U38  ( .A1(_add_98_4_n87 ), .A2(_add_98_4_n88 ), .A3(_add_98_4_n12 ), .ZN(_add_98_4_n86 ) );
NOR2_X2 _add_98_4_U37  ( .A1(_add_98_4_n211 ), .A2(_add_98_4_n210 ), .ZN(_add_98_4_n291 ) );
NAND3_X2 _add_98_4_U36  ( .A1(_add_98_4_n291 ), .A2(_add_98_4_n134 ), .A3(_add_98_4_n260 ), .ZN(_add_98_4_n88 ) );
OR2_X4 _add_98_4_U35  ( .A1(rnd_q[32]), .A2(cv_q[32]), .ZN(_add_98_4_n382 ));
NOR2_X1 _add_98_4_U34  ( .A1(cv_q[42]), .A2(rnd_q[42]), .ZN(_add_98_4_n357 ));
NOR2_X1 _add_98_4_U33  ( .A1(cv_q[34]), .A2(rnd_q[34]), .ZN(_add_98_4_n79 ));
NOR2_X1 _add_98_4_U32  ( .A1(cv_q[35]), .A2(rnd_q[35]), .ZN(_add_98_4_n76 ));
OR2_X4 _add_98_4_U31  ( .A1(rnd_q[43]), .A2(cv_q[43]), .ZN(_add_98_4_n315 ));
NOR2_X1 _add_98_4_U30  ( .A1(cv_q[42]), .A2(rnd_q[42]), .ZN(_add_98_4_n352 ));
AND2_X4 _add_98_4_U29  ( .A1(_add_98_4_n382 ), .A2(_add_98_4_n221 ), .ZN(N125) );
AND2_X4 _add_98_4_U28  ( .A1(_add_98_4_n151 ), .A2(_add_98_4_n101 ), .ZN(_add_98_4_n27 ) );
AND2_X4 _add_98_4_U27  ( .A1(_add_98_4_n199 ), .A2(_add_98_4_n204 ), .ZN(_add_98_4_n26 ) );
AND2_X4 _add_98_4_U26  ( .A1(_add_98_4_n159 ), .A2(_add_98_4_n162 ), .ZN(_add_98_4_n25 ) );
OR2_X4 _add_98_4_U25  ( .A1(_add_98_4_n310 ), .A2(_add_98_4_n329 ), .ZN(_add_98_4_n24 ) );
AND2_X4 _add_98_4_U24  ( .A1(_add_98_4_n127 ), .A2(_add_98_4_n196 ), .ZN(_add_98_4_n23 ) );
OR2_X4 _add_98_4_U23  ( .A1(_add_98_4_n309 ), .A2(_add_98_4_n310 ), .ZN(_add_98_4_n22 ) );
AND2_X4 _add_98_4_U22  ( .A1(_add_98_4_n149 ), .A2(_add_98_4_n104 ), .ZN(_add_98_4_n21 ) );
AND2_X4 _add_98_4_U21  ( .A1(_add_98_4_n109 ), .A2(_add_98_4_n110 ), .ZN(_add_98_4_n20 ) );
AND2_X4 _add_98_4_U20  ( .A1(_add_98_4_n373 ), .A2(_add_98_4_n3 ), .ZN(_add_98_4_n19 ) );
AND3_X4 _add_98_4_U19  ( .A1(_add_98_4_n31 ), .A2(_add_98_4_n150 ), .A3(_add_98_4_n163 ), .ZN(_add_98_4_n18 ) );
OR2_X4 _add_98_4_U18  ( .A1(_add_98_4_n235 ), .A2(_add_98_4_n229 ), .ZN(_add_98_4_n17 ) );
AND2_X4 _add_98_4_U17  ( .A1(rnd_q[47]), .A2(cv_q[47]), .ZN(_add_98_4_n16 ));
OR2_X4 _add_98_4_U16  ( .A1(_add_98_4_n352 ), .A2(_add_98_4_n353 ), .ZN(_add_98_4_n15 ) );
AND2_X4 _add_98_4_U15  ( .A1(_add_98_4_n215 ), .A2(_add_98_4_n341 ), .ZN(_add_98_4_n14 ) );
AND2_X4 _add_98_4_U14  ( .A1(_add_98_4_n103 ), .A2(_add_98_4_n104 ), .ZN(_add_98_4_n13 ) );
AND3_X4 _add_98_4_U13  ( .A1(_add_98_4_n103 ), .A2(_add_98_4_n94 ), .A3(_add_98_4_n104 ), .ZN(_add_98_4_n12 ) );
AND2_X4 _add_98_4_U12  ( .A1(_add_98_4_n153 ), .A2(_add_98_4_n151 ), .ZN(_add_98_4_n11 ) );
OR2_X4 _add_98_4_U11  ( .A1(cv_q[46]), .A2(rnd_q[46]), .ZN(_add_98_4_n10 ));
OR2_X4 _add_98_4_U10  ( .A1(_add_98_4_n178 ), .A2(_add_98_4_n179 ), .ZN(_add_98_4_n9 ) );
OR2_X4 _add_98_4_U9  ( .A1(cv_q[33]), .A2(rnd_q[33]), .ZN(_add_98_4_n8 ) );
OR3_X4 _add_98_4_U8  ( .A1(_add_98_4_n327 ), .A2(_add_98_4_n19 ), .A3(_add_98_4_n328 ), .ZN(_add_98_4_n7 ) );
OR2_X4 _add_98_4_U7  ( .A1(cv_q[38]), .A2(rnd_q[38]), .ZN(_add_98_4_n6 ) );
OR2_X4 _add_98_4_U6  ( .A1(cv_q[35]), .A2(rnd_q[35]), .ZN(_add_98_4_n5 ) );
OR2_X4 _add_98_4_U5  ( .A1(cv_q[45]), .A2(rnd_q[45]), .ZN(_add_98_4_n4 ) );
OR2_X4 _add_98_4_U4  ( .A1(cv_q[39]), .A2(rnd_q[39]), .ZN(_add_98_4_n3 ) );
OR2_X4 _add_98_4_U3  ( .A1(cv_q[34]), .A2(rnd_q[34]), .ZN(_add_98_4_n2 ) );
AND3_X4 _add_98_4_U2  ( .A1(_add_98_4_n2 ), .A2(_add_98_4_n5 ), .A3(_add_98_4_n8 ), .ZN(_add_98_4_n1 ) );
endmodule
