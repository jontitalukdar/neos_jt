module s35932(blif_clk_net, blif_reset_net, DATA_0_31, DATA_0_30,DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24,DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18,DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12,DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7, DATA_0_6,DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2, DATA_0_1, DATA_0_0, RESET,TM1, TM0, DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27,DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21,DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15,DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9,DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3,DATA_9_2, DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1,CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11,CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15,CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19,CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23,CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27,CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31,CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4,CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9,CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17,CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21,CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25,CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29,CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2,CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7,CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11,CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19,CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23,CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27,CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31,CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4,CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9,CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13,CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21,CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25,CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29,CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2,CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7,CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11,CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15,CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27,CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31,CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4,CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9,CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13,CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17,CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21,CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29,CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2,CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7,CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11,CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15,CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19,CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23,CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31,CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4,CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9,CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13,CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17,CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21,CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25,CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2,CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11,CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15,CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19,CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23,CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27,CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31);
input blif_clk_net, blif_reset_net, DATA_0_31, DATA_0_30, DATA_0_29,DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24,DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19,DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14,DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8,DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2,DATA_0_1, DATA_0_0, RESET, TM1, TM0;
output DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27,DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22,DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17,DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12,DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6,DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2, DATA_9_1, DATA_9_0,CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4,CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9,CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13,CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17,CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21,CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29,CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1,CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6,CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10,CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14,CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26,CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30,CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2,CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7,CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11,CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19,CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23,CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27,CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31,CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4,CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9,CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13,CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21,CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25,CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29,CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1,CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6,CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10,CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18,CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22,CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26,CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30,CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2,CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7,CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11,CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15,CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19,CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23,CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27,CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31,CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4,CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9,CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17,CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21,CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25,CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29,CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1,CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6,CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10,CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14,CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18,CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22,CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26,CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30,CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2,CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11,CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15,CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19,CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23,CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27,CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31;
wire blif_clk_net, blif_reset_net, DATA_0_31, DATA_0_30, DATA_0_29,DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24,DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19,DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14,DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8,DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2,DATA_0_1, DATA_0_0, RESET, TM1, TM0;
wire DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27,DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22,DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17,DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12,DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6,DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2, DATA_9_1, DATA_9_0,CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4,CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9,CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13,CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17,CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21,CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29,CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1,CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6,CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10,CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14,CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26,CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30,CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2,CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7,CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11,CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19,CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23,CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27,CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31,CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4,CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9,CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13,CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21,CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25,CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29,CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1,CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6,CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10,CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18,CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22,CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26,CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30,CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2,CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7,CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11,CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15,CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19,CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23,CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27,CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31,CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4,CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9,CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17,CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21,CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25,CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29,CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1,CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6,CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10,CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14,CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18,CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22,CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26,CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30,CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2,CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11,CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15,CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19,CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23,CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27,CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31;
wire WX485, WX487, WX489, WX491, WX493, WX495, WX497, WX499;
wire WX501, WX503, WX505, WX507, WX509, WX511, WX513, WX515;
wire WX517, WX519, WX521, WX523, WX525, WX527, WX529, WX531;
wire WX533, WX535, WX537, WX539, WX541, WX543, WX545, WX547;
wire WX645, WX647, WX649, WX651, WX653, WX655, WX657, WX659;
wire WX661, WX663, WX665, WX667, WX669, WX671, WX673, WX675;
wire WX677, WX679, WX681, WX683, WX685, WX687, WX689, WX691;
wire WX693, WX695, WX697, WX699, WX701, WX703, WX705, WX707;
wire WX709, WX711, WX713, WX715, WX717, WX719, WX721, WX723;
wire WX725, WX727, WX729, WX731, WX733, WX735, WX737, WX739;
wire WX741, WX743, WX745, WX747, WX749, WX751, WX753, WX755;
wire WX757, WX759, WX761, WX763, WX765, WX767, WX769, WX771;
wire WX773, WX775, WX777, WX779, WX781, WX783, WX785, WX787;
wire WX789, WX791, WX793, WX795, WX797, WX799, WX801, WX803;
wire WX805, WX807, WX809, WX811, WX813, WX815, WX817, WX819;
wire WX821, WX823, WX825, WX827, WX829, WX831, WX833, WX835;
wire WX837, WX839, WX841, WX843, WX845, WX847, WX849, WX851;
wire WX853, WX855, WX857, WX859, WX861, WX863, WX865, WX867;
wire WX869, WX871, WX873, WX875, WX877, WX879, WX881, WX883;
wire WX885, WX887, WX889, WX891, WX893, WX895, WX897, WX899;
wire WX1778, WX1780, WX1782, WX1784, WX1786, WX1788, WX1790, WX1792;
wire WX1794, WX1796, WX1798, WX1800, WX1802, WX1804, WX1806, WX1808;
wire WX1810, WX1812, WX1814, WX1816, WX1818, WX1820, WX1822, WX1824;
wire WX1826, WX1828, WX1830, WX1832, WX1834, WX1836, WX1838, WX1840;
wire WX1938, WX1940, WX1942, WX1944, WX1946, WX1948, WX1950, WX1952;
wire WX1954, WX1956, WX1958, WX1960, WX1962, WX1964, WX1966, WX1968;
wire WX1970, WX1972, WX1974, WX1976, WX1978, WX1980, WX1982, WX1984;
wire WX1986, WX1988, WX1990, WX1992, WX1994, WX1996, WX1998, WX2000;
wire WX2002, WX2004, WX2006, WX2008, WX2010, WX2012, WX2014, WX2016;
wire WX2018, WX2020, WX2022, WX2024, WX2026, WX2028, WX2030, WX2032;
wire WX2034, WX2036, WX2038, WX2040, WX2042, WX2044, WX2046, WX2048;
wire WX2050, WX2052, WX2054, WX2056, WX2058, WX2060, WX2062, WX2064;
wire WX2066, WX2068, WX2070, WX2072, WX2074, WX2076, WX2078, WX2080;
wire WX2082, WX2084, WX2086, WX2088, WX2090, WX2092, WX2094, WX2096;
wire WX2098, WX2100, WX2102, WX2104, WX2106, WX2108, WX2110, WX2112;
wire WX2114, WX2116, WX2118, WX2120, WX2122, WX2124, WX2126, WX2128;
wire WX2130, WX2132, WX2134, WX2136, WX2138, WX2140, WX2142, WX2144;
wire WX2146, WX2148, WX2150, WX2152, WX2154, WX2156, WX2158, WX2160;
wire WX2162, WX2164, WX2166, WX2168, WX2170, WX2172, WX2174, WX2176;
wire WX2178, WX2180, WX2182, WX2184, WX2186, WX2188, WX2190, WX2192;
wire WX3071, WX3073, WX3075, WX3077, WX3079, WX3081, WX3083, WX3085;
wire WX3087, WX3089, WX3091, WX3093, WX3095, WX3097, WX3099, WX3101;
wire WX3103, WX3105, WX3107, WX3109, WX3111, WX3113, WX3115, WX3117;
wire WX3119, WX3121, WX3123, WX3125, WX3127, WX3129, WX3131, WX3133;
wire WX3231, WX3233, WX3235, WX3237, WX3239, WX3241, WX3243, WX3245;
wire WX3247, WX3249, WX3251, WX3253, WX3255, WX3257, WX3259, WX3261;
wire WX3263, WX3265, WX3267, WX3269, WX3271, WX3273, WX3275, WX3277;
wire WX3279, WX3281, WX3283, WX3285, WX3287, WX3289, WX3291, WX3293;
wire WX3295, WX3297, WX3299, WX3301, WX3303, WX3305, WX3307, WX3309;
wire WX3311, WX3313, WX3315, WX3317, WX3319, WX3321, WX3323, WX3325;
wire WX3327, WX3329, WX3331, WX3333, WX3335, WX3337, WX3339, WX3341;
wire WX3343, WX3345, WX3347, WX3349, WX3351, WX3353, WX3355, WX3357;
wire WX3359, WX3361, WX3363, WX3365, WX3367, WX3369, WX3371, WX3373;
wire WX3375, WX3377, WX3379, WX3381, WX3383, WX3385, WX3387, WX3389;
wire WX3391, WX3393, WX3395, WX3397, WX3399, WX3401, WX3403, WX3405;
wire WX3407, WX3409, WX3411, WX3413, WX3415, WX3417, WX3419, WX3421;
wire WX3423, WX3425, WX3427, WX3429, WX3431, WX3433, WX3435, WX3437;
wire WX3439, WX3441, WX3443, WX3445, WX3447, WX3449, WX3451, WX3453;
wire WX3455, WX3457, WX3459, WX3461, WX3463, WX3465, WX3467, WX3469;
wire WX3471, WX3473, WX3475, WX3477, WX3479, WX3481, WX3483, WX3485;
wire WX4364, WX4366, WX4368, WX4370, WX4372, WX4374, WX4376, WX4378;
wire WX4380, WX4382, WX4384, WX4386, WX4388, WX4390, WX4392, WX4394;
wire WX4396, WX4398, WX4400, WX4402, WX4404, WX4406, WX4408, WX4410;
wire WX4412, WX4414, WX4416, WX4418, WX4420, WX4422, WX4424, WX4426;
wire WX4524, WX4526, WX4528, WX4530, WX4532, WX4534, WX4536, WX4538;
wire WX4540, WX4542, WX4544, WX4546, WX4548, WX4550, WX4552, WX4554;
wire WX4556, WX4558, WX4560, WX4562, WX4564, WX4566, WX4568, WX4570;
wire WX4572, WX4574, WX4576, WX4578, WX4580, WX4582, WX4584, WX4586;
wire WX4588, WX4590, WX4592, WX4594, WX4596, WX4598, WX4600, WX4602;
wire WX4604, WX4606, WX4608, WX4610, WX4612, WX4614, WX4616, WX4618;
wire WX4620, WX4622, WX4624, WX4626, WX4628, WX4630, WX4632, WX4634;
wire WX4636, WX4638, WX4640, WX4642, WX4644, WX4646, WX4648, WX4650;
wire WX4652, WX4654, WX4656, WX4658, WX4660, WX4662, WX4664, WX4666;
wire WX4668, WX4670, WX4672, WX4674, WX4676, WX4678, WX4680, WX4682;
wire WX4684, WX4686, WX4688, WX4690, WX4692, WX4694, WX4696, WX4698;
wire WX4700, WX4702, WX4704, WX4706, WX4708, WX4710, WX4712, WX4714;
wire WX4716, WX4718, WX4720, WX4722, WX4724, WX4726, WX4728, WX4730;
wire WX4732, WX4734, WX4736, WX4738, WX4740, WX4742, WX4744, WX4746;
wire WX4748, WX4750, WX4752, WX4754, WX4756, WX4758, WX4760, WX4762;
wire WX4764, WX4766, WX4768, WX4770, WX4772, WX4774, WX4776, WX4778;
wire WX5657, WX5659, WX5661, WX5663, WX5665, WX5667, WX5669, WX5671;
wire WX5673, WX5675, WX5677, WX5679, WX5681, WX5683, WX5685, WX5687;
wire WX5689, WX5691, WX5693, WX5695, WX5697, WX5699, WX5701, WX5703;
wire WX5705, WX5707, WX5709, WX5711, WX5713, WX5715, WX5717, WX5719;
wire WX5817, WX5819, WX5821, WX5823, WX5825, WX5827, WX5829, WX5831;
wire WX5833, WX5835, WX5837, WX5839, WX5841, WX5843, WX5845, WX5847;
wire WX5849, WX5851, WX5853, WX5855, WX5857, WX5859, WX5861, WX5863;
wire WX5865, WX5867, WX5869, WX5871, WX5873, WX5875, WX5877, WX5879;
wire WX5881, WX5883, WX5885, WX5887, WX5889, WX5891, WX5893, WX5895;
wire WX5897, WX5899, WX5901, WX5903, WX5905, WX5907, WX5909, WX5911;
wire WX5913, WX5915, WX5917, WX5919, WX5921, WX5923, WX5925, WX5927;
wire WX5929, WX5931, WX5933, WX5935, WX5937, WX5939, WX5941, WX5943;
wire WX5945, WX5947, WX5949, WX5951, WX5953, WX5955, WX5957, WX5959;
wire WX5961, WX5963, WX5965, WX5967, WX5969, WX5971, WX5973, WX5975;
wire WX5977, WX5979, WX5981, WX5983, WX5985, WX5987, WX5989, WX5991;
wire WX5993, WX5995, WX5997, WX5999, WX6001, WX6003, WX6005, WX6007;
wire WX6009, WX6011, WX6013, WX6015, WX6017, WX6019, WX6021, WX6023;
wire WX6025, WX6027, WX6029, WX6031, WX6033, WX6035, WX6037, WX6039;
wire WX6041, WX6043, WX6045, WX6047, WX6049, WX6051, WX6053, WX6055;
wire WX6057, WX6059, WX6061, WX6063, WX6065, WX6067, WX6069, WX6071;
wire WX6950, WX6952, WX6954, WX6956, WX6958, WX6960, WX6962, WX6964;
wire WX6966, WX6968, WX6970, WX6972, WX6974, WX6976, WX6978, WX6980;
wire WX6982, WX6984, WX6986, WX6988, WX6990, WX6992, WX6994, WX6996;
wire WX6998, WX7000, WX7002, WX7004, WX7006, WX7008, WX7010, WX7012;
wire WX7110, WX7112, WX7114, WX7116, WX7118, WX7120, WX7122, WX7124;
wire WX7126, WX7128, WX7130, WX7132, WX7134, WX7136, WX7138, WX7140;
wire WX7142, WX7144, WX7146, WX7148, WX7150, WX7152, WX7154, WX7156;
wire WX7158, WX7160, WX7162, WX7164, WX7166, WX7168, WX7170, WX7172;
wire WX7174, WX7176, WX7178, WX7180, WX7182, WX7184, WX7186, WX7188;
wire WX7190, WX7192, WX7194, WX7196, WX7198, WX7200, WX7202, WX7204;
wire WX7206, WX7208, WX7210, WX7212, WX7214, WX7216, WX7218, WX7220;
wire WX7222, WX7224, WX7226, WX7228, WX7230, WX7232, WX7234, WX7236;
wire WX7238, WX7240, WX7242, WX7244, WX7246, WX7248, WX7250, WX7252;
wire WX7254, WX7256, WX7258, WX7260, WX7262, WX7264, WX7266, WX7268;
wire WX7270, WX7272, WX7274, WX7276, WX7278, WX7280, WX7282, WX7284;
wire WX7286, WX7288, WX7290, WX7292, WX7294, WX7296, WX7298, WX7300;
wire WX7302, WX7304, WX7306, WX7308, WX7310, WX7312, WX7314, WX7316;
wire WX7318, WX7320, WX7322, WX7324, WX7326, WX7328, WX7330, WX7332;
wire WX7334, WX7336, WX7338, WX7340, WX7342, WX7344, WX7346, WX7348;
wire WX7350, WX7352, WX7354, WX7356, WX7358, WX7360, WX7362, WX7364;
wire WX8243, WX8245, WX8247, WX8249, WX8251, WX8253, WX8255, WX8257;
wire WX8259, WX8261, WX8263, WX8265, WX8267, WX8269, WX8271, WX8273;
wire WX8275, WX8277, WX8279, WX8281, WX8283, WX8285, WX8287, WX8289;
wire WX8291, WX8293, WX8295, WX8297, WX8299, WX8301, WX8303, WX8305;
wire WX8403, WX8405, WX8407, WX8409, WX8411, WX8413, WX8415, WX8417;
wire WX8419, WX8421, WX8423, WX8425, WX8427, WX8429, WX8431, WX8433;
wire WX8435, WX8437, WX8439, WX8441, WX8443, WX8445, WX8447, WX8449;
wire WX8451, WX8453, WX8455, WX8457, WX8459, WX8461, WX8463, WX8465;
wire WX8467, WX8469, WX8471, WX8473, WX8475, WX8477, WX8479, WX8481;
wire WX8483, WX8485, WX8487, WX8489, WX8491, WX8493, WX8495, WX8497;
wire WX8499, WX8501, WX8503, WX8505, WX8507, WX8509, WX8511, WX8513;
wire WX8515, WX8517, WX8519, WX8521, WX8523, WX8525, WX8527, WX8529;
wire WX8531, WX8533, WX8535, WX8537, WX8539, WX8541, WX8543, WX8545;
wire WX8547, WX8549, WX8551, WX8553, WX8555, WX8557, WX8559, WX8561;
wire WX8563, WX8565, WX8567, WX8569, WX8571, WX8573, WX8575, WX8577;
wire WX8579, WX8581, WX8583, WX8585, WX8587, WX8589, WX8591, WX8593;
wire WX8595, WX8597, WX8599, WX8601, WX8603, WX8605, WX8607, WX8609;
wire WX8611, WX8613, WX8615, WX8617, WX8619, WX8621, WX8623, WX8625;
wire WX8627, WX8629, WX8631, WX8633, WX8635, WX8637, WX8639, WX8641;
wire WX8643, WX8645, WX8647, WX8649, WX8651, WX8653, WX8655, WX8657;
wire WX9536, WX9538, WX9540, WX9542, WX9544, WX9546, WX9548, WX9550;
wire WX9552, WX9554, WX9556, WX9558, WX9560, WX9562, WX9564, WX9566;
wire WX9568, WX9570, WX9572, WX9574, WX9576, WX9578, WX9580, WX9582;
wire WX9584, WX9586, WX9588, WX9590, WX9592, WX9594, WX9596, WX9598;
wire WX9696, WX9698, WX9700, WX9702, WX9704, WX9706, WX9708, WX9710;
wire WX9712, WX9714, WX9716, WX9718, WX9720, WX9722, WX9724, WX9726;
wire WX9728, WX9730, WX9732, WX9734, WX9736, WX9738, WX9740, WX9742;
wire WX9744, WX9746, WX9748, WX9750, WX9752, WX9754, WX9756, WX9758;
wire WX9760, WX9762, WX9764, WX9766, WX9768, WX9770, WX9772, WX9774;
wire WX9776, WX9778, WX9780, WX9782, WX9784, WX9786, WX9788, WX9790;
wire WX9792, WX9794, WX9796, WX9798, WX9800, WX9802, WX9804, WX9806;
wire WX9808, WX9810, WX9812, WX9814, WX9816, WX9818, WX9820, WX9822;
wire WX9824, WX9826, WX9828, WX9830, WX9832, WX9834, WX9836, WX9838;
wire WX9840, WX9842, WX9844, WX9846, WX9848, WX9850, WX9852, WX9854;
wire WX9856, WX9858, WX9860, WX9862, WX9864, WX9866, WX9868, WX9870;
wire WX9872, WX9874, WX9876, WX9878, WX9880, WX9882, WX9884, WX9886;
wire WX9888, WX9890, WX9892, WX9894, WX9896, WX9898, WX9900, WX9902;
wire WX9904, WX9906, WX9908, WX9910, WX9912, WX9914, WX9916, WX9918;
wire WX9920, WX9922, WX9924, WX9926, WX9928, WX9930, WX9932, WX9934;
wire WX9936, WX9938, WX9940, WX9942, WX9944, WX9946, WX9948, WX9950;
wire WX10829, WX10831, WX10833, WX10835, WX10837, WX10839, WX10841,WX10843;
wire WX10845, WX10847, WX10849, WX10851, WX10853, WX10855, WX10857,WX10859;
wire WX10861, WX10863, WX10865, WX10867, WX10869, WX10871, WX10873,WX10875;
wire WX10877, WX10879, WX10881, WX10883, WX10885, WX10887, WX10889,WX10891;
wire WX10989, WX10991, WX10993, WX10995, WX10997, WX10999, WX11001,WX11003;
wire WX11005, WX11007, WX11009, WX11011, WX11013, WX11015, WX11017,WX11019;
wire WX11021, WX11023, WX11025, WX11027, WX11029, WX11031, WX11033,WX11035;
wire WX11037, WX11039, WX11041, WX11043, WX11045, WX11047, WX11049,WX11051;
wire WX11053, WX11055, WX11057, WX11059, WX11061, WX11063, WX11065,WX11067;
wire WX11069, WX11071, WX11073, WX11075, WX11077, WX11079, WX11081,WX11083;
wire WX11085, WX11087, WX11089, WX11091, WX11093, WX11095, WX11097,WX11099;
wire WX11101, WX11103, WX11105, WX11107, WX11109, WX11111, WX11113,WX11115;
wire WX11117, WX11119, WX11121, WX11123, WX11125, WX11127, WX11129,WX11131;
wire WX11133, WX11135, WX11137, WX11139, WX11141, WX11143, WX11145,WX11147;
wire WX11149, WX11151, WX11153, WX11155, WX11157, WX11159, WX11161,WX11163;
wire WX11165, WX11167, WX11169, WX11171, WX11173, WX11175, WX11177,WX11179;
wire WX11181, WX11183, WX11185, WX11187, WX11189, WX11191, WX11193,WX11195;
wire WX11197, WX11199, WX11201, WX11203, WX11205, WX11207, WX11209,WX11211;
wire WX11213, WX11215, WX11217, WX11219, WX11221, WX11223, WX11225,WX11227;
wire WX11229, WX11231, WX11233, WX11235, WX11237, WX11239, WX11241,WX11243;
wire _2077_, _2078_, _2079_, _2080_, _2081_, _2082_, _2083_, _2084_;
wire _2085_, _2086_, _2087_, _2088_, _2089_, _2090_, _2091_, _2092_;
wire _2093_, _2094_, _2095_, _2096_, _2097_, _2098_, _2099_, _2100_;
wire _2101_, _2102_, _2103_, _2104_, _2105_, _2106_, _2107_, _2108_;
wire _2109_, _2110_, _2111_, _2112_, _2113_, _2114_, _2115_, _2116_;
wire _2117_, _2118_, _2119_, _2120_, _2121_, _2122_, _2123_, _2124_;
wire _2125_, _2126_, _2127_, _2128_, _2129_, _2130_, _2131_, _2132_;
wire _2133_, _2134_, _2135_, _2136_, _2137_, _2138_, _2139_, _2140_;
wire _2141_, _2142_, _2143_, _2144_, _2145_, _2146_, _2147_, _2148_;
wire _2149_, _2150_, _2151_, _2152_, _2153_, _2154_, _2155_, _2156_;
wire _2157_, _2158_, _2159_, _2160_, _2161_, _2162_, _2163_, _2164_;
wire _2165_, _2166_, _2167_, _2168_, _2169_, _2170_, _2171_, _2172_;
wire _2173_, _2174_, _2175_, _2176_, _2177_, _2178_, _2179_, _2180_;
wire _2181_, _2182_, _2183_, _2184_, _2185_, _2186_, _2187_, _2188_;
wire _2189_, _2190_, _2191_, _2192_, _2193_, _2194_, _2195_, _2196_;
wire _2197_, _2198_, _2199_, _2200_, _2201_, _2202_, _2203_, _2204_;
wire _2205_, _2206_, _2207_, _2208_, _2209_, _2210_, _2211_, _2212_;
wire _2213_, _2214_, _2215_, _2216_, _2217_, _2218_, _2219_, _2220_;
wire _2221_, _2222_, _2223_, _2224_, _2225_, _2226_, _2227_, _2228_;
wire _2229_, _2230_, _2231_, _2232_, _2233_, _2234_, _2235_, _2236_;
wire _2237_, _2238_, _2239_, _2240_, _2241_, _2242_, _2243_, _2244_;
wire _2245_, _2246_, _2247_, _2248_, _2249_, _2250_, _2251_, _2252_;
wire _2253_, _2254_, _2255_, _2256_, _2257_, _2258_, _2259_, _2260_;
wire _2261_, _2262_, _2263_, _2264_, _2265_, _2266_, _2267_, _2268_;
wire _2269_, _2270_, _2271_, _2272_, _2273_, _2274_, _2275_, _2276_;
wire _2277_, _2278_, _2279_, _2280_, _2281_, _2282_, _2283_, _2284_;
wire _2285_, _2286_, _2287_, _2288_, _2289_, _2290_, _2291_, _2292_;
wire _2293_, _2294_, _2295_, _2296_, _2297_, _2298_, _2299_, _2300_;
wire _2301_, _2302_, _2303_, _2304_, _2305_, _2306_, _2307_, _2308_;
wire _2309_, _2310_, _2311_, _2312_, _2313_, _2314_, _2315_, _2316_;
wire _2317_, _2318_, _2319_, _2320_, _2321_, _2322_, _2323_, _2324_;
wire _2325_, _2326_, _2327_, _2328_, _2329_, _2330_, _2331_, _2332_;
wire _2333_, _2334_, _2335_, _2336_, _2337_, _2338_, _2339_, _2340_;
wire _2341_, _2342_, _2343_, _2344_, _2345_, _2346_, _2347_, _2348_;
wire _2349_, _2350_, _2351_, _2352_, _2353_, _2354_, _2355_, _2356_;
wire _2357_, _2358_, _2359_, _2360_, _2361_, _2362_, _2363_, _2364_;
wire n_0, n_2, n_3, n_4, n_5, n_12, n_14, n_16;
wire n_18, n_19, n_20, n_21, n_24, n_27, n_28, n_32;
wire n_33, n_35, n_36, n_38, n_40, n_41, n_43, n_44;
wire n_46, n_48, n_49, n_51, n_52, n_56, n_58, n_63;
wire n_65, n_67, n_68, n_69, n_70, n_71, n_73, n_79;
wire n_81, n_83, n_85, n_87, n_89, n_95, n_96, n_98;
wire n_100, n_101, n_104, n_105, n_106, n_108, n_109, n_111;
wire n_112, n_113, n_117, n_118, n_119, n_120, n_124, n_126;
wire n_127, n_129, n_130, n_131, n_133, n_135, n_136, n_137;
wire n_139, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
wire n_180, n_181, n_183, n_184, n_185, n_186, n_187, n_188;
wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_197;
wire n_198, n_199, n_200, n_201, n_204, n_205, n_206, n_207;
wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_219;
wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
wire n_233, n_235, n_236, n_241, n_244, n_247, n_252, n_254;
wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_264;
wire n_266, n_268, n_271, n_273, n_276, n_278, n_280, n_282;
wire n_283, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
wire n_292, n_293, n_294, n_295, n_296, n_297, n_298, n_299;
wire n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307;
wire n_308, n_310, n_311, n_312, n_313, n_314, n_315, n_316;
wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
wire n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332;
wire n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340;
wire n_341, n_342, n_343, n_344, n_345, n_346, n_347, n_348;
wire n_349, n_350, n_351, n_352, n_353, n_354, n_356, n_357;
wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
wire n_398, n_399, n_401, n_402, n_403, n_404, n_405, n_406;
wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
wire n_415, n_416, n_417, n_418, n_419, n_420, n_422, n_423;
wire n_424, n_426, n_427, n_428, n_429, n_431, n_433, n_434;
wire n_436, n_438, n_440, n_442, n_443, n_447, n_448, n_450;
wire n_451, n_453, n_454, n_456, n_457, n_458, n_460, n_461;
wire n_462, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
wire n_471, n_472, n_473, n_474, n_476, n_478, n_479, n_480;
wire n_482, n_484, n_486, n_488, n_489, n_490, n_491, n_492;
wire n_495, n_496, n_497, n_499, n_500, n_501, n_502, n_503;
wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_514;
wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
wire n_523, n_524, n_525, n_526, n_527, n_529, n_530, n_531;
wire n_532, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
wire n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581;
wire n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589;
wire n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597;
wire n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605;
wire n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613;
wire n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621;
wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
wire n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677;
wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685;
wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
wire n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702;
wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
wire n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718;
wire n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726;
wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
wire n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742;
wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
wire n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
wire n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790;
wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814;
wire n_815, n_816, n_817, n_823, n_830, n_831, n_836, n_842;
wire n_846, n_847, n_848, n_849, n_850, n_852, n_853, n_857;
wire n_858, n_860, n_866, n_867, n_868, n_869, n_873, n_874;
wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
wire n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898;
wire n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906;
wire n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
wire n_915, n_916, n_918, n_919, n_920, n_921, n_922, n_923;
wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931;
wire n_932, n_933, n_935, n_937, n_938, n_939, n_940, n_941;
wire n_942, n_943, n_944, n_945, n_947, n_948, n_949, n_950;
wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
wire n_959, n_960, n_962, n_963, n_964, n_965, n_966, n_967;
wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
wire n_977, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
wire n_986, n_987, n_988, n_990, n_991, n_992, n_993, n_994;
wire n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002;
wire n_1003, n_1004, n_1005, n_1006, n_1007, n_1009, n_1011, n_1012;
wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020;
wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044;
wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052;
wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060;
wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100;
wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132;
wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140;
wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148;
wire n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156;
wire n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164;
wire n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172;
wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180;
wire n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228;
wire n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
wire n_1237, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
wire n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261;
wire n_1262, n_1263, n_1264, n_1265, n_1267, n_1268, n_1272, n_1275;
wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
wire n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291;
wire n_1294, n_1297, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
wire n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318;
wire n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326;
wire n_1327, n_1328, n_1329, n_1330, n_1332, n_1333, n_1334, n_1335;
wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1344;
wire n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
wire n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360;
wire n_1362, n_1364, n_1365, n_1366, n_1367, n_1369, n_1370, n_1371;
wire n_1372, n_1373, n_1374, n_1375, n_1377, n_1378, n_1379, n_1380;
wire n_1381, n_1382, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
wire n_1391, n_1393, n_1395, n_1396, n_1398, n_1399, n_1400, n_1402;
wire n_1403, n_1404, n_1405, n_1407, n_1409, n_1410, n_1411, n_1412;
wire n_1413, n_1414, n_1415, n_1417, n_1418, n_1419, n_1420, n_1421;
wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
wire n_1430, n_1431, n_1432, n_1433, n_1435, n_1436, n_1437, n_1438;
wire n_1440, n_1441, n_1442, n_1443, n_1444, n_1446, n_1447, n_1448;
wire n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1456, n_1458;
wire n_1459, n_1460, n_1461, n_1462, n_1464, n_1465, n_1470, n_1471;
wire n_1472, n_1473, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481;
wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
wire n_1498, n_1499, n_1500, n_1502, n_1503, n_1504, n_1506, n_1507;
wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
wire n_1516, n_1517, n_1518, n_1519, n_1521, n_1522, n_1523, n_1524;
wire n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1533;
wire n_1534, n_1535, n_1536, n_1537, n_1539, n_1540, n_1541, n_1542;
wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1550, n_1551, n_1552;
wire n_1553, n_1554, n_1555, n_1557, n_1558, n_1559, n_1560, n_1561;
wire n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1570, n_1571;
wire n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1579, n_1580;
wire n_1581, n_1582, n_1583, n_1584, n_1585, n_1587, n_1588, n_1590;
wire n_1591, n_1592, n_1593, n_1594, n_1595, n_1597, n_1598, n_1599;
wire n_1600, n_1601, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608;
wire n_1609, n_1611, n_1612, n_1613, n_1614, n_1615, n_1617, n_1618;
wire n_1619, n_1620, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627;
wire n_1628, n_1629, n_1631, n_1632, n_1633, n_1635, n_1636, n_1637;
wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1644, n_1645, n_1646;
wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1654, n_1655;
wire n_1656, n_1658, n_1659, n_1660, n_1661, n_1662, n_1664, n_1665;
wire n_1666, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1675;
wire n_1676, n_1677, n_1678, n_1679, n_1681, n_1682, n_1684, n_1685;
wire n_1687, n_1688, n_1690, n_1691, n_1693, n_1694, n_1696, n_1697;
wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1706, n_1707, n_1708;
wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
wire n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732;
wire n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740;
wire n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748;
wire n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756;
wire n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764;
wire n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772;
wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
wire n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796;
wire n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804;
wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
wire n_1837, n_1838, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845;
wire n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853;
wire n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861;
wire n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869;
wire n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877;
wire n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885;
wire n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893;
wire n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901;
wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909;
wire n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917;
wire n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925;
wire n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933;
wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
wire n_1950, n_1951, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958;
wire n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966;
wire n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974;
wire n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982;
wire n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990;
wire n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998;
wire n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
wire n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014;
wire n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022;
wire n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030;
wire n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038;
wire n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046;
wire n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054;
wire n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062;
wire n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070;
wire n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078;
wire n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086;
wire n_2087, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
wire n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103;
wire n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111;
wire n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
wire n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127;
wire n_2128, n_2129, n_2130, n_2132, n_2133, n_2134, n_2135, n_2136;
wire n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144;
wire n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152;
wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176;
wire n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2185;
wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
wire n_2194, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202;
wire n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210;
wire n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218;
wire n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226;
wire n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234;
wire n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242;
wire n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250;
wire n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258;
wire n_2259, n_2260, n_2261, n_2262, n_2264, n_2266, n_2267, n_2268;
wire n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276;
wire n_2277, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285;
wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
wire n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302;
wire n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310;
wire n_2311, n_2312, n_2313, n_2315, n_2316, n_2317, n_2318, n_2320;
wire n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2328, n_2329;
wire n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337;
wire n_2338, n_2339, n_2340, n_2341, n_2343, n_2344, n_2345, n_2346;
wire n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2355;
wire n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363;
wire n_2364, n_2365, n_2366, n_2368, n_2369, n_2370, n_2371, n_2372;
wire n_2373, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2382;
wire n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390;
wire n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398;
wire n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406;
wire n_2408, n_2409, n_2412, n_2419, n_2420, n_2421, n_2422, n_2423;
wire n_2424, n_2425, n_2428, n_2431, n_2433, n_2434, n_2437, n_2438;
wire n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446;
wire n_2447, n_2448, n_2452, n_2453, n_2454, n_2457, n_2458, n_2459;
wire n_2462, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471;
wire n_2472, n_2473, n_2475, n_2476, n_2477, n_2480, n_2481, n_2484;
wire n_2487, n_2488, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498;
wire n_2499, n_2500, n_2503, n_2504, n_2505, n_2508, n_2511, n_2512;
wire n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520;
wire n_2521, n_2522, n_2523, n_2524, n_2525, n_2527, n_2528, n_2529;
wire n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537;
wire n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545;
wire n_2546, n_2547, n_2548, n_2551, n_2552, n_2553, n_2554, n_2555;
wire n_2556, n_2557, n_2558, n_2559, n_2562, n_2563, n_2564, n_2565;
wire n_2566, n_2567, n_2568, n_2570, n_2571, n_2572, n_2573, n_2574;
wire n_2575, n_2576, n_2577, n_2579, n_2581, n_2582, n_2583, n_2584;
wire n_2585, n_2587, n_2588, n_2589, n_2590, n_2591, n_2593, n_2594;
wire n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602;
wire n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610;
wire n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618;
wire n_2619, n_2620, n_2621, n_2622, n_2624, n_2625, n_2626, n_2627;
wire n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635;
wire n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643;
wire n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
wire n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659;
wire n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667;
wire n_2668, n_2669, n_2670, n_2671, n_2673, n_2675, n_2676, n_2677;
wire n_2678, n_2680, n_2681, n_2682, n_2684, n_2685, n_2686, n_2687;
wire n_2689, n_2690, n_2691, n_2692, n_2694, n_2695, n_2696, n_2697;
wire n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705;
wire n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713;
wire n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721;
wire n_2722, n_2724, n_2725, n_2726, n_2728, n_2729, n_2730, n_2731;
wire n_2732, n_2733, n_2734, n_2736, n_2737, n_2738, n_2739, n_2741;
wire n_2742, n_2743, n_2744, n_2745, n_2746, n_2749, n_2750, n_2752;
wire n_2754, n_2755, n_2756, n_2757, n_2759, n_2760, n_2761, n_2762;
wire n_2763, n_2765, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772;
wire n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2780, n_2782;
wire n_2783, n_2784, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791;
wire n_2792, n_2793, n_2794, n_2795, n_2797, n_2798, n_2799, n_2800;
wire n_2801, n_2803, n_2805, n_2806, n_2807, n_2809, n_2810, n_2811;
wire n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2820;
wire n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829;
wire n_2830, n_2831, n_2833, n_2835, n_2836, n_2837, n_2838, n_2839;
wire n_2840, n_2843, n_2844, n_2846, n_2847, n_2848, n_2849, n_2850;
wire n_2851, n_2852, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859;
wire n_2860, n_2861, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868;
wire n_2870, n_2872, n_2873, n_2875, n_2876, n_2878, n_2879, n_2881;
wire n_2882, n_2883, n_2884, n_2885, n_2887, n_2888, n_2889, n_2892;
wire n_2893, n_2894, n_2897, n_2898, n_2900, n_2902, n_2903, n_2905;
wire n_2906, n_2907, n_2908, n_2909, n_2911, n_2912, n_2914, n_2916;
wire n_2917, n_2920, n_2921, n_2922, n_2924, n_2925, n_2926, n_2927;
wire n_2928, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936;
wire n_2937, n_2938, n_2939, n_2940, n_2941, n_2943, n_2944, n_2945;
wire n_2946, n_2947, n_2948, n_2949, n_2950, n_2952, n_2953, n_2954;
wire n_2955, n_2957, n_2958, n_2960, n_2961, n_2963, n_2965, n_2966;
wire n_2967, n_2968, n_2969, n_2971, n_2972, n_2974, n_2975, n_2976;
wire n_2978, n_2979, n_2981, n_2982, n_2984, n_2985, n_2986, n_2987;
wire n_2988, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996;
wire n_2997, n_2998, n_2999, n_3000, n_3001, n_3003, n_3004, n_3005;
wire n_3007, n_3009, n_3011, n_3012, n_3014, n_3015, n_3017, n_3018;
wire n_3020, n_3021, n_3022, n_3023, n_3024, n_3026, n_3027, n_3028;
wire n_3029, n_3030, n_3031, n_3032, n_3034, n_3037, n_3038, n_3039;
wire n_3040, n_3041, n_3043, n_3044, n_3045, n_3047, n_3048, n_3049;
wire n_3051, n_3052, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059;
wire n_3061, n_3062, n_3064, n_3065, n_3066, n_3068, n_3069, n_3071;
wire n_3072, n_3074, n_3075, n_3076, n_3077, n_3080, n_3081, n_3083;
wire n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3092, n_3093;
wire n_3095, n_3096, n_3098, n_3099, n_3101, n_3102, n_3103, n_3104;
wire n_3105, n_3106, n_3107, n_3108, n_3110, n_3111, n_3113, n_3114;
wire n_3115, n_3116, n_3117, n_3118, n_3120, n_3121, n_3123, n_3125;
wire n_3126, n_3127, n_3128, n_3131, n_3134, n_3135, n_3136, n_3137;
wire n_3138, n_3139, n_3140, n_3141, n_3142, n_3145, n_3147, n_3149;
wire n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158;
wire n_3162, n_3163, n_3167, n_3168, n_3169, n_3173, n_3177, n_3178;
wire n_3179, n_3180, n_3181, n_3183, n_3186, n_3187, n_3188, n_3189;
wire n_3190, n_3191, n_3192, n_3194, n_3195, n_3197, n_3198, n_3199;
wire n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3207, n_3208;
wire n_3210, n_3211, n_3212, n_3213, n_3215, n_3216, n_3217, n_3218;
wire n_3219, n_3221, n_3222, n_3223, n_3224, n_3225, n_3227, n_3230;
wire n_3231, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239;
wire n_3240, n_3241, n_3242, n_3243, n_3244, n_3249, n_3250, n_3253;
wire n_3254, n_3255, n_3256, n_3257, n_3260, n_3261, n_3262, n_3263;
wire n_3264, n_3265, n_3268, n_3269, n_3272, n_3273, n_3276, n_3278;
wire n_3280, n_3281, n_3282, n_3285, n_3286, n_3287, n_3290, n_3291;
wire n_3292, n_3293, n_3296, n_3297, n_3299, n_3300, n_3301, n_3302;
wire n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310;
wire n_3311, n_3312, n_3313, n_3314, n_3315, n_3318, n_3319, n_3320;
wire n_3321, n_3322, n_3323, n_3324, n_3327, n_3330, n_3333, n_3334;
wire n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342;
wire n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3352;
wire n_3353, n_3356, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364;
wire n_3365, n_3366, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374;
wire n_3375, n_3376, n_3377, n_3378, n_3379, n_3382, n_3383, n_3384;
wire n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3393, n_3394;
wire n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402;
wire n_3403, n_3404, n_3405, n_3408, n_3409, n_3410, n_3411, n_3414;
wire n_3421, n_3426, n_3428, n_3431, n_3433, n_3434, n_3435, n_3436;
wire n_3437, n_3439, n_3443, n_3447, n_3449, n_3450, n_3451, n_3452;
wire n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460;
wire n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468;
wire n_3469, n_3470, n_3471, n_3472, n_3474, n_3475, n_3476, n_3477;
wire n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485;
wire n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493;
wire n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501;
wire n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509;
wire n_3510, n_3511, n_3512, n_3513, n_3514, n_3516, n_3517, n_3518;
wire n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526;
wire n_3527, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535;
wire n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543;
wire n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551;
wire n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559;
wire n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567;
wire n_3568, n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575;
wire n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, n_3582, n_3583;
wire n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3591, n_3592;
wire n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600;
wire n_3601, n_3604, n_3605, n_3606, n_3609, n_3612, n_3614, n_3616;
wire n_3620, n_3621, n_3622, n_3626, n_3628, n_3632, n_3633, n_3637;
wire n_3639, n_3642, n_3643, n_3647, n_3648, n_3650, n_3652, n_3653;
wire n_3658, n_3663, n_3664, n_3666, n_3669, n_3670, n_3676, n_3678;
wire n_3679, n_3681, n_3682, n_3684, n_3685, n_3686, n_3688, n_3689;
wire n_3690, n_3691, n_3692, n_3694, n_3695, n_3696, n_3698, n_3699;
wire n_3701, n_3702, n_3703, n_3707, n_3708, n_3709, n_3710, n_3711;
wire n_3712, n_3713, n_3714, n_3715, n_3716, n_3718, n_3719, n_3722;
wire n_3724, n_3726, n_3729, n_3731, n_3732, n_3733, n_3734, n_3735;
wire n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3744;
wire n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753;
wire n_3755, n_3757, n_3758, n_3759, n_3761, n_3762, n_3764, n_3765;
wire n_3766, n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773;
wire n_3774, n_3775, n_3776, n_3778, n_3781, n_3782, n_3783, n_3785;
wire n_3786, n_3787, n_3790, n_3792, n_3793, n_3795, n_3796, n_3798;
wire n_3799, n_3800, n_3801, n_3802, n_3804, n_3805, n_3806, n_3807;
wire n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3815, n_3816;
wire n_3817, n_3818, n_3819, n_3821, n_3822, n_3824, n_3826, n_3827;
wire n_3828, n_3829, n_3830, n_3831, n_3833, n_3834, n_3835, n_3836;
wire n_3837, n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845;
wire n_3846, n_3848, n_3850, n_3853, n_3854, n_3855, n_3856, n_3857;
wire n_3859, n_3860, n_3863, n_3864, n_3865, n_3868, n_3870, n_3871;
wire n_3872, n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880;
wire n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888;
wire n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3898;
wire n_3900, n_3901, n_3903, n_3906, n_3908, n_3910, n_3911, n_3912;
wire n_3913, n_3914, n_3915, n_3916, n_3917, n_3919, n_3920, n_3921;
wire n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3930, n_3932;
wire n_3933, n_3934, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941;
wire n_3942, n_3943, n_3944, n_3945, n_3947, n_3948, n_3951, n_3952;
wire n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960;
wire n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968;
wire n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976;
wire n_3977, n_3979, n_3980, n_3981, n_3982, n_3984, n_3985, n_3987;
wire n_3988, n_3990, n_3991, n_3992, n_3993, n_3994, n_3995, n_3996;
wire n_3997, n_3998, n_3999, n_4000, n_4001, n_4002, n_4005, n_4006;
wire n_4007, n_4009, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016;
wire n_4017, n_4018, n_4019, n_4021, n_4023, n_4025, n_4026, n_4027;
wire n_4029, n_4031, n_4033, n_4035, n_4037, n_4038, n_4039, n_4040;
wire n_4041, n_4043, n_4044, n_4045, n_4047, n_4049, n_4050, n_4051;
wire n_4052, n_4053, n_4055, n_4057, n_4058, n_4060, n_4061, n_4062;
wire n_4064, n_4066, n_4068, n_4069, n_4070, n_4071, n_4072, n_4075;
wire n_4076, n_4077, n_4078, n_4079, n_4080, n_4082, n_4083, n_4084;
wire n_4086, n_4087, n_4088, n_4090, n_4092, n_4093, n_4094, n_4095;
wire n_4096, n_4099, n_4100, n_4101, n_4103, n_4104, n_4105, n_4106;
wire n_4107, n_4108, n_4109, n_4111, n_4112, n_4113, n_4114, n_4115;
wire n_4116, n_4117, n_4119, n_4121, n_4122, n_4123, n_4124, n_4125;
wire n_4126, n_4127, n_4128, n_4129, n_4130, n_4131, n_4132, n_4133;
wire n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4140, n_4141;
wire n_4142, n_4143, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149;
wire n_4150, n_4151, n_4152, n_4153, n_4154, n_4155, n_4156, n_4157;
wire n_4158, n_4159, n_4160, n_4161, n_4162, n_4163, n_4164, n_4165;
wire n_4166, n_4167, n_4168, n_4169, n_4170, n_4171, n_4172, n_4173;
wire n_4174, n_4175, n_4176, n_4177, n_4178, n_4179, n_4180, n_4181;
wire n_4182, n_4183, n_4184, n_4185, n_4186, n_4187, n_4188, n_4190;
wire n_4191, n_4192, n_4193, n_4194, n_4195, n_4197, n_4198, n_4199;
wire n_4201, n_4203, n_4204, n_4205, n_4207, n_4208, n_4209, n_4210;
wire n_4211, n_4213, n_4215, n_4218, n_4219, n_4220, n_4221, n_4222;
wire n_4223, n_4224, n_4225, n_4227, n_4228, n_4229, n_4230, n_4231;
wire n_4232, n_4233, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240;
wire n_4241, n_4243, n_4244, n_4245, n_4247, n_4248, n_4249, n_4250;
wire n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257, n_4258;
wire n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265, n_4266;
wire n_4267, n_4269, n_4271, n_4272, n_4273, n_4274, n_4275, n_4276;
wire n_4277, n_4279, n_4280, n_4281, n_4282, n_4283, n_4285, n_4286;
wire n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293, n_4294;
wire n_4295, n_4297, n_4298, n_4299, n_4301, n_4302, n_4303, n_4304;
wire n_4305, n_4307, n_4308, n_4309, n_4310, n_4311, n_4312, n_4313;
wire n_4314, n_4315, n_4316, n_4317, n_4318, n_4319, n_4320, n_4322;
wire n_4323, n_4324, n_4325, n_4326, n_4327, n_4328, n_4329, n_4330;
wire n_4331, n_4332, n_4333, n_4334, n_4335, n_4336, n_4337, n_4338;
wire n_4339, n_4340, n_4341, n_4342, n_4343, n_4345, n_4346, n_4347;
wire n_4348, n_4349, n_4350, n_4351, n_4353, n_4354, n_4355, n_4356;
wire n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364;
wire n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372;
wire n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380;
wire n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388;
wire n_4389, n_4390, n_4392, n_4394, n_4395, n_4396, n_4398, n_4399;
wire n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4408;
wire n_4409, n_4410, n_4411, n_4412, n_4413, n_4414, n_4415, n_4416;
wire n_4417, n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424;
wire n_4425, n_4426, n_4427, n_4428, n_4429, n_4430, n_4431, n_4432;
wire n_4433, n_4434, n_4435, n_4436, n_4437, n_4438, n_4439, n_4440;
wire n_4441, n_4442, n_4444, n_4446, n_4447, n_4448, n_4449, n_4450;
wire n_4451, n_4452, n_4454, n_4455, n_4456, n_4457, n_4458, n_4459;
wire n_4460, n_4461, n_4462, n_4463, n_4464, n_4465, n_4466, n_4467;
wire n_4468, n_4469, n_4471, n_4472, n_4473, n_4474, n_4476, n_4477;
wire n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485;
wire n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493;
wire n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501;
wire n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509;
wire n_4510, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517, n_4518;
wire n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526;
wire n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534;
wire n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542;
wire n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549, n_4551;
wire n_4552, n_4553, n_4554, n_4555, n_4556, n_4557, n_4558, n_4559;
wire n_4560, n_4562, n_4563, n_4564, n_4565, n_4566, n_4567, n_4568;
wire n_4569, n_4570, n_4571, n_4572, n_4573, n_4574, n_4575, n_4577;
wire n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584, n_4586;
wire n_4587, n_4588, n_4589, n_4590, n_4591, n_4592, n_4593, n_4594;
wire n_4595, n_4596, n_4597, n_4598, n_4599, n_4600, n_4601, n_4602;
wire n_4603, n_4604, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610;
wire n_4611, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618, n_4620;
wire n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629;
wire n_4630, n_4631, n_4633, n_4634, n_4636, n_4638, n_4639, n_4640;
wire n_4641, n_4642, n_4643, n_4644, n_4645, n_4646, n_4647, n_4648;
wire n_4649, n_4650, n_4651, n_4652, n_4653, n_4654, n_4655, n_4656;
wire n_4657, n_4658, n_4659, n_4660, n_4661, n_4662, n_4665, n_4667;
wire n_4669, n_4670, n_4671, n_4672, n_4673, n_4674, n_4676, n_4677;
wire n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685;
wire n_4686, n_4687, n_4688, n_4689, n_4690, n_4692, n_4693, n_4695;
wire n_4696, n_4697, n_4698, n_4702, n_4704, n_4706, n_4711, n_4714;
wire n_4715, n_4716, n_4717, n_4719, n_4720, n_4721, n_4722, n_4723;
wire n_4725, n_4727, n_4728, n_4729, n_4730, n_4731, n_4733, n_4734;
wire n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742;
wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
wire n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758;
wire n_4759, n_4760, n_4761, n_4762, n_4765, n_4766, n_4768, n_4769;
wire n_4770, n_4771, n_4772, n_4773, n_4774, n_4775, n_4777, n_4778;
wire n_4779, n_4780, n_4781, n_4783, n_4784, n_4785, n_4786, n_4788;
wire n_4790, n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797;
wire n_4798, n_4799, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806;
wire n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814;
wire n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822;
wire n_4823, n_4824, n_4825, n_4827, n_4828, n_4829, n_4830, n_4832;
wire n_4833, n_4834, n_4835, n_4837, n_4838, n_4839, n_4840, n_4841;
wire n_4842, n_4844, n_4845, n_4848, n_4851, n_4852, n_4853, n_4854;
wire n_4857, n_4858, n_4859, n_4860, n_4861, n_4863, n_4864, n_4865;
wire n_4866, n_4867, n_4868, n_4869, n_4870, n_4871, n_4873, n_4874;
wire n_4875, n_4876, n_4877, n_4879, n_4880, n_4881, n_4882, n_4883;
wire n_4884, n_4887, n_4888, n_4890, n_4891, n_4893, n_4899, n_4902;
wire n_4903, n_4904, n_4905, n_4906, n_4907, n_4908, n_4909, n_4911;
wire n_4912, n_4913, n_4915, n_4916, n_4917, n_4918, n_4920, n_4921;
wire n_4922, n_4923, n_4924, n_4925, n_4927, n_4930, n_4934, n_4935;
wire n_4936, n_4938, n_4939, n_4941, n_4942, n_4943, n_4944, n_4945;
wire n_4946, n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953;
wire n_4954, n_4955, n_4956, n_4958, n_4959, n_4960, n_4961, n_4962;
wire n_4963, n_4964, n_4966, n_4968, n_4970, n_4973, n_4974, n_4976;
wire n_4978, n_4979, n_4980, n_4984, n_4985, n_4986, n_4988, n_4991;
wire n_4992, n_4994, n_4995, n_4996, n_4997, n_4998, n_4999, n_5001;
wire n_5003, n_5004, n_5005, n_5007, n_5009, n_5010, n_5011, n_5012;
wire n_5016, n_5017, n_5020, n_5022, n_5024, n_5025, n_5027, n_5028;
wire n_5030, n_5034, n_5035, n_5036, n_5037, n_5038, n_5039, n_5040;
wire n_5041, n_5042, n_5043, n_5045, n_5046, n_5047, n_5050, n_5052;
wire n_5053, n_5054, n_5055, n_5056, n_5059, n_5060, n_5062, n_5063;
wire n_5064, n_5065, n_5066, n_5067, n_5069, n_5071, n_5072, n_5073;
wire n_5074, n_5075, n_5076, n_5078, n_5079, n_5080, n_5081, n_5082;
wire n_5083, n_5084, n_5085, n_5086, n_5087, n_5088, n_5089, n_5090;
wire n_5092, n_5095, n_5097, n_5100, n_5102, n_5104, n_5105, n_5106;
wire n_5107, n_5109, n_5110, n_5111, n_5112, n_5113, n_5115, n_5116;
wire n_5117, n_5118, n_5119, n_5121, n_5122, n_5123, n_5126, n_5127;
wire n_5128, n_5129, n_5132, n_5133, n_5135, n_5136, n_5139, n_5141;
wire n_5143, n_5144, n_5145, n_5146, n_5148, n_5149, n_5150, n_5152;
wire n_5153, n_5154, n_5156, n_5157, n_5158, n_5159, n_5160, n_5161;
wire n_5162, n_5164, n_5165, n_5166, n_5169, n_5171, n_5173, n_5177;
wire n_5179, n_5180, n_5181, n_5182, n_5183, n_5184, n_5185, n_5186;
wire n_5187, n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5196;
wire n_5197, n_5198, n_5199, n_5200, n_5201, n_5203, n_5204, n_5207;
wire n_5208, n_5210, n_5211, n_5212, n_5213, n_5214, n_5217, n_5219;
wire n_5222, n_5224, n_5225, n_5226, n_5227, n_5228, n_5230, n_5232;
wire n_5233, n_5234, n_5235, n_5236, n_5237, n_5238, n_5239, n_5240;
wire n_5241, n_5242, n_5243, n_5245, n_5247, n_5249, n_5250, n_5251;
wire n_5252, n_5253, n_5254, n_5255, n_5256, n_5257, n_5259, n_5261;
wire n_5263, n_5264, n_5265, n_5267, n_5269, n_5271, n_5272, n_5273;
wire n_5274, n_5275, n_5276, n_5278, n_5279, n_5281, n_5282, n_5285;
wire n_5287, n_5288, n_5289, n_5291, n_5293, n_5294, n_5297, n_5300;
wire n_5304, n_5305, n_5307, n_5309, n_5310, n_5311, n_5313, n_5314;
wire n_5316, n_5317, n_5318, n_5319, n_5320, n_5321, n_5323, n_5325;
wire n_5328, n_5330, n_5331, n_5333, n_5334, n_5335, n_5336, n_5338;
wire n_5342, n_5343, n_5345, n_5347, n_5348, n_5350, n_5352, n_5353;
wire n_5354, n_5355, n_5356, n_5358, n_5360, n_5361, n_5362, n_5365;
wire n_5366, n_5367, n_5368, n_5369, n_5370, n_5371, n_5376, n_5377;
wire n_5380, n_5382, n_5384, n_5385, n_5386, n_5388, n_5389, n_5390;
wire n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398, n_5401;
wire n_5403, n_5404, n_5407, n_5409, n_5410, n_5411, n_5413, n_5414;
wire n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5424;
wire n_5425, n_5426, n_5427, n_5429, n_5430, n_5432, n_5434, n_5436;
wire n_5437, n_5438, n_5439, n_5440, n_5442, n_5445, n_5446, n_5448;
wire n_5450, n_5453, n_5454, n_5456, n_5458, n_5459, n_5460, n_5461;
wire n_5462, n_5463, n_5464, n_5465, n_5467, n_5468, n_5469, n_5471;
wire n_5472, n_5473, n_5474, n_5475, n_5477, n_5478, n_5479, n_5480;
wire n_5481, n_5482, n_5483, n_5485, n_5486, n_5488, n_5489, n_5490;
wire n_5491, n_5492, n_5493, n_5494, n_5496, n_5497, n_5499, n_5500;
wire n_5503, n_5505, n_5507, n_5509, n_5511, n_5512, n_5513, n_5514;
wire n_5517, n_5518, n_5519, n_5521, n_5523, n_5525, n_5528, n_5529;
wire n_5530, n_5532, n_5533, n_5534, n_5535, n_5536, n_5537, n_5539;
wire n_5540, n_5541, n_5543, n_5545, n_5546, n_5547, n_5548, n_5549;
wire n_5550, n_5551, n_5553, n_5554, n_5555, n_5556, n_5557, n_5558;
wire n_5560, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
wire n_5569, n_5573, n_5576, n_5577, n_5578, n_5579, n_5580, n_5584;
wire n_5588, n_5591, n_5592, n_5594, n_5595, n_5596, n_5597, n_5598;
wire n_5599, n_5600, n_5601, n_5603, n_5604, n_5605, n_5606, n_5608;
wire n_5609, n_5610, n_5612, n_5616, n_5617, n_5618, n_5619, n_5620;
wire n_5621, n_5622, n_5623, n_5625, n_5627, n_5628, n_5629, n_5630;
wire n_5631, n_5633, n_5634, n_5637, n_5638, n_5641, n_5642, n_5643;
wire n_5644, n_5646, n_5648, n_5649, n_5650, n_5651, n_5652, n_5654;
wire n_5657, n_5658, n_5660, n_5661, n_5662, n_5664, n_5665, n_5666;
wire n_5667, n_5669, n_5670, n_5671, n_5672, n_5674, n_5676, n_5678;
wire n_5682, n_5685, n_5686, n_5687, n_5688, n_5689, n_5690, n_5693;
wire n_5694, n_5695, n_5699, n_5700, n_5701, n_5702, n_5703, n_5705;
wire n_5706, n_5707, n_5708, n_5709, n_5711, n_5712, n_5713, n_5714;
wire n_5716, n_5719, n_5720, n_5721, n_5722, n_5723, n_5724, n_5725;
wire n_5727, n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5735;
wire n_5737, n_5738, n_5742, n_5743, n_5744, n_5745, n_5747, n_5748;
wire n_5749, n_5750, n_5751, n_5752, n_5753, n_5754, n_5755, n_5759;
wire n_5760, n_5763, n_5765, n_5766, n_5767, n_5768, n_5769, n_5770;
wire n_5771, n_5773, n_5774, n_5776, n_5777, n_5781, n_5784, n_5788;
wire n_5789, n_5790, n_5791, n_5792, n_5794, n_5796, n_5798, n_5800;
wire n_5801, n_5802, n_5803, n_5804, n_5806, n_5807, n_5809, n_5811;
wire n_5812, n_5813, n_5814, n_5815, n_5816, n_5818, n_5820, n_5821;
wire n_5822, n_5823, n_5824, n_5825, n_5826, n_5828, n_5830, n_5831;
wire n_5833, n_5834, n_5835, n_5837, n_5838, n_5840, n_5841, n_5842;
wire n_5843, n_5844, n_5845, n_5846, n_5847, n_5848, n_5849, n_5851;
wire n_5853, n_5854, n_5855, n_5856, n_5857, n_5858, n_5860, n_5862;
wire n_5865, n_5866, n_5867, n_5869, n_5871, n_5872, n_5873, n_5876;
wire n_5878, n_5879, n_5880, n_5881, n_5882, n_5883, n_5884, n_5885;
wire n_5886, n_5887, n_5888, n_5889, n_5890, n_5891, n_5892, n_5893;
wire n_5894, n_5896, n_5898, n_5899, n_5901, n_5903, n_5905, n_5907;
wire n_5910, n_5912, n_5914, n_5915, n_5916, n_5917, n_5918, n_5919;
wire n_5921, n_5922, n_5924, n_5925, n_5926, n_5927, n_5928, n_5929;
wire n_5931, n_5933, n_5934, n_5936, n_5937, n_5938, n_5939, n_5940;
wire n_5941, n_5942, n_5944, n_5947, n_5948, n_5949, n_5950, n_5951;
wire n_5952, n_5954, n_5956, n_5959, n_5961, n_5963, n_5964, n_5965;
wire n_5966, n_5967, n_5968, n_5969, n_5970, n_5971, n_5973, n_5974;
wire n_5976, n_5977, n_5978, n_5981, n_5982, n_5983, n_5985, n_5986;
wire n_5987, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993, n_5995;
wire n_5996, n_5998, n_5999, n_6000, n_6001, n_6002, n_6003, n_6004;
wire n_6007, n_6008, n_6010, n_6011, n_6012, n_6013, n_6014, n_6015;
wire n_6017, n_6019, n_6020, n_6021, n_6022, n_6023, n_6024, n_6025;
wire n_6027, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6036;
wire n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6046, n_6047;
wire n_6048, n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6057;
wire n_6058, n_6059, n_6060, n_6061, n_6063, n_6064, n_6066, n_6067;
wire n_6068, n_6069, n_6070, n_6072, n_6074, n_6075, n_6076, n_6078;
wire n_6079, n_6080, n_6081, n_6083, n_6084, n_6085, n_6086, n_6087;
wire n_6088, n_6090, n_6091, n_6092, n_6093, n_6095, n_6096, n_6097;
wire n_6099, n_6100, n_6102, n_6103, n_6104, n_6105, n_6106, n_6107;
wire n_6108, n_6109, n_6110, n_6111, n_6112, n_6114, n_6115, n_6116;
wire n_6117, n_6118, n_6120, n_6121, n_6122, n_6123, n_6126, n_6127;
wire n_6128, n_6130, n_6131, n_6132, n_6133, n_6136, n_6137, n_6138;
wire n_6139, n_6141, n_6142, n_6143, n_6146, n_6147, n_6148, n_6150;
wire n_6152, n_6153, n_6154, n_6155, n_6156, n_6157, n_6158, n_6160;
wire n_6161, n_6162, n_6163, n_6167, n_6168, n_6169, n_6171, n_6172;
wire n_6173, n_6177, n_6178, n_6179, n_6180, n_6181, n_6182, n_6183;
wire n_6184, n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191;
wire n_6192, n_6193, n_6194, n_6195, n_6196, n_6197, n_6198, n_6199;
wire n_6200, n_6201, n_6202, n_6203, n_6204, n_6205, n_6206, n_6207;
wire n_6208, n_6209, n_6210, n_6212, n_6213, n_6214, n_6215, n_6216;
wire n_6217, n_6218, n_6219, n_6220, n_6221, n_6222, n_6223, n_6224;
wire n_6225, n_6226, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232;
wire n_6422, n_6423, n_6424, n_6425, n_6428, n_6429, n_6430, n_6431;
wire n_6432, n_6433, n_6437, n_6438, n_6439, n_6440, n_6446, n_6447;
wire n_6448, n_6449, n_6450, n_6451, n_6452, n_6454, n_6455, n_6456;
wire n_6457, n_6458, n_6465, n_6466, n_6467, n_6468, n_6469, n_6471;
wire n_6472, n_6473, n_6474, n_6475, n_6479, n_6480, n_6482, n_6484;
wire n_6485, n_6486, n_6487, n_6488, n_6491, n_6492, n_6493, n_6494;
wire n_6495, n_6497, n_6501, n_6503, n_6504, n_6505, n_6507, n_6508;
wire n_6510, n_6511, n_6512, n_6513, n_6514, n_6515, n_6519, n_6520;
wire n_6521, n_6523, n_6524, n_6528, n_6529, n_6530, n_6532, n_6533;
wire n_6536, n_6537, n_6538, n_6540, n_6541, n_6544, n_6545, n_6546;
wire n_6548, n_6549, n_6550, n_6551, n_6552, n_6553, n_6555, n_6556;
wire n_6557, n_6558, n_6560, n_6561, n_6570, n_6571, n_6572, n_6573;
wire n_6575, n_6576, n_6577, n_6578, n_6580, n_6581, n_6583, n_6584;
wire n_6585, n_6586, n_6588, n_6589, n_6598, n_6599, n_6600, n_6601;
wire n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617;
wire n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6626;
wire n_6628, n_6629, n_6630, n_6631, n_6632, n_6633, n_6642, n_6643;
wire n_6644, n_6645, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663;
wire n_6664, n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671;
wire n_6672, n_6673, n_6674, n_6675, n_6676, n_6677, n_6678, n_6679;
wire n_6680, n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687;
wire n_6688, n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695;
wire n_6696, n_6697, n_6698, n_6699, n_6882, n_6883, n_6884, n_6885;
wire n_6886, n_7059, n_7060, n_7061, n_7062, n_7063, n_7064, n_7065;
wire n_7066, n_7067, n_7068, n_7069, n_7070, n_7071, n_7072, n_7073;
wire n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7080, n_7081;
wire n_7082, n_7083, n_7084, n_7085, n_7086, n_7087, n_7088, n_7089;
wire n_7090, n_7092, n_7093, n_7094, n_7281, n_7282, n_7480, n_7481;
wire n_7482, n_7483, n_7484, n_7485, n_7487, n_7488, n_7490, n_7504;
wire n_7505, n_7506, n_7507, n_7508, n_7509, n_7510, n_7511, n_8314;
wire n_8315, n_8316, n_8317, n_8318, n_8319, n_8320, n_8321, n_8322;
wire n_8323, n_8324, n_8325, n_8326, n_8327, n_8328, n_8329, n_8330;
wire n_8331, n_8332, n_8333, n_8334, n_8335, n_8336, n_8337, n_8338;
wire n_8339, n_8340, n_8341, n_8342, n_8343, n_8344, n_8345, n_8346;
wire n_8347, n_8348, n_8349, n_8350, n_8351, n_8352, n_8353, n_8354;
wire n_8355, n_8538, n_8539, n_8540, n_8541, n_8542, n_8543, n_8544;
wire n_8545, n_8546, n_8547, n_8548, n_8549, n_8550, n_8551, n_8552;
wire n_8553, n_8554, n_9384, n_9385, n_9386, n_9387, n_9388, n_9389;
wire n_9390, n_9391, n_9392, n_9393, n_9394, n_9395, n_9396, n_9397;
wire n_9398, n_9399, n_9400, n_9401, n_9402, n_9403, n_9404, n_9405;
wire n_9406, n_9407, n_9408, n_9409, n_9410, n_9411, n_9412, n_9413;
wire n_9414, n_9415, n_9416, n_9418, n_9419, n_9420, n_9421, n_9422;
wire n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430;
wire n_9431, n_9432, n_9433, n_9434, n_9435, n_9436, n_9437, n_9438;
wire n_9797, n_9798, n_9799, n_9800, n_9814, n_9815, n_9816, n_9817;
wire n_9818, n_9819, n_9820, n_9821, n_9822, n_9823, n_9824, n_10712;
wire n_10713, n_10714, n_10716, n_10717, n_10718, n_10719, n_10720,n_10721;
wire n_10722, n_10723, n_10724, n_10725, n_10726, n_10727, n_10728,n_10729;
wire n_10730, n_10731, n_10732, n_10733, n_10734, n_10735, n_10736,n_10737;
wire n_10738, n_10739, n_10740, n_10741, n_10742, n_10743, n_10744,n_10745;
wire n_10746, n_10747, n_11595, n_11596, n_11597, n_11599, n_11600,n_11601;
wire n_11602, n_11603, n_11604, n_11605, n_11607, n_11608, n_11609,n_11611;
wire n_11612, n_11613, n_11614, n_11615, n_11616, n_11617, n_11618,n_11619;
wire n_11621, n_11623, n_11625, n_11626, n_12492, n_12493, n_12494,n_15851;
wire n_15852, n_15853, n_15854, n_15855, n_15856, n_15857, n_15858,n_15859;
wire n_15860, n_15861, n_15862, n_15863, n_15864, n_15865, n_15866,n_15867;
wire n_15868;
DFFSRX1 WX651_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6173), .Q (WX651), .QN ());
NAND2X2 g55802(.A (n_6172), .B (n_4727), .Y (n_6173));
NAND2X1 g55823(.A (n_6615), .B (n_8328), .Y (n_6172));
DFFSRX1 WX653_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6169), .Q (WX653), .QN ());
OAI21X1 g55843(.A0 (n_6167), .A1 (n_5889), .B0 (n_6156), .Y (n_8328));
NAND2X2 g55841(.A (n_6168), .B (n_4725), .Y (n_6169));
NAND2X1 g55878(.A (n_6555), .B (n_8329), .Y (n_6168));
INVX1 g55905(.A (DATA_9_28), .Y (n_6167));
DFFSRX1 WX655_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6163), .Q (WX655), .QN ());
OAI21X1 g55906(.A0 (n_6162), .A1 (n_5242), .B0 (n_4070), .Y(DATA_9_28));
OAI21X1 g55903(.A0 (n_6160), .A1 (n_5889), .B0 (n_6146), .Y (n_8329));
NAND2X2 g55901(.A (n_6161), .B (n_4723), .Y (n_6163));
DFFSRX1 WX489_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6158), .Q (WX489), .QN ());
MX2X1 g55963(.A (n_6157), .B (WX491), .S0 (n_4069), .Y (n_6162));
NAND2X1 g55938(.A (n_6155), .B (n_6583), .Y (n_6161));
INVX1 g55964(.A (DATA_9_27), .Y (n_6160));
NOR2X1 g55992(.A (n_1425), .B (n_6157), .Y (n_6158));
OR2X1 g55996(.A (n_6157), .B (n_5990), .Y (n_6156));
OAI21X1 g55965(.A0 (n_6153), .A1 (n_6091), .B0 (n_4041), .Y(DATA_9_27));
DFFSRX1 WX657_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6154), .Q (WX657), .QN ());
OAI21X1 g55962(.A0 (n_6150), .A1 (n_5889), .B0 (n_6137), .Y (n_6155));
INVX1 g56007(.A (WX491), .Y (n_6157));
NAND2X2 g55960(.A (n_6152), .B (n_4722), .Y (n_6154));
DFFSRX1 WX491_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6148), .Q (WX491), .QN ());
MX2X1 g56022(.A (n_6147), .B (WX493), .S0 (n_4040), .Y (n_6153));
NAND2X2 g55997(.A (n_6583), .B (n_6882), .Y (n_6152));
INVX1 g56023(.A (DATA_9_26), .Y (n_6150));
NOR2X1 g56051(.A (n_1425), .B (n_6147), .Y (n_6148));
OR2X1 g56055(.A (n_6147), .B (n_5968), .Y (n_6146));
OAI21X1 g56024(.A0 (n_6142), .A1 (n_5242), .B0 (n_4023), .Y(DATA_9_26));
DFFSRX1 WX659_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6143), .Q (WX659), .QN ());
INVX1 g56068(.A (WX493), .Y (n_6147));
OAI21X1 g56021(.A0 (n_6141), .A1 (n_5889), .B0 (n_6126), .Y (n_6882));
DFFSRX1 WX493_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6139), .Q (WX493), .QN ());
NAND2X1 g56019(.A (n_6136), .B (n_4721), .Y (n_6143));
MX2X1 g56081(.A (n_6138), .B (WX495), .S0 (n_7066), .Y (n_6142));
INVX1 g56082(.A (DATA_9_25), .Y (n_6141));
NOR2X1 g56110(.A (n_5181), .B (n_6138), .Y (n_6139));
OR2X1 g56114(.A (n_6138), .B (n_5990), .Y (n_6137));
NAND2X1 g56056(.A (n_6555), .B (n_8330), .Y (n_6136));
OAI21X1 g56083(.A0 (n_6132), .A1 (n_6091), .B0 (n_4072), .Y(DATA_9_25));
DFFSRX1 WX661_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6133), .Q (WX661), .QN ());
OAI21X1 g56080(.A0 (n_6130), .A1 (n_5889), .B0 (n_6116), .Y (n_8330));
INVX1 g56123(.A (WX495), .Y (n_6138));
NAND2X1 g56078(.A (n_6131), .B (n_4720), .Y (n_6133));
DFFSRX1 WX495_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6128), .Q (WX495), .QN ());
MX2X1 g56140(.A (n_6127), .B (WX497), .S0 (n_4071), .Y (n_6132));
NAND2X1 g56115(.A (n_6583), .B (n_6883), .Y (n_6131));
INVX1 g56141(.A (DATA_9_24), .Y (n_6130));
NOR2X1 g56169(.A (n_5181), .B (n_6127), .Y (n_6128));
OR2X1 g56173(.A (n_6127), .B (n_5990), .Y (n_6126));
OAI21X1 g56142(.A0 (n_6122), .A1 (n_5242), .B0 (n_4055), .Y(DATA_9_24));
DFFSRX1 WX663_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6123), .Q (WX663), .QN ());
OAI21X1 g56139(.A0 (n_6120), .A1 (n_5889), .B0 (n_6095), .Y (n_6883));
INVX1 g56184(.A (WX497), .Y (n_6127));
NAND2X1 g56137(.A (n_6121), .B (n_4719), .Y (n_6123));
DFFSRX1 WX497_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6118), .Q (WX497), .QN ());
DFFSRX1 WX10993_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6115), .Q (WX10993), .QN ());
DFFSRX1 WX1942_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6114), .Q (WX1942), .QN ());
MX2X1 g56199(.A (n_6117), .B (WX499), .S0 (n_10727), .Y (n_6122));
NAND2X1 g56174(.A (n_6110), .B (n_6555), .Y (n_6121));
INVX1 g56200(.A (DATA_9_23), .Y (n_6120));
NOR2X1 g56228(.A (n_5181), .B (n_6117), .Y (n_6118));
OR2X1 g56232(.A (n_6117), .B (n_3828), .Y (n_6116));
OAI21X1 g55842(.A0 (n_3841), .A1 (n_6106), .B0 (n_6111), .Y (n_6115));
OAI21X1 g55836(.A0 (n_4283), .A1 (n_5415), .B0 (n_6112), .Y (n_6114));
OAI21X1 g56201(.A0 (n_6108), .A1 (n_6091), .B0 (n_4043), .Y(DATA_9_23));
DFFSRX1 WX665_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6109), .Q (WX665), .QN ());
OAI21X1 g55865(.A0 (n_6102), .A1 (n_4195), .B0 (n_5722), .Y (n_6112));
OAI21X1 g55866(.A0 (n_4551), .A1 (n_6177), .B0 (n_5722), .Y (n_6111));
OAI21X1 g56198(.A0 (n_6099), .A1 (n_5889), .B0 (n_6078), .Y (n_6110));
INVX1 g56243(.A (WX499), .Y (n_6117));
DFFSRX1 WX10995_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6105), .Q (WX10995), .QN ());
DFFSRX1 WX1944_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6107), .Q (WX1944), .QN ());
NAND2X1 g56196(.A (n_6100), .B (n_4717), .Y (n_6109));
DFFSRX1 WX499_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6097), .Q (WX499), .QN ());
DFFSRX1 WX10831_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6104), .Q (WX10831), .QN ());
DFFSRX1 WX1780_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6103), .Q (WX1780), .QN ());
MX2X1 g56258(.A (n_6096), .B (WX501), .S0 (n_7062), .Y (n_6108));
OAI21X1 g55896(.A0 (n_4558), .A1 (n_6106), .B0 (n_6092), .Y (n_6107));
OAI21X1 g55902(.A0 (n_3834), .A1 (n_6050), .B0 (n_6093), .Y (n_6105));
NOR2X1 g55916(.A (WX10833), .B (n_1648), .Y (n_6104));
NOR2X1 g55920(.A (WX1782), .B (n_5181), .Y (n_6103));
NOR2X1 g55923(.A (WX1782), .B (n_5500), .Y (n_6102));
NOR2X1 g55924(.A (WX10833), .B (n_5811), .Y (n_6177));
NAND2X1 g56233(.A (n_6090), .B (n_6583), .Y (n_6100));
INVX1 g56259(.A (DATA_9_22), .Y (n_6099));
NOR2X1 g56287(.A (n_2849), .B (n_6096), .Y (n_6097));
OR2X1 g56291(.A (n_6096), .B (n_5990), .Y (n_6095));
OAI21X1 g55926(.A0 (n_4549), .A1 (n_6184), .B0 (n_5722), .Y (n_6093));
OAI21X1 g55925(.A0 (n_6083), .A1 (n_4193), .B0 (n_4947), .Y (n_6092));
OAI21X1 g56260(.A0 (n_6081), .A1 (n_6091), .B0 (n_4033), .Y(DATA_9_22));
DFFSRX1 WX10997_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6087), .Q (WX10997), .QN ());
DFFSRX1 WX1946_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6088), .Q (WX1946), .QN ());
DFFSRX1 WX667_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6086), .Q (WX667), .QN ());
DFFSRX1 WX10833_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6085), .Q (), .QN (WX10833));
DFFSRX1 WX1782_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6084), .Q (), .QN (WX1782));
OAI21X1 g56257(.A0 (n_6072), .A1 (n_5889), .B0 (n_6053), .Y (n_6090));
INVX1 g56303(.A (WX501), .Y (n_6096));
OAI21X1 g55955(.A0 (n_4556), .A1 (n_5600), .B0 (n_6076), .Y (n_6088));
OAI21X1 g55961(.A0 (n_3839), .A1 (n_6106), .B0 (n_6075), .Y (n_6087));
NAND2X1 g56255(.A (n_6074), .B (n_4716), .Y (n_6086));
DFFSRX1 WX501_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6080), .Q (WX501), .QN ());
NOR2X1 g55975(.A (WX10835), .B (n_2605), .Y (n_6085));
NOR2X1 g55978(.A (WX1784), .B (n_1648), .Y (n_6084));
NOR2X1 g55982(.A (WX1784), .B (n_5479), .Y (n_6083));
NOR2X1 g55984(.A (WX10835), .B (n_5811), .Y (n_6184));
MX2X1 g56317(.A (n_6079), .B (WX503), .S0 (n_7070), .Y (n_6081));
NOR2X1 g56346(.A (n_5181), .B (n_6079), .Y (n_6080));
OR2X1 g56350(.A (n_6079), .B (n_5990), .Y (n_6078));
OAI21X1 g55983(.A0 (n_6064), .A1 (n_4191), .B0 (n_5460), .Y (n_6076));
OAI21X1 g55987(.A0 (n_4547), .A1 (n_6209), .B0 (n_5619), .Y (n_6075));
NAND2X1 g56292(.A (n_6068), .B (n_6615), .Y (n_6074));
DFFSRX1 WX10999_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6069), .Q (WX10999), .QN ());
DFFSRX1 WX1948_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6070), .Q (WX1948), .QN ());
INVX1 g56318(.A (DATA_9_21), .Y (n_6072));
DFFSRX1 WX10835_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6067), .Q (), .QN (WX10835));
DFFSRX1 WX1784_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6066), .Q (), .QN (WX1784));
DFFSRX1 WX669_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6063), .Q (WX669), .QN ());
OAI21X1 g56319(.A0 (n_6061), .A1 (n_6091), .B0 (n_4025), .Y(DATA_9_21));
INVX1 g56362(.A (WX503), .Y (n_6079));
OAI21X1 g56014(.A0 (n_4554), .A1 (n_4803), .B0 (n_6060), .Y (n_6070));
OAI21X1 g56020(.A0 (n_3837), .A1 (n_5482), .B0 (n_6059), .Y (n_6069));
OAI21X1 g56316(.A0 (n_6057), .A1 (n_5889), .B0 (n_6033), .Y (n_6068));
DFFSRX1 WX503_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6055), .Q (WX503), .QN ());
NOR2X1 g56034(.A (WX10837), .B (n_1648), .Y (n_6067));
NOR2X1 g56036(.A (WX1786), .B (n_2605), .Y (n_6066));
NOR2X1 g56041(.A (WX1786), .B (n_5811), .Y (n_6064));
NAND2X1 g56314(.A (n_6058), .B (n_4715), .Y (n_6063));
NOR2X1 g56045(.A (WX10837), .B (n_5811), .Y (n_6209));
MX2X1 g56376(.A (n_6054), .B (WX505), .S0 (n_6553), .Y (n_6061));
DFFSRX1 WX11001_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6051), .Q (WX11001), .QN ());
DFFSRX1 WX1950_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6052), .Q (WX1950), .QN ());
OAI21X1 g56044(.A0 (n_6046), .A1 (n_4188), .B0 (n_4860), .Y (n_6060));
OAI21X1 g56048(.A0 (n_4545), .A1 (n_6210), .B0 (n_5460), .Y (n_6059));
DFFSRX1 WX10837_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6048), .Q (), .QN (WX10837));
NAND2X1 g56351(.A (n_6555), .B (n_8331), .Y (n_6058));
DFFSRX1 WX1786_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6047), .Q (), .QN (WX1786));
INVX1 g56377(.A (DATA_9_20), .Y (n_6057));
NOR2X1 g56405(.A (n_2849), .B (n_6054), .Y (n_6055));
OR2X1 g56409(.A (n_6054), .B (n_5990), .Y (n_6053));
OAI21X1 g56073(.A0 (n_4522), .A1 (n_5928), .B0 (n_6042), .Y (n_6052));
OAI21X1 g56378(.A0 (n_6040), .A1 (n_5242), .B0 (n_4082), .Y(DATA_9_20));
OAI21X1 g56079(.A0 (n_3822), .A1 (n_6050), .B0 (n_6041), .Y (n_6051));
DFFSRX1 WX671_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6043), .Q (WX671), .QN ());
OAI21X1 g56375(.A0 (n_6038), .A1 (n_5889), .B0 (n_6013), .Y (n_8331));
NOR2X1 g56093(.A (WX10839), .B (n_2620), .Y (n_6048));
NOR2X1 g56095(.A (WX1788), .B (n_5181), .Y (n_6047));
INVX1 g56423(.A (WX505), .Y (n_6054));
NOR2X1 g56102(.A (WX1788), .B (n_5811), .Y (n_6046));
NOR2X1 g56106(.A (WX10839), .B (n_5811), .Y (n_6210));
NAND2X1 g56373(.A (n_6039), .B (n_4714), .Y (n_6043));
DFFSRX1 WX505_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6036), .Q (WX505), .QN ());
OAI21X1 g56105(.A0 (n_6027), .A1 (n_4186), .B0 (n_5722), .Y (n_6042));
OAI21X1 g56107(.A0 (n_4543), .A1 (n_6178), .B0 (n_4860), .Y (n_6041));
DFFSRX1 WX11003_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6031), .Q (WX11003), .QN ());
DFFSRX1 WX1952_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6032), .Q (WX1952), .QN ());
MX2X1 g56435(.A (n_6034), .B (WX507), .S0 (n_6645), .Y (n_6040));
DFFSRX1 WX10839_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6030), .Q (), .QN (WX10839));
DFFSRX1 WX1788_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6029), .Q (), .QN (WX1788));
NAND2X1 g56410(.A (n_6025), .B (n_6583), .Y (n_6039));
INVX1 g56436(.A (DATA_9_19), .Y (n_6038));
NOR2X1 g56464(.A (n_5181), .B (n_6034), .Y (n_6036));
OR2X1 g56468(.A (n_6034), .B (n_5990), .Y (n_6033));
OAI21X1 g56133(.A0 (n_4496), .A1 (n_5918), .B0 (n_6024), .Y (n_6032));
OAI21X1 g56138(.A0 (n_3836), .A1 (n_5879), .B0 (n_6023), .Y (n_6031));
OAI21X1 g56437(.A0 (n_6021), .A1 (n_5843), .B0 (n_4075), .Y(DATA_9_19));
NOR2X1 g56152(.A (WX10841), .B (n_1648), .Y (n_6030));
NOR2X1 g56154(.A (WX1790), .B (n_1648), .Y (n_6029));
NOR2X1 g56163(.A (WX1790), .B (n_5822), .Y (n_6027));
NOR2X1 g56165(.A (WX10841), .B (n_5479), .Y (n_6178));
DFFSRX1 WX673_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6022), .Q (WX673), .QN ());
OAI21X1 g56434(.A0 (n_6017), .A1 (n_5889), .B0 (n_5991), .Y (n_6025));
INVX1 g56477(.A (WX507), .Y (n_6034));
OAI21X1 g56164(.A0 (n_6010), .A1 (n_4183), .B0 (n_5566), .Y (n_6024));
OAI21X1 g56166(.A0 (n_4541), .A1 (n_6179), .B0 (n_5722), .Y (n_6023));
DFFSRX1 WX11005_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6019), .Q (WX11005), .QN ());
DFFSRX1 WX1954_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6020), .Q (WX1954), .QN ());
NAND2X1 g56432(.A (n_15853), .B (n_15854), .Y (n_6022));
DFFSRX1 WX507_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6015), .Q (WX507), .QN ());
DFFSRX1 WX10841_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6012), .Q (), .QN (WX10841));
DFFSRX1 WX1790_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6011), .Q (), .QN (WX1790));
MX2X1 g56494(.A (n_6014), .B (WX509), .S0 (n_10731), .Y (n_6021));
OAI21X1 g56192(.A0 (n_4488), .A1 (n_5834), .B0 (n_6008), .Y (n_6020));
OAI21X1 g56197(.A0 (n_3827), .A1 (n_5841), .B0 (n_6007), .Y (n_6019));
NAND2X1 g56469(.A (n_6615), .B (n_8332), .Y (n_15854));
INVX1 g56495(.A (DATA_9_18), .Y (n_6017));
NOR2X1 g56523(.A (n_1425), .B (n_6014), .Y (n_6015));
OR2X1 g56527(.A (n_6014), .B (n_5968), .Y (n_6013));
NOR2X1 g56211(.A (WX10843), .B (n_5712), .Y (n_6012));
NOR2X1 g56213(.A (WX1792), .B (n_2620), .Y (n_6011));
NOR2X1 g56222(.A (WX1792), .B (n_5427), .Y (n_6010));
NOR2X1 g56224(.A (WX10843), .B (n_5822), .Y (n_6179));
OAI21X1 g56496(.A0 (n_6001), .A1 (n_5965), .B0 (n_4064), .Y(DATA_9_18));
OAI21X1 g56223(.A0 (n_5998), .A1 (n_4181), .B0 (n_4860), .Y (n_6008));
OAI21X1 g56225(.A0 (n_4537), .A1 (n_6439), .B0 (n_6497), .Y (n_6007));
DFFSRX1 WX11007_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6002), .Q (WX11007), .QN ());
DFFSRX1 WX1956_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6003), .Q (WX1956), .QN ());
DFFSRX1 WX675_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6004), .Q (WX675), .QN ());
OAI21X1 g56493(.A0 (n_5995), .A1 (n_5889), .B0 (n_5969), .Y (n_8332));
INVX1 g56536(.A (WX509), .Y (n_6014));
DFFSRX1 WX10843_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6000), .Q (), .QN (WX10843));
DFFSRX1 WX1792_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5999), .Q (), .QN (WX1792));
NAND2X2 g56491(.A (n_5996), .B (n_4711), .Y (n_6004));
DFFSRX1 WX509_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5993), .Q (WX509), .QN ());
OAI21X1 g56251(.A0 (n_4253), .A1 (n_5439), .B0 (n_5989), .Y (n_6003));
OAI21X1 g56256(.A0 (n_3830), .A1 (n_5845), .B0 (n_5988), .Y (n_6002));
MX2X1 g56553(.A (n_5992), .B (WX511), .S0 (n_7074), .Y (n_6001));
NOR2X1 g56270(.A (WX10845), .B (n_1648), .Y (n_6000));
NOR2X1 g56272(.A (WX1794), .B (n_5181), .Y (n_5999));
NOR2X1 g56281(.A (WX1794), .B (n_5662), .Y (n_5998));
NAND2X1 g56528(.A (n_5987), .B (n_6575), .Y (n_5996));
INVX1 g56554(.A (DATA_9_17), .Y (n_5995));
NOR2X1 g56582(.A (n_1425), .B (n_5992), .Y (n_5993));
OR2X1 g56587(.A (n_5992), .B (n_5990), .Y (n_5991));
OAI21X1 g56282(.A0 (n_5981), .A1 (n_4179), .B0 (n_5566), .Y (n_5989));
OAI21X1 g56285(.A0 (n_4625), .A1 (n_6216), .B0 (n_4860), .Y (n_5988));
DFFSRX1 WX11009_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5985), .Q (WX11009), .QN ());
DFFSRX1 WX1958_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5986), .Q (WX1958), .QN ());
OAI21X1 g56555(.A0 (n_5978), .A1 (n_5965), .B0 (n_4057), .Y(DATA_9_17));
DFFSRX1 WX677_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6524), .Q (WX677), .QN ());
DFFSRX1 WX10845_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5983), .Q (), .QN (WX10845));
DFFSRX1 WX1794_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5982), .Q (), .QN (WX1794));
OAI21X1 g56552(.A0 (n_5973), .A1 (n_5889), .B0 (n_5940), .Y (n_5987));
INVX1 g56597(.A (WX511), .Y (n_5992));
OAI21X1 g56310(.A0 (n_4251), .A1 (n_5630), .B0 (n_5977), .Y (n_5986));
OAI21X1 g56315(.A0 (n_3833), .A1 (n_5882), .B0 (n_5976), .Y (n_5985));
DFFSRX1 WX511_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5971), .Q (WX511), .QN ());
DFFSRX1 WX9718_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5974), .Q (WX9718), .QN ());
NOR2X1 g56329(.A (WX10847), .B (n_5712), .Y (n_5983));
NOR2X1 g56331(.A (WX1796), .B (n_1425), .Y (n_5982));
NOR2X1 g56340(.A (WX1796), .B (n_5662), .Y (n_5981));
NOR2X1 g56342(.A (WX10847), .B (n_5811), .Y (n_6216));
MX2X1 g56612(.A (n_5970), .B (WX513), .S0 (n_9800), .Y (n_5978));
DFFSRX1 WX11011_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5966), .Q (WX11011), .QN ());
DFFSRX1 WX1960_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5967), .Q (WX1960), .QN ());
OAI21X1 g56341(.A0 (n_5961), .A1 (n_4176), .B0 (n_7087), .Y (n_5977));
OAI21X1 g56345(.A0 (n_4535), .A1 (n_6217), .B0 (n_5722), .Y (n_5976));
DFFSRX1 WX10847_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5964), .Q (), .QN (WX10847));
DFFSRX1 WX1796_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5963), .Q (), .QN (WX1796));
OAI21X1 g55798(.A0 (n_4534), .A1 (n_5183), .B0 (n_5959), .Y (n_5974));
INVX1 g56613(.A (DATA_9_16), .Y (n_5973));
NOR2X1 g56641(.A (n_1425), .B (n_5970), .Y (n_5971));
OR2X1 g56647(.A (n_5970), .B (n_5968), .Y (n_5969));
OAI21X1 g56369(.A0 (n_4474), .A1 (n_5418), .B0 (n_5956), .Y (n_5967));
OAI21X1 g56374(.A0 (n_3819), .A1 (n_5892), .B0 (n_5954), .Y (n_5966));
OAI21X1 g56614(.A0 (n_5951), .A1 (n_5965), .B0 (n_4049), .Y(DATA_9_16));
DFFSRX1 WX679_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6561), .Q (WX679), .QN ());
NOR2X1 g56388(.A (WX10849), .B (n_5712), .Y (n_5964));
NOR2X1 g56390(.A (WX1798), .B (n_1648), .Y (n_5963));
NOR2X1 g56399(.A (WX1798), .B (n_5427), .Y (n_5961));
NOR2X1 g56403(.A (WX10849), .B (n_5479), .Y (n_6217));
OAI21X1 g55820(.A0 (n_4592), .A1 (n_6218), .B0 (n_3183), .Y (n_5959));
INVX1 g56656(.A (WX513), .Y (n_5970));
DFFSRX1 WX8427_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5952), .Q (WX8427), .QN ());
DFFSRX1 WX9720_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5950), .Q (WX9720), .QN ());
OAI21X1 g56400(.A0 (n_5936), .A1 (n_4174), .B0 (n_5722), .Y (n_5956));
OAI21X1 g56404(.A0 (n_4533), .A1 (n_6180), .B0 (n_5722), .Y (n_5954));
DFFSRX1 WX513_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5942), .Q (WX513), .QN ());
DFFSRX1 WX9556_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5947), .Q (WX9556), .QN ());
DFFSRX1 WX11013_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5948), .Q (WX11013), .QN ());
DFFSRX1 WX1962_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5949), .Q (WX1962), .QN ());
OAI21X1 g55797(.A0 (n_4591), .A1 (n_5886), .B0 (n_5939), .Y (n_5952));
DFFSRX1 WX10849_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5938), .Q (), .QN (WX10849));
DFFSRX1 WX1798_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5937), .Q (), .QN (WX1798));
MX2X1 g56671(.A (n_5941), .B (WX515), .S0 (n_7078), .Y (n_5951));
OAI21X1 g55837(.A0 (n_4532), .A1 (n_5892), .B0 (n_5934), .Y (n_5950));
OAI21X1 g56428(.A0 (n_4464), .A1 (n_5879), .B0 (n_5933), .Y (n_5949));
OAI21X1 g56433(.A0 (n_3844), .A1 (n_5928), .B0 (n_5931), .Y (n_5948));
AND2X1 g55867(.A (WX9558), .B (n_2383), .Y (n_5947));
AND2X1 g55869(.A (WX9558), .B (n_5828), .Y (n_6218));
INVX1 g56672(.A (DATA_9_15), .Y (n_5944));
NOR2X1 g56700(.A (n_1425), .B (n_5941), .Y (n_5942));
OR2X1 g56706(.A (n_5941), .B (n_4882), .Y (n_5940));
OAI21X1 g55818(.A0 (n_4364), .A1 (n_6658), .B0 (n_5619), .Y (n_5939));
NOR2X1 g56447(.A (WX10851), .B (n_1425), .Y (n_5938));
NOR2X1 g56449(.A (WX1800), .B (n_1648), .Y (n_5937));
NOR2X1 g56458(.A (WX1800), .B (n_5838), .Y (n_5936));
NOR2X1 g56462(.A (WX10851), .B (n_5479), .Y (n_6180));
OAI21X1 g55870(.A0 (n_4590), .A1 (n_6185), .B0 (n_5556), .Y (n_5934));
OAI21X1 g56673(.A0 (n_5917), .A1 (n_5242), .B0 (n_4045), .Y(DATA_9_15));
DFFSRX1 WX7136_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5929), .Q (WX7136), .QN ());
DFFSRX1 WX8429_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5925), .Q (WX8429), .QN ());
DFFSRX1 WX9722_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5926), .Q (WX9722), .QN ());
DFFSRX1 WX681_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5927), .Q (WX681), .QN ());
OAI21X1 g56459(.A0 (n_5910), .A1 (n_4172), .B0 (n_5722), .Y (n_5933));
OAI21X1 g56463(.A0 (n_4531), .A1 (n_6214), .B0 (n_4860), .Y (n_5931));
DFFSRX1 WX9558_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5924), .Q (WX9558), .QN ());
INVX1 g56715(.A (WX515), .Y (n_5941));
DFFSRX1 WX8265_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5922), .Q (WX8265), .QN ());
DFFSRX1 WX11015_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5919), .Q (WX11015), .QN ());
DFFSRX1 WX1964_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5921), .Q (WX1964), .QN ());
DFFSRX1 WX10851_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5914), .Q (), .QN (WX10851));
DFFSRX1 WX1800_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5912), .Q (), .QN (WX1800));
OAI21X1 g55801(.A0 (n_4363), .A1 (n_5928), .B0 (n_5907), .Y (n_5929));
NAND2X1 g56668(.A (n_5905), .B (n_4706), .Y (n_5927));
DFFSRX1 WX515_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5901), .Q (WX515), .QN ());
OAI21X1 g55897(.A0 (n_4530), .A1 (n_5598), .B0 (n_5916), .Y (n_5926));
OAI21X1 g55835(.A0 (n_4589), .A1 (n_5493), .B0 (n_5915), .Y (n_5925));
NOR2X1 g55927(.A (WX9560), .B (n_5712), .Y (n_5924));
NOR2X1 g55929(.A (WX9560), .B (n_5479), .Y (n_6185));
AND2X1 g55858(.A (WX8267), .B (n_2396), .Y (n_5922));
OAI21X1 g56487(.A0 (n_4241), .A1 (n_5830), .B0 (n_5896), .Y (n_5921));
AND2X1 g55861(.A (WX8267), .B (n_5873), .Y (n_6658));
OAI21X1 g56492(.A0 (n_3812), .A1 (n_5918), .B0 (n_5894), .Y (n_5919));
MX2X1 g56730(.A (n_5899), .B (WX517), .S0 (n_4044), .Y (n_5917));
OAI21X1 g55930(.A0 (n_4588), .A1 (n_6187), .B0 (n_5460), .Y (n_5916));
OAI21X1 g55862(.A0 (n_5884), .A1 (n_4362), .B0 (n_5722), .Y (n_5915));
NOR2X1 g56507(.A (WX10853), .B (n_5712), .Y (n_5914));
NOR2X1 g56508(.A (WX1802), .B (n_5712), .Y (n_5912));
NOR2X1 g56517(.A (WX1802), .B (n_5500), .Y (n_5910));
NOR2X1 g56521(.A (WX10853), .B (n_5500), .Y (n_6214));
OAI21X1 g55824(.A0 (n_4413), .A1 (n_6186), .B0 (n_5722), .Y (n_5907));
NAND2X1 g56707(.A (n_5890), .B (n_6575), .Y (n_5905));
INVX1 g56731(.A (DATA_9_14), .Y (n_5903));
NOR2X1 g56758(.A (n_1425), .B (n_5899), .Y (n_5901));
OR2X1 g56764(.A (n_5899), .B (n_5968), .Y (n_5898));
DFFSRX1 WX5845_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5893), .Q (WX5845), .QN ());
DFFSRX1 WX7138_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5887), .Q (WX7138), .QN ());
DFFSRX1 WX8431_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5888), .Q (WX8431), .QN ());
DFFSRX1 WX9724_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5891), .Q (WX9724), .QN ());
DFFSRX1 WX9560_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5878), .Q (), .QN (WX9560));
OAI21X1 g56518(.A0 (n_5865), .A1 (n_4170), .B0 (n_4947), .Y (n_5896));
OAI21X1 g56522(.A0 (n_4529), .A1 (n_6215), .B0 (n_7087), .Y (n_5894));
DFFSRX1 WX8267_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5885), .Q (WX8267), .QN ());
OAI21X1 g56732(.A0 (n_5858), .A1 (n_5965), .B0 (n_4039), .Y(DATA_9_14));
DFFSRX1 WX4554_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5883), .Q (WX4554), .QN ());
DFFSRX1 WX6974_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5876), .Q (WX6974), .QN ());
DFFSRX1 WX11017_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5880), .Q (WX11017), .QN ());
DFFSRX1 WX1966_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5881), .Q (WX1966), .QN ());
DFFSRX1 WX683_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5872), .Q (WX683), .QN ());
OAI21X1 g55800(.A0 (n_4412), .A1 (n_5892), .B0 (n_5869), .Y (n_5893));
OAI21X1 g55956(.A0 (n_4273), .A1 (n_5841), .B0 (n_5862), .Y (n_5891));
DFFSRX1 WX10853_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5867), .Q (), .QN (WX10853));
DFFSRX1 WX1802_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5866), .Q (), .QN (WX1802));
OAI21X1 g56729(.A0 (n_5853), .A1 (n_5889), .B0 (n_5790), .Y (n_5890));
OAI21X1 g55895(.A0 (n_4303), .A1 (n_5750), .B0 (n_5871), .Y (n_5888));
INVX1 g56775(.A (WX517), .Y (n_5899));
OAI21X1 g55840(.A0 (n_4361), .A1 (n_5886), .B0 (n_5860), .Y (n_5887));
NOR2X1 g55917(.A (WX8269), .B (n_5712), .Y (n_5885));
NOR2X1 g55921(.A (WX8269), .B (n_5838), .Y (n_5884));
OAI21X1 g55799(.A0 (n_4478), .A1 (n_5882), .B0 (n_5857), .Y (n_5883));
OAI21X1 g56547(.A0 (n_4460), .A1 (n_5235), .B0 (n_5856), .Y (n_5881));
OAI21X1 g56551(.A0 (n_3829), .A1 (n_5879), .B0 (n_5855), .Y (n_5880));
NOR2X1 g55985(.A (WX9562), .B (n_1648), .Y (n_5878));
AND2X1 g55879(.A (WX6976), .B (n_2383), .Y (n_5876));
NOR2X1 g55988(.A (WX9562), .B (n_5811), .Y (n_6187));
AND2X1 g55881(.A (WX6976), .B (n_5873), .Y (n_6186));
NAND2X2 g56727(.A (n_5854), .B (n_4704), .Y (n_5872));
DFFSRX1 WX517_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5851), .Q (WX517), .QN ());
OAI21X1 g55922(.A0 (n_4360), .A1 (n_6189), .B0 (n_5722), .Y (n_5871));
OAI21X1 g55822(.A0 (n_4479), .A1 (n_6188), .B0 (n_5566), .Y (n_5869));
NOR2X1 g56567(.A (WX10855), .B (n_2851), .Y (n_5867));
NOR2X1 g56568(.A (WX1804), .B (n_2851), .Y (n_5866));
NOR2X1 g56577(.A (WX1804), .B (n_5427), .Y (n_5865));
NOR2X1 g56581(.A (WX10855), .B (n_5811), .Y (n_6215));
OAI21X1 g55989(.A0 (n_5823), .A1 (n_4302), .B0 (n_6497), .Y (n_5862));
OAI21X1 g55882(.A0 (n_4411), .A1 (n_6665), .B0 (n_5619), .Y (n_5860));
MX2X1 g56789(.A (n_5849), .B (WX519), .S0 (n_4038), .Y (n_5858));
DFFSRX1 WX5847_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5842), .Q (WX5847), .QN ());
DFFSRX1 WX7140_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5844), .Q (WX7140), .QN ());
DFFSRX1 WX8433_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5847), .Q (WX8433), .QN ());
DFFSRX1 WX9726_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5846), .Q (WX9726), .QN ());
DFFSRX1 WX8269_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5837), .Q (), .QN (WX8269));
OAI21X1 g55821(.A0 (n_4623), .A1 (n_6219), .B0 (n_5556), .Y (n_5857));
OAI21X1 g56580(.A0 (n_5813), .A1 (n_4168), .B0 (n_5460), .Y (n_5856));
OAI21X1 g56583(.A0 (n_5812), .A1 (n_4272), .B0 (n_5722), .Y (n_5855));
DFFSRX1 WX9562_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5824), .Q (), .QN (WX9562));
DFFSRX1 WX6976_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5840), .Q (WX6976), .QN ());
NAND2X1 g56765(.A (n_6575), .B (n_8333), .Y (n_5854));
INVX1 g56790(.A (DATA_9_13), .Y (n_5853));
DFFSRX1 WX4556_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5826), .Q (WX4556), .QN ());
DFFSRX1 WX5683_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5833), .Q (WX5683), .QN ());
NOR2X1 g56815(.A (n_5181), .B (n_5849), .Y (n_5851));
DFFSRX1 WX1968_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5835), .Q (WX1968), .QN ());
DFFSRX1 WX11019_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5831), .Q (WX11019), .QN ());
OR2X1 g56822(.A (n_5849), .B (n_5990), .Y (n_5848));
OAI21X1 g55954(.A0 (n_4584), .A1 (n_5825), .B0 (n_5818), .Y (n_5847));
DFFSRX1 WX10855_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5816), .Q (), .QN (WX10855));
DFFSRX1 WX1804_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5815), .Q (), .QN (WX1804));
OAI21X1 g56015(.A0 (n_4526), .A1 (n_5845), .B0 (n_5809), .Y (n_5846));
OAI21X1 g55900(.A0 (n_4357), .A1 (n_5879), .B0 (n_5821), .Y (n_5844));
OAI21X1 g56791(.A0 (n_5803), .A1 (n_5843), .B0 (n_4035), .Y(DATA_9_13));
DFFSRX1 WX4392_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5820), .Q (WX4392), .QN ());
DFFSRX1 WX685_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6533), .Q (WX685), .QN ());
OAI21X1 g55839(.A0 (n_4410), .A1 (n_5841), .B0 (n_5814), .Y (n_5842));
NOR2X1 g55939(.A (WX6978), .B (n_2620), .Y (n_5840));
NOR2X1 g55941(.A (WX6978), .B (n_5838), .Y (n_6665));
NOR2X1 g55976(.A (WX8271), .B (n_2620), .Y (n_5837));
OAI21X1 g56607(.A0 (n_4452), .A1 (n_5834), .B0 (n_5806), .Y (n_5835));
AND2X1 g55874(.A (WX5685), .B (n_2378), .Y (n_5833));
NOR2X1 g55980(.A (WX8271), .B (n_5838), .Y (n_6189));
OAI21X1 g56610(.A0 (n_3826), .A1 (n_5830), .B0 (n_5804), .Y (n_5831));
AND2X1 g55875(.A (WX5685), .B (n_5828), .Y (n_6188));
OAI21X1 g56788(.A0 (n_5796), .A1 (n_5889), .B0 (n_5743), .Y (n_8333));
OAI21X1 g55838(.A0 (n_4476), .A1 (n_5825), .B0 (n_5807), .Y (n_5826));
INVX1 g56834(.A (WX519), .Y (n_5849));
NOR2X1 g56042(.A (WX9564), .B (n_5712), .Y (n_5824));
NOR2X1 g56046(.A (WX9564), .B (n_5822), .Y (n_5823));
OAI21X1 g55942(.A0 (n_4409), .A1 (n_6671), .B0 (n_5556), .Y (n_5821));
AND2X1 g55868(.A (WX4394), .B (n_2529), .Y (n_5820));
AND2X1 g55871(.A (WX4394), .B (n_5828), .Y (n_6219));
OAI21X1 g55981(.A0 (n_4356), .A1 (n_6220), .B0 (n_5722), .Y (n_5818));
NOR2X1 g56627(.A (WX10857), .B (n_3188), .Y (n_5816));
NOR2X1 g56628(.A (WX1806), .B (n_1648), .Y (n_5815));
OAI21X1 g55876(.A0 (n_4477), .A1 (n_6190), .B0 (n_4860), .Y (n_5814));
NOR2X1 g56639(.A (WX1806), .B (n_5427), .Y (n_5813));
NOR2X1 g56642(.A (WX10857), .B (n_5811), .Y (n_5812));
DFFSRX1 WX3263_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5794), .Q (WX3263), .QN ());
DFFSRX1 WX5849_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5798), .Q (WX5849), .QN ());
DFFSRX1 WX7142_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5801), .Q (WX7142), .QN ());
DFFSRX1 WX8435_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5800), .Q (WX8435), .QN ());
DFFSRX1 WX9728_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5802), .Q (WX9728), .QN ());
DFFSRX1 WX519_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5792), .Q (WX519), .QN ());
OAI21X1 g56047(.A0 (n_4583), .A1 (n_6659), .B0 (n_5722), .Y (n_5809));
DFFSRX1 WX9564_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5789), .Q (), .QN (WX9564));
DFFSRX1 WX6978_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5781), .Q (), .QN (WX6978));
OAI21X1 g55872(.A0 (n_5771), .A1 (n_9405), .B0 (n_5556), .Y (n_5807));
OAI21X1 g56640(.A0 (n_5765), .A1 (n_4166), .B0 (n_5460), .Y (n_5806));
OAI21X1 g56644(.A0 (n_4525), .A1 (n_6181), .B0 (n_5722), .Y (n_5804));
DFFSRX1 WX8271_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5776), .Q (), .QN (WX8271));
DFFSRX1 WX5685_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5788), .Q (WX5685), .QN ());
DFFSRX1 WX4558_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5777), .Q (WX4558), .QN ());
DFFSRX1 WX11021_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_7094), .Q (WX11021), .QN ());
DFFSRX1 WX1970_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5784), .Q (WX1970), .QN ());
MX2X1 g56848(.A (n_5791), .B (WX521), .S0 (n_6573), .Y (n_5803));
OAI21X1 g56074(.A0 (n_4271), .A1 (n_5841), .B0 (n_5769), .Y (n_5802));
OAI21X1 g55959(.A0 (n_4123), .A1 (n_5576), .B0 (n_5766), .Y (n_5801));
DFFSRX1 WX10857_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5768), .Q (), .QN (WX10857));
DFFSRX1 WX1806_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5767), .Q (), .QN (WX1806));
DFFSRX1 WX4394_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5773), .Q (WX4394), .QN ());
OAI21X1 g56013(.A0 (n_4582), .A1 (n_5439), .B0 (n_5763), .Y (n_5800));
OAI21X1 g55899(.A0 (n_4408), .A1 (n_5549), .B0 (n_5770), .Y (n_5798));
INVX1 g56849(.A (DATA_9_12), .Y (n_5796));
OAI21X1 g55795(.A0 (n_4622), .A1 (n_5183), .B0 (n_5774), .Y (n_5794));
NOR2X1 g56873(.A (n_5181), .B (n_5791), .Y (n_5792));
OR2X1 g56881(.A (n_5791), .B (n_5968), .Y (n_5790));
NOR2X1 g56100(.A (WX9566), .B (n_5181), .Y (n_5789));
NOR2X1 g55934(.A (WX5687), .B (n_5181), .Y (n_5788));
NOR2X1 g55935(.A (WX5687), .B (n_5838), .Y (n_6190));
NOR2X1 g56103(.A (WX9566), .B (n_5500), .Y (n_6659));
OAI21X1 g56666(.A0 (n_4231), .A1 (n_5468), .B0 (n_5759), .Y (n_5784));
NOR2X1 g55998(.A (WX6980), .B (n_2620), .Y (n_5781));
NOR2X1 g56000(.A (WX6980), .B (n_5838), .Y (n_6671));
OAI21X1 g55898(.A0 (n_4249), .A1 (n_5892), .B0 (n_5760), .Y (n_5777));
DFFSRX1 WX687_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5755), .Q (WX687), .QN ());
NOR2X1 g56035(.A (WX8273), .B (n_1425), .Y (n_5776));
NOR2X1 g56039(.A (WX8273), .B (n_5500), .Y (n_6220));
OAI21X1 g56850(.A0 (n_5748), .A1 (n_5709), .B0 (n_4029), .Y(DATA_9_12));
OAI21X1 g55816(.A0 (n_4230), .A1 (n_8538), .B0 (n_4860), .Y (n_5774));
NOR2X1 g55928(.A (WX4396), .B (n_5712), .Y (n_5773));
NOR2X1 g55931(.A (WX4396), .B (n_5479), .Y (n_5771));
OAI21X1 g55936(.A0 (n_5732), .A1 (n_9421), .B0 (n_4860), .Y (n_5770));
OAI21X1 g56104(.A0 (n_4581), .A1 (n_6685), .B0 (n_5722), .Y (n_5769));
NOR2X1 g56686(.A (WX10859), .B (n_5181), .Y (n_5768));
NOR2X1 g56687(.A (WX1808), .B (n_3188), .Y (n_5767));
OAI21X1 g56001(.A0 (n_5747), .A1 (n_9423), .B0 (n_5706), .Y (n_5766));
NOR2X1 g56698(.A (WX1808), .B (n_4882), .Y (n_5765));
NOR2X1 g56702(.A (WX10859), .B (n_5838), .Y (n_6181));
DFFSRX1 WX3265_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5751), .Q (WX3265), .QN ());
DFFSRX1 WX5851_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5752), .Q (WX5851), .QN ());
DFFSRX1 WX7144_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5749), .Q (WX7144), .QN ());
DFFSRX1 WX8437_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5754), .Q (WX8437), .QN ());
DFFSRX1 WX9730_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5753), .Q (WX9730), .QN ());
OAI21X1 g56040(.A0 (n_4122), .A1 (n_9814), .B0 (n_4947), .Y (n_5763));
INVX1 g56893(.A (WX521), .Y (n_5791));
DFFSRX1 WX8273_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5742), .Q (), .QN (WX8273));
OAI21X1 g55932(.A0 (n_15855), .A1 (n_15856), .B0 (n_5722), .Y(n_5760));
DFFSRX1 WX5687_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5733), .Q (), .QN (WX5687));
DFFSRX1 WX9566_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5737), .Q (), .QN (WX9566));
OAI21X1 g56699(.A0 (n_5711), .A1 (n_4164), .B0 (n_4860), .Y (n_5759));
DFFSRX1 WX6980_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5725), .Q (), .QN (WX6980));
DFFSRX1 WX3101_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5735), .Q (WX3101), .QN ());
DFFSRX1 WX4560_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5738), .Q (WX4560), .QN ());
DFFSRX1 WX11023_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5730), .Q (WX11023), .QN ());
DFFSRX1 WX1972_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5731), .Q (WX1972), .QN ());
NAND2X1 g56845(.A (n_5728), .B (n_4702), .Y (n_5755));
DFFSRX1 WX521_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5745), .Q (WX521), .QN ());
OAI21X1 g56072(.A0 (n_4577), .A1 (n_4868), .B0 (n_5723), .Y (n_5754));
DFFSRX1 WX4396_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5719), .Q (), .QN (WX4396));
OAI21X1 g56132(.A0 (n_4524), .A1 (n_5825), .B0 (n_5720), .Y (n_5753));
OAI21X1 g55958(.A0 (n_4406), .A1 (n_5834), .B0 (n_5716), .Y (n_5752));
OAI21X1 g55834(.A0 (n_4322), .A1 (n_5750), .B0 (n_5721), .Y (n_5751));
DFFSRX1 WX10859_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5714), .Q (), .QN (WX10859));
DFFSRX1 WX1808_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5713), .Q (), .QN (WX1808));
OAI21X1 g56018(.A0 (n_4353), .A1 (n_5393), .B0 (n_5724), .Y (n_5749));
MX2X1 g56907(.A (n_5744), .B (WX523), .S0 (n_10735), .Y (n_5748));
NOR2X1 g56059(.A (WX6982), .B (n_5838), .Y (n_5747));
NOR2X1 g56931(.A (n_1425), .B (n_5744), .Y (n_5745));
OR2X1 g56939(.A (n_5744), .B (n_5990), .Y (n_5743));
NOR2X1 g56094(.A (WX8275), .B (n_3188), .Y (n_5742));
NOR2X1 g56098(.A (WX8275), .B (n_5500), .Y (n_9814));
NOR2X1 g55857(.A (WX3103), .B (n_5479), .Y (n_8538));
OAI21X1 g55957(.A0 (n_4247), .A1 (n_5841), .B0 (n_5708), .Y (n_5738));
NOR2X1 g56159(.A (WX9568), .B (n_3188), .Y (n_5737));
NOR2X1 g56161(.A (WX9568), .B (n_5427), .Y (n_6685));
NOR2X1 g55880(.A (WX3103), .B (n_1648), .Y (n_5735));
NOR2X1 g55993(.A (WX5689), .B (n_5712), .Y (n_5733));
NOR2X1 g55994(.A (WX5689), .B (n_5838), .Y (n_5732));
OAI21X1 g56724(.A0 (n_4450), .A1 (n_5729), .B0 (n_5707), .Y (n_5731));
OAI21X1 g56728(.A0 (n_3824), .A1 (n_5729), .B0 (n_5705), .Y (n_5730));
NAND2X1 g56882(.A (n_6575), .B (n_8334), .Y (n_5728));
INVX1 g56908(.A (DATA_9_11), .Y (n_5727));
NOR2X1 g56057(.A (WX6982), .B (n_1648), .Y (n_5725));
OAI21X1 g56060(.A0 (n_4405), .A1 (n_6686), .B0 (n_4860), .Y (n_5724));
OAI21X1 g56099(.A0 (n_5689), .A1 (n_9407), .B0 (n_5722), .Y (n_5723));
OAI21X1 g55859(.A0 (n_4449), .A1 (n_9815), .B0 (n_5566), .Y (n_5721));
OAI21X1 g56162(.A0 (n_5687), .A1 (n_9409), .B0 (n_4947), .Y (n_5720));
NOR2X1 g55986(.A (WX4398), .B (n_3188), .Y (n_5719));
NOR2X1 g55990(.A (WX4398), .B (n_5662), .Y (n_15856));
OAI21X1 g55995(.A0 (n_4248), .A1 (n_8539), .B0 (n_4860), .Y (n_5716));
NOR2X1 g56745(.A (WX10861), .B (n_1648), .Y (n_5714));
NOR2X1 g56746(.A (WX1810), .B (n_5712), .Y (n_5713));
NOR2X1 g56756(.A (WX1810), .B (n_5838), .Y (n_5711));
DFFSRX1 WX3267_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5700), .Q (WX3267), .QN ());
DFFSRX1 WX5853_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5699), .Q (WX5853), .QN ());
DFFSRX1 WX7146_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5703), .Q (WX7146), .QN ());
DFFSRX1 WX8439_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5702), .Q (WX8439), .QN ());
DFFSRX1 WX9732_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5701), .Q (WX9732), .QN ());
DFFSRX1 WX689_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6581), .Q (WX689), .QN ());
OAI21X1 g56909(.A0 (n_5695), .A1 (n_5709), .B0 (n_4027), .Y(DATA_9_11));
DFFSRX1 WX6982_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5693), .Q (), .QN (WX6982));
INVX1 g56952(.A (WX523), .Y (n_5744));
DFFSRX1 WX8275_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5690), .Q (), .QN (WX8275));
DFFSRX1 WX9568_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5688), .Q (), .QN (WX9568));
OAI21X1 g55991(.A0 (n_5660), .A1 (n_9411), .B0 (n_4947), .Y (n_5708));
DFFSRX1 WX3103_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5694), .Q (), .QN (WX3103));
DFFSRX1 WX5689_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5682), .Q (), .QN (WX5689));
OAI21X1 g56757(.A0 (n_5664), .A1 (n_4162), .B0 (n_5706), .Y (n_5707));
OAI21X1 g56761(.A0 (n_4523), .A1 (n_7504), .B0 (n_5619), .Y (n_5705));
DFFSRX1 WX4562_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5686), .Q (WX4562), .QN ());
DFFSRX1 WX11025_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6467), .Q (WX11025), .QN ());
DFFSRX1 WX1974_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5685), .Q (WX1974), .QN ());
OAI21X1 g56906(.A0 (n_5676), .A1 (n_5889), .B0 (n_5608), .Y (n_8334));
DFFSRX1 WX523_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5674), .Q (WX523), .QN ());
OAI21X1 g56077(.A0 (n_4121), .A1 (n_5235), .B0 (n_5670), .Y (n_5703));
OAI21X1 g56131(.A0 (n_4575), .A1 (n_5830), .B0 (n_5669), .Y (n_5702));
OAI21X1 g56191(.A0 (n_4269), .A1 (n_5834), .B0 (n_5667), .Y (n_5701));
DFFSRX1 WX4398_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5661), .Q (), .QN (WX4398));
OAI21X1 g55894(.A0 (n_4620), .A1 (n_5439), .B0 (n_5678), .Y (n_5700));
OAI21X1 g56017(.A0 (n_4404), .A1 (n_6106), .B0 (n_5658), .Y (n_5699));
DFFSRX1 WX10861_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5666), .Q (), .QN (WX10861));
DFFSRX1 WX1810_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5665), .Q (), .QN (WX1810));
NOR2X1 g55918(.A (WX3105), .B (n_5427), .Y (n_9815));
MX2X1 g56966(.A (n_5672), .B (WX525), .S0 (n_4026), .Y (n_5695));
NOR2X1 g55940(.A (WX3105), .B (n_5712), .Y (n_5694));
NOR2X1 g56116(.A (WX6984), .B (n_2851), .Y (n_5693));
NOR2X1 g56118(.A (WX6984), .B (n_5838), .Y (n_6686));
NOR2X1 g56153(.A (WX8277), .B (n_3690), .Y (n_5690));
NOR2X1 g56157(.A (WX8277), .B (n_5838), .Y (n_5689));
NOR2X1 g56218(.A (WX9570), .B (n_5712), .Y (n_5688));
NOR2X1 g56220(.A (WX9570), .B (n_5811), .Y (n_5687));
OAI21X1 g56016(.A0 (n_4245), .A1 (n_5535), .B0 (n_5654), .Y (n_5686));
OAI21X1 g56783(.A0 (n_4448), .A1 (n_5535), .B0 (n_5657), .Y (n_5685));
NOR2X1 g56052(.A (WX5691), .B (n_1648), .Y (n_5682));
NOR2X1 g56053(.A (WX5691), .B (n_5427), .Y (n_8539));
OAI21X1 g55919(.A0 (n_5638), .A1 (n_4447), .B0 (n_5460), .Y (n_5678));
INVX1 g56967(.A (DATA_9_10), .Y (n_5676));
NOR2X1 g56989(.A (n_5181), .B (n_5672), .Y (n_5674));
OR2X1 g56997(.A (n_5672), .B (n_5990), .Y (n_5671));
OAI21X1 g56119(.A0 (n_4403), .A1 (n_9816), .B0 (n_4947), .Y (n_5670));
OAI21X1 g56158(.A0 (n_15857), .A1 (n_15858), .B0 (n_7087), .Y(n_5669));
OAI21X1 g56221(.A0 (n_4574), .A1 (n_6687), .B0 (n_5460), .Y (n_5667));
NOR2X1 g56804(.A (WX10863), .B (n_1425), .Y (n_5666));
NOR2X1 g56805(.A (WX1812), .B (n_5712), .Y (n_5665));
NOR2X1 g56814(.A (WX1812), .B (n_5811), .Y (n_5664));
DFFSRX1 WX3269_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5651), .Q (WX3269), .QN ());
DFFSRX1 WX5855_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5652), .Q (WX5855), .QN ());
DFFSRX1 WX8441_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5648), .Q (WX8441), .QN ());
DFFSRX1 WX7148_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5650), .Q (WX7148), .QN ());
DFFSRX1 WX9734_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5646), .Q (WX9734), .QN ());
NOR2X1 g56818(.A (WX10863), .B (n_5662), .Y (n_7504));
NOR2X1 g56043(.A (WX4400), .B (n_2620), .Y (n_5661));
NOR2X1 g56049(.A (WX4400), .B (n_5811), .Y (n_5660));
OAI21X1 g56054(.A0 (n_5642), .A1 (n_11608), .B0 (n_3183), .Y(n_5658));
DFFSRX1 WX5691_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5643), .Q (), .QN (WX5691));
OAI21X1 g56968(.A0 (n_5628), .A1 (n_6091), .B0 (n_4021), .Y(DATA_9_10));
DFFSRX1 WX3105_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5634), .Q (), .QN (WX3105));
DFFSRX1 WX6984_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5641), .Q (), .QN (WX6984));
DFFSRX1 WX8277_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5637), .Q (), .QN (WX8277));
DFFSRX1 WX9570_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5633), .Q (), .QN (WX9570));
DFFSRX1 WX4564_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5644), .Q (WX4564), .QN ());
OAI21X1 g56816(.A0 (n_5616), .A1 (n_4160), .B0 (n_6497), .Y (n_5657));
DFFSRX1 WX11027_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5629), .Q (WX11027), .QN ());
DFFSRX1 WX1976_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5631), .Q (WX1976), .QN ());
DFFSRX1 WX691_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6541), .Q (WX691), .QN ());
OAI21X1 g56050(.A0 (n_4316), .A1 (n_8547), .B0 (n_6497), .Y (n_5654));
DFFSRX1 WX4400_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5627), .Q (), .QN (WX4400));
OAI21X1 g56076(.A0 (n_4402), .A1 (n_5254), .B0 (n_5625), .Y (n_5652));
INVX1 g57013(.A (WX525), .Y (n_5672));
OAI21X1 g55953(.A0 (n_4317), .A1 (n_5649), .B0 (n_5622), .Y (n_5651));
OAI21X1 g56136(.A0 (n_4349), .A1 (n_5649), .B0 (n_5623), .Y (n_5650));
OAI21X1 g56190(.A0 (n_4299), .A1 (n_5841), .B0 (n_5621), .Y (n_5648));
OAI21X1 g56250(.A0 (n_4267), .A1 (n_5439), .B0 (n_5620), .Y (n_5646));
DFFSRX1 WX10863_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5618), .Q (), .QN (WX10863));
DFFSRX1 WX1812_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5617), .Q (), .QN (WX1812));
OAI21X1 g56075(.A0 (n_4472), .A1 (n_5493), .B0 (n_5606), .Y (n_5644));
DFFSRX1 WX525_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5610), .Q (WX525), .QN ());
NOR2X1 g56111(.A (WX5693), .B (n_3188), .Y (n_5643));
NOR2X1 g56112(.A (WX5693), .B (n_5662), .Y (n_5642));
NOR2X1 g56175(.A (WX6986), .B (n_1648), .Y (n_5641));
NOR2X1 g56177(.A (WX6986), .B (n_5500), .Y (n_9816));
NOR2X1 g55977(.A (WX3107), .B (n_5811), .Y (n_5638));
NOR2X1 g56212(.A (WX8279), .B (n_1425), .Y (n_5637));
NOR2X1 g56216(.A (WX8279), .B (n_5811), .Y (n_15858));
NOR2X1 g55999(.A (WX3107), .B (n_3690), .Y (n_5634));
NOR2X1 g56277(.A (WX9572), .B (n_5181), .Y (n_5633));
NOR2X1 g56279(.A (WX9572), .B (n_4882), .Y (n_6687));
DFFSRX1 WX3235_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5605), .Q (WX3235), .QN ());
OAI21X1 g56843(.A0 (n_4229), .A1 (n_5630), .B0 (n_5604), .Y (n_5631));
OAI21X1 g56846(.A0 (n_3821), .A1 (n_5630), .B0 (n_5603), .Y (n_5629));
MX2X1 g57025(.A (n_5609), .B (WX527), .S0 (n_10739), .Y (n_5628));
NOR2X1 g56101(.A (WX4402), .B (n_1425), .Y (n_5627));
NOR2X1 g56108(.A (WX4402), .B (n_5052), .Y (n_8547));
OAI21X1 g56113(.A0 (n_4244), .A1 (n_8540), .B0 (n_5722), .Y (n_5625));
OAI21X1 g56178(.A0 (n_4401), .A1 (n_6683), .B0 (n_5619), .Y (n_5623));
OAI21X1 g55979(.A0 (n_4228), .A1 (n_9817), .B0 (n_4947), .Y (n_5622));
OAI21X1 g56217(.A0 (n_4348), .A1 (n_6688), .B0 (n_5566), .Y (n_5621));
OAI21X1 g56280(.A0 (n_4298), .A1 (n_9818), .B0 (n_5619), .Y (n_5620));
DFFSRX1 WX3271_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5597), .Q (WX3271), .QN ());
DFFSRX1 WX5857_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5601), .Q (WX5857), .QN ());
DFFSRX1 WX7150_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5599), .Q (WX7150), .QN ());
DFFSRX1 WX8443_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5596), .Q (WX8443), .QN ());
DFFSRX1 WX9736_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5595), .Q (WX9736), .QN ());
NOR2X1 g56863(.A (WX10865), .B (n_5712), .Y (n_5618));
NOR2X1 g56864(.A (WX1814), .B (n_3188), .Y (n_5617));
NOR2X1 g56874(.A (WX1814), .B (n_5052), .Y (n_5616));
INVX1 g57026(.A (DATA_9_9), .Y (n_5612));
NOR2X1 g57048(.A (n_1425), .B (n_5609), .Y (n_5610));
OR2X1 g57056(.A (n_5609), .B (n_4882), .Y (n_5608));
OAI21X1 g56109(.A0 (n_5568), .A1 (n_4314), .B0 (n_6479), .Y (n_5606));
DFFSRX1 WX5693_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5591), .Q (), .QN (WX5693));
DFFSRX1 WX6986_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5588), .Q (), .QN (WX6986));
DFFSRX1 WX8279_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5584), .Q (), .QN (WX8279));
DFFSRX1 WX3107_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5594), .Q (), .QN (WX3107));
DFFSRX1 WX4566_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5592), .Q (WX4566), .QN ());
DFFSRX1 WX11029_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5577), .Q (WX11029), .QN ());
DFFSRX1 WX1978_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5579), .Q (WX1978), .QN ());
DFFSRX1 WX9572_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5578), .Q (), .QN (WX9572));
OAI21X1 g56844(.A0 (n_4359), .A1 (n_5630), .B0 (n_5580), .Y (n_5605));
OAI21X1 g56877(.A0 (n_5573), .A1 (n_4158), .B0 (n_5460), .Y (n_5604));
OAI21X1 g56879(.A0 (n_4266), .A1 (n_7506), .B0 (n_4860), .Y (n_5603));
OAI21X1 g57027(.A0 (n_5554), .A1 (n_5843), .B0 (n_4019), .Y(DATA_9_9));
DFFSRX1 WX4402_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5569), .Q (), .QN (WX4402));
OAI21X1 g56135(.A0 (n_4400), .A1 (n_5600), .B0 (n_5567), .Y (n_5601));
OAI21X1 g56195(.A0 (n_4119), .A1 (n_5598), .B0 (n_5565), .Y (n_5599));
OAI21X1 g56012(.A0 (n_4315), .A1 (n_5841), .B0 (n_5563), .Y (n_5597));
OAI21X1 g56249(.A0 (n_4573), .A1 (n_5841), .B0 (n_5564), .Y (n_5596));
DFFSRX1 WX693_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6589), .Q (WX693), .QN ());
OAI21X1 g56309(.A0 (n_4518), .A1 (n_4803), .B0 (n_5562), .Y (n_5595));
DFFSRX1 WX10865_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5560), .Q (), .QN (WX10865));
DFFSRX1 WX1814_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5558), .Q (), .QN (WX1814));
NOR2X1 g56058(.A (WX3109), .B (n_1648), .Y (n_5594));
INVX1 g57072(.A (WX527), .Y (n_5609));
OAI21X1 g56134(.A0 (n_4243), .A1 (n_5600), .B0 (n_5553), .Y (n_5592));
NOR2X1 g56170(.A (WX5695), .B (n_1648), .Y (n_5591));
NOR2X1 g56171(.A (WX5695), .B (n_5479), .Y (n_8540));
NOR2X1 g56234(.A (WX6988), .B (n_1648), .Y (n_5588));
NOR2X1 g56236(.A (WX6988), .B (n_5500), .Y (n_6683));
NOR2X1 g56271(.A (WX8281), .B (n_5712), .Y (n_5584));
NOR2X1 g56275(.A (WX8281), .B (n_5427), .Y (n_6688));
DFFSRX1 WX4528_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5551), .Q (WX4528), .QN ());
DFFSRX1 WX3237_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5550), .Q (WX3237), .QN ());
NOR2X1 g56037(.A (WX3109), .B (n_5479), .Y (n_9817));
OAI21X1 g56886(.A0 (n_5547), .A1 (n_4282), .B0 (n_4947), .Y (n_5580));
OAI21X1 g56901(.A0 (n_4227), .A1 (n_5535), .B0 (n_5557), .Y (n_5579));
NOR2X1 g56336(.A (WX9574), .B (n_1648), .Y (n_5578));
OAI21X1 g56905(.A0 (n_3817), .A1 (n_5576), .B0 (n_5555), .Y (n_5577));
NOR2X1 g56338(.A (WX9574), .B (n_5427), .Y (n_9818));
NOR2X1 g56935(.A (WX1816), .B (n_5479), .Y (n_5573));
NOR2X1 g56937(.A (WX10867), .B (n_5479), .Y (n_7506));
DFFSRX1 WX527_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5541), .Q (WX527), .QN ());
NOR2X1 g56160(.A (WX4404), .B (n_1425), .Y (n_5569));
NOR2X1 g56167(.A (WX4404), .B (n_5662), .Y (n_5568));
OAI21X1 g56172(.A0 (n_5518), .A1 (n_9427), .B0 (n_5566), .Y (n_5567));
OAI21X1 g56237(.A0 (n_4399), .A1 (n_9819), .B0 (n_5275), .Y (n_5565));
OAI21X1 g56276(.A0 (n_5513), .A1 (n_11614), .B0 (n_5619), .Y(n_5564));
DFFSRX1 WX3273_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5546), .Q (WX3273), .QN ());
DFFSRX1 WX5859_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5537), .Q (WX5859), .QN ());
DFFSRX1 WX7152_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5536), .Q (WX7152), .QN ());
DFFSRX1 WX8445_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5534), .Q (WX8445), .QN ());
DFFSRX1 WX9738_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5545), .Q (WX9738), .QN ());
DFFSRX1 WX3073_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5548), .Q (), .QN (WX3073));
OAI21X1 g56038(.A0 (n_5525), .A1 (n_11612), .B0 (n_5566), .Y(n_5563));
OAI21X1 g56339(.A0 (n_4572), .A1 (n_9820), .B0 (n_4947), .Y (n_5562));
NOR2X1 g56921(.A (WX10867), .B (n_3690), .Y (n_5560));
NOR2X1 g56922(.A (WX1816), .B (n_2605), .Y (n_5558));
OAI21X1 g56936(.A0 (n_5509), .A1 (n_4156), .B0 (n_5556), .Y (n_5557));
OAI21X1 g56938(.A0 (n_4517), .A1 (n_7505), .B0 (n_4860), .Y (n_5555));
DFFSRX1 WX9574_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5528), .Q (), .QN (WX9574));
DFFSRX1 WX3109_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5523), .Q (), .QN (WX3109));
MX2X1 g57084(.A (n_5540), .B (WX529), .S0 (n_4018), .Y (n_5554));
OAI21X1 g56168(.A0 (n_4310), .A1 (n_8548), .B0 (n_5460), .Y (n_5553));
DFFSRX1 WX5695_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5519), .Q (), .QN (WX5695));
DFFSRX1 WX6988_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5517), .Q (), .QN (WX6988));
DFFSRX1 WX4568_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5521), .Q (WX4568), .QN ());
DFFSRX1 WX11031_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5529), .Q (WX11031), .QN ());
DFFSRX1 WX1980_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5530), .Q (WX1980), .QN ());
DFFSRX1 WX8281_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5514), .Q (), .QN (WX8281));
OAI21X1 g56898(.A0 (n_4520), .A1 (n_5334), .B0 (n_5533), .Y (n_5551));
OAI21X1 g56903(.A0 (n_4355), .A1 (n_5549), .B0 (n_5532), .Y (n_5550));
NOR2X1 g56943(.A (WX3075), .B (n_5181), .Y (n_5548));
NOR2X1 g56944(.A (WX3075), .B (n_5427), .Y (n_5547));
DFFSRX1 WX10867_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5512), .Q (), .QN (WX10867));
DFFSRX1 WX1816_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5511), .Q (), .QN (WX1816));
OAI21X1 g56071(.A0 (n_4311), .A1 (n_5185), .B0 (n_5505), .Y (n_5546));
OAI21X1 g56368(.A0 (n_4516), .A1 (n_4866), .B0 (n_5507), .Y (n_5545));
INVX1 g57085(.A (DATA_9_8), .Y (n_5543));
NOR2X1 g57107(.A (n_1425), .B (n_5540), .Y (n_5541));
OR2X1 g57115(.A (n_5540), .B (n_3828), .Y (n_5539));
DFFSRX1 WX4404_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5503), .Q (), .QN (WX4404));
OAI21X1 g56194(.A0 (n_4220), .A1 (n_5490), .B0 (n_5499), .Y (n_5537));
OAI21X1 g56254(.A0 (n_4345), .A1 (n_5535), .B0 (n_5497), .Y (n_5536));
OAI21X1 g56308(.A0 (n_4293), .A1 (n_5845), .B0 (n_5496), .Y (n_5534));
OAI21X1 g56928(.A0 (n_5480), .A1 (n_4358), .B0 (n_5722), .Y (n_5533));
OAI21X1 g56945(.A0 (n_5477), .A1 (n_4557), .B0 (n_3183), .Y (n_5532));
OAI21X1 g56960(.A0 (n_4425), .A1 (n_5535), .B0 (n_5489), .Y (n_5530));
OAI21X1 g56964(.A0 (n_3816), .A1 (n_5474), .B0 (n_5488), .Y (n_5529));
NOR2X1 g56395(.A (WX9576), .B (n_1648), .Y (n_5528));
NOR2X1 g56398(.A (WX9576), .B (n_5427), .Y (n_9820));
NOR2X1 g56096(.A (WX3111), .B (n_3218), .Y (n_5525));
OAI21X1 g57086(.A0 (n_5473), .A1 (n_5965), .B0 (n_4080), .Y(DATA_9_8));
NOR2X1 g56117(.A (WX3111), .B (n_5712), .Y (n_5523));
OAI21X1 g56193(.A0 (n_4469), .A1 (n_5235), .B0 (n_5485), .Y (n_5521));
NOR2X1 g56229(.A (WX5697), .B (n_1425), .Y (n_5519));
NOR2X1 g56230(.A (WX5697), .B (n_5500), .Y (n_5518));
NOR2X1 g56293(.A (WX6990), .B (n_2620), .Y (n_5517));
DFFSRX1 WX5821_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5492), .Q (WX5821), .QN ());
DFFSRX1 WX4530_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5494), .Q (WX4530), .QN ());
DFFSRX1 WX3239_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5491), .Q (WX3239), .QN ());
DFFSRX1 WX695_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5486), .Q (WX695), .QN ());
NOR2X1 g56295(.A (WX6990), .B (n_5500), .Y (n_9819));
NOR2X1 g56330(.A (WX8283), .B (n_5712), .Y (n_5514));
NOR2X1 g56334(.A (WX8283), .B (n_5500), .Y (n_5513));
DFFSRX1 WX3075_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5478), .Q (), .QN (WX3075));
NOR2X1 g56980(.A (WX10869), .B (n_2849), .Y (n_5512));
NOR2X1 g56981(.A (WX1818), .B (n_2849), .Y (n_5511));
NOR2X1 g56993(.A (WX1818), .B (n_5838), .Y (n_5509));
NOR2X1 g56995(.A (WX10869), .B (n_5662), .Y (n_7505));
OAI21X1 g56397(.A0 (n_4292), .A1 (n_8549), .B0 (n_5722), .Y (n_5507));
OAI21X1 g56097(.A0 (n_4424), .A1 (n_9821), .B0 (n_5722), .Y (n_5505));
INVX1 g57123(.A (WX529), .Y (n_5540));
NOR2X1 g56219(.A (WX4406), .B (n_2851), .Y (n_5503));
NOR2X1 g56226(.A (WX4406), .B (n_5500), .Y (n_8548));
OAI21X1 g56231(.A0 (n_5437), .A1 (n_11616), .B0 (n_4947), .Y(n_5499));
DFFSRX1 WX3275_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5472), .Q (WX3275), .QN ());
DFFSRX1 WX5861_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5471), .Q (WX5861), .QN ());
DFFSRX1 WX7154_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5469), .Q (WX7154), .QN ());
DFFSRX1 WX8447_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5483), .Q (WX8447), .QN ());
DFFSRX1 WX9740_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5475), .Q (WX9740), .QN ());
DFFSRX1 WX4366_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5481), .Q (), .QN (WX4366));
OAI21X1 g56296(.A0 (n_5465), .A1 (n_4219), .B0 (n_4947), .Y (n_5497));
OAI21X1 g56335(.A0 (n_5459), .A1 (n_9429), .B0 (n_5460), .Y (n_5496));
DFFSRX1 WX8283_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5462), .Q (), .QN (WX8283));
OAI21X1 g56957(.A0 (n_4508), .A1 (n_5493), .B0 (n_5464), .Y (n_5494));
OAI21X1 g56959(.A0 (n_4442), .A1 (n_5415), .B0 (n_5463), .Y (n_5492));
OAI21X1 g56962(.A0 (n_4351), .A1 (n_5490), .B0 (n_5461), .Y (n_5491));
OAI21X1 g56994(.A0 (n_5429), .A1 (n_4154), .B0 (n_5722), .Y (n_5489));
OAI21X1 g56996(.A0 (n_4515), .A1 (n_6678), .B0 (n_4860), .Y (n_5488));
DFFSRX1 WX9576_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5453), .Q (), .QN (WX9576));
NAND2X1 g57081(.A (n_5454), .B (n_4698), .Y (n_5486));
DFFSRX1 WX529_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5448), .Q (WX529), .QN ());
DFFSRX1 WX3111_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5442), .Q (), .QN (WX3111));
OAI21X1 g56227(.A0 (n_4308), .A1 (n_8550), .B0 (n_5556), .Y (n_5485));
DFFSRX1 WX5697_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5438), .Q (), .QN (WX5697));
DFFSRX1 WX4570_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5440), .Q (WX4570), .QN ());
DFFSRX1 WX11033_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5456), .Q (WX11033), .QN ());
DFFSRX1 WX1982_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5458), .Q (WX1982), .QN ());
DFFSRX1 WX6990_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5467), .Q (), .QN (WX6990));
OAI21X1 g56367(.A0 (n_4291), .A1 (n_5482), .B0 (n_5434), .Y (n_5483));
NOR2X1 g56983(.A (WX4368), .B (n_5181), .Y (n_5481));
NOR2X1 g56985(.A (WX4368), .B (n_5479), .Y (n_5480));
NOR2X1 g57002(.A (WX3077), .B (n_5181), .Y (n_5478));
NOR2X1 g57003(.A (WX3077), .B (n_5662), .Y (n_5477));
DFFSRX1 WX10869_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5432), .Q (), .QN (WX10869));
DFFSRX1 WX1818_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5430), .Q (), .QN (WX1818));
OAI21X1 g56427(.A0 (n_4514), .A1 (n_5474), .B0 (n_5426), .Y (n_5475));
MX2X1 g57143(.A (n_5446), .B (WX531), .S0 (n_4079), .Y (n_5473));
OAI21X1 g56130(.A0 (n_4309), .A1 (n_5105), .B0 (n_5425), .Y (n_5472));
DFFSRX1 WX4406_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5424), .Q (), .QN (WX4406));
OAI21X1 g56253(.A0 (n_4218), .A1 (n_4803), .B0 (n_5421), .Y (n_5471));
OAI21X1 g56313(.A0 (n_4117), .A1 (n_5468), .B0 (n_5436), .Y (n_5469));
NOR2X1 g56352(.A (WX6992), .B (n_2851), .Y (n_5467));
NOR2X1 g56354(.A (WX6992), .B (n_5052), .Y (n_5465));
OAI21X1 g56986(.A0 (n_4354), .A1 (n_6191), .B0 (n_5722), .Y (n_5464));
OAI21X1 g56992(.A0 (n_5403), .A1 (n_4519), .B0 (n_3183), .Y (n_5463));
NOR2X1 g56389(.A (WX8285), .B (n_1425), .Y (n_5462));
OAI21X1 g57004(.A0 (n_4555), .A1 (n_6673), .B0 (n_5460), .Y (n_5461));
NOR2X1 g56393(.A (WX8285), .B (n_5500), .Y (n_5459));
OAI21X1 g57019(.A0 (n_4418), .A1 (n_5415), .B0 (n_5414), .Y (n_5458));
OAI21X1 g57023(.A0 (n_3815), .A1 (n_5892), .B0 (n_5413), .Y (n_5456));
NAND2X1 g57117(.A (n_5411), .B (n_6615), .Y (n_5454));
NOR2X1 g56454(.A (WX9578), .B (n_5181), .Y (n_5453));
NOR2X1 g56456(.A (WX9578), .B (n_5427), .Y (n_8549));
INVX1 g57144(.A (DATA_9_7), .Y (n_5450));
NOR2X1 g57167(.A (n_1425), .B (n_5446), .Y (n_5448));
OR2X1 g57175(.A (n_5446), .B (n_4882), .Y (n_5445));
NOR2X1 g56155(.A (WX3113), .B (n_5500), .Y (n_9821));
NOR2X1 g56176(.A (WX3113), .B (n_5712), .Y (n_5442));
OAI21X1 g56252(.A0 (n_4466), .A1 (n_5439), .B0 (n_5410), .Y (n_5440));
NOR2X1 g56288(.A (WX5699), .B (n_1648), .Y (n_5438));
NOR2X1 g56289(.A (WX5699), .B (n_3218), .Y (n_5437));
DFFSRX1 WX5823_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5419), .Q (WX5823), .QN ());
DFFSRX1 WX4532_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5420), .Q (WX4532), .QN ());
DFFSRX1 WX7114_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5417), .Q (WX7114), .QN ());
DFFSRX1 WX3241_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5416), .Q (WX3241), .QN ());
OAI21X1 g56355(.A0 (n_5386), .A1 (n_11618), .B0 (n_5722), .Y(n_5436));
DFFSRX1 WX4368_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5407), .Q (), .QN (WX4368));
DFFSRX1 WX3077_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5401), .Q (), .QN (WX3077));
OAI21X1 g56394(.A0 (n_4116), .A1 (n_8551), .B0 (n_4860), .Y (n_5434));
NOR2X1 g57040(.A (WX10871), .B (n_3188), .Y (n_5432));
NOR2X1 g57041(.A (WX1820), .B (n_1648), .Y (n_5430));
NOR2X1 g57052(.A (WX1820), .B (n_5838), .Y (n_5429));
NOR2X1 g57054(.A (WX10871), .B (n_5427), .Y (n_6678));
OAI21X1 g56457(.A0 (n_4290), .A1 (n_8552), .B0 (n_5722), .Y (n_5426));
OAI21X1 g57145(.A0 (n_5377), .A1 (n_5965), .B0 (n_4077), .Y(DATA_9_7));
OAI21X1 g56156(.A0 (n_4417), .A1 (n_6689), .B0 (n_5722), .Y (n_5425));
NOR2X1 g56278(.A (WX4408), .B (n_5181), .Y (n_5424));
NOR2X1 g56284(.A (WX4408), .B (n_3218), .Y (n_8550));
OAI21X1 g56290(.A0 (n_4467), .A1 (n_6690), .B0 (n_4947), .Y (n_5421));
DFFSRX1 WX3277_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5395), .Q (WX3277), .QN ());
DFFSRX1 WX5863_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5394), .Q (WX5863), .QN ());
DFFSRX1 WX7156_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5409), .Q (WX7156), .QN ());
DFFSRX1 WX8449_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5398), .Q (WX8449), .QN ());
DFFSRX1 WX9742_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5396), .Q (WX9742), .QN ());
DFFSRX1 WX5659_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5404), .Q (), .QN (WX5659));
DFFSRX1 WX697_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5397), .Q (WX697), .QN ());
DFFSRX1 WX6992_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5388), .Q (), .QN (WX6992));
OAI21X1 g57017(.A0 (n_4502), .A1 (n_5841), .B0 (n_5390), .Y (n_5420));
OAI21X1 g57018(.A0 (n_4440), .A1 (n_5418), .B0 (n_5389), .Y (n_5419));
OAI21X1 g57020(.A0 (n_4381), .A1 (n_5439), .B0 (n_5385), .Y (n_5417));
OAI21X1 g57021(.A0 (n_4347), .A1 (n_5415), .B0 (n_5384), .Y (n_5416));
OAI21X1 g57053(.A0 (n_5365), .A1 (n_4152), .B0 (n_5556), .Y (n_5414));
OAI21X1 g57055(.A0 (n_4513), .A1 (n_6679), .B0 (n_4860), .Y (n_5413));
DFFSRX1 WX8285_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5380), .Q (), .QN (WX8285));
OAI21X1 g57142(.A0 (n_5360), .A1 (n_5889), .B0 (n_5256), .Y (n_5411));
DFFSRX1 WX9578_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5376), .Q (), .QN (WX9578));
INVX1 g57184(.A (WX531), .Y (n_5446));
DFFSRX1 WX3113_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5371), .Q (), .QN (WX3113));
DFFSRX1 WX11035_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6486), .Q (WX11035), .QN ());
OAI21X1 g56286(.A0 (n_15851), .A1 (n_15852), .B0 (n_5722), .Y(n_5410));
DFFSRX1 WX4572_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5370), .Q (WX4572), .QN ());
DFFSRX1 WX1984_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5382), .Q (WX1984), .QN ());
DFFSRX1 WX5699_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5392), .Q (), .QN (WX5699));
OAI21X1 g56372(.A0 (n_4341), .A1 (n_5105), .B0 (n_5368), .Y (n_5409));
NOR2X1 g57042(.A (WX4370), .B (n_1648), .Y (n_5407));
NOR2X1 g57045(.A (WX4370), .B (n_5662), .Y (n_6191));
NOR2X1 g57049(.A (WX5661), .B (n_1648), .Y (n_5404));
NOR2X1 g57050(.A (WX5661), .B (n_5838), .Y (n_5403));
NOR2X1 g57061(.A (WX3079), .B (n_5181), .Y (n_5401));
NOR2X1 g57062(.A (WX3079), .B (n_5479), .Y (n_6673));
DFFSRX1 WX10871_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5367), .Q (), .QN (WX10871));
DFFSRX1 WX1820_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5366), .Q (), .QN (WX1820));
OAI21X1 g56426(.A0 (n_4289), .A1 (n_5105), .B0 (n_5362), .Y (n_5398));
NAND2X2 g57140(.A (n_5361), .B (n_4695), .Y (n_5397));
DFFSRX1 WX531_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5358), .Q (WX531), .QN ());
OAI21X1 g56486(.A0 (n_4512), .A1 (n_5649), .B0 (n_5354), .Y (n_5396));
OAI21X1 g56189(.A0 (n_4307), .A1 (n_5841), .B0 (n_5353), .Y (n_5395));
DFFSRX1 WX4408_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5352), .Q (), .QN (WX4408));
OAI21X1 g56312(.A0 (n_4396), .A1 (n_5393), .B0 (n_5369), .Y (n_5394));
NOR2X1 g56347(.A (WX5701), .B (n_1425), .Y (n_5392));
NOR2X1 g56348(.A (WX5701), .B (n_5479), .Y (n_6690));
OAI21X1 g57047(.A0 (n_5331), .A1 (n_4350), .B0 (n_5556), .Y (n_5390));
OAI21X1 g57051(.A0 (n_4507), .A1 (n_6666), .B0 (n_4860), .Y (n_5389));
NOR2X1 g56411(.A (WX6994), .B (n_5181), .Y (n_5388));
NOR2X1 g56413(.A (WX6994), .B (n_5838), .Y (n_5386));
OAI21X1 g57060(.A0 (n_4441), .A1 (n_6192), .B0 (n_5722), .Y (n_5385));
OAI21X1 g57063(.A0 (n_4553), .A1 (n_6193), .B0 (n_4860), .Y (n_5384));
OAI21X1 g57078(.A0 (n_4225), .A1 (n_5918), .B0 (n_5342), .Y (n_5382));
NOR2X1 g56448(.A (WX8287), .B (n_1425), .Y (n_5380));
NOR2X1 g56452(.A (WX8287), .B (n_5838), .Y (n_8551));
MX2X1 g57204(.A (n_5356), .B (WX533), .S0 (n_4076), .Y (n_5377));
NOR2X1 g56513(.A (WX9580), .B (n_1648), .Y (n_5376));
NOR2X1 g56515(.A (WX9580), .B (n_5427), .Y (n_8552));
DFFSRX1 WX5825_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5347), .Q (WX5825), .QN ());
NOR2X1 g56214(.A (WX3115), .B (n_5811), .Y (n_6689));
NOR2X1 g56235(.A (WX3115), .B (n_5181), .Y (n_5371));
DFFSRX1 WX8407_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5350), .Q (WX8407), .QN ());
DFFSRX1 WX4534_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5348), .Q (WX4534), .QN ());
DFFSRX1 WX7116_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5345), .Q (WX7116), .QN ());
DFFSRX1 WX3243_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5343), .Q (WX3243), .QN ());
OAI21X1 g56311(.A0 (n_4462), .A1 (n_5393), .B0 (n_5338), .Y (n_5370));
OAI21X1 g56349(.A0 (n_4465), .A1 (n_6691), .B0 (n_5460), .Y (n_5369));
OAI21X1 g56414(.A0 (n_4395), .A1 (n_6692), .B0 (n_5722), .Y (n_5368));
DFFSRX1 WX4370_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5333), .Q (), .QN (WX4370));
DFFSRX1 WX5661_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5330), .Q (), .QN (WX5661));
DFFSRX1 WX3079_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5325), .Q (), .QN (WX3079));
NOR2X1 g57099(.A (WX10873), .B (n_1648), .Y (n_5367));
NOR2X1 g57100(.A (WX1822), .B (n_1425), .Y (n_5366));
NOR2X1 g57111(.A (WX1822), .B (n_5662), .Y (n_5365));
NOR2X1 g57113(.A (WX10873), .B (n_5662), .Y (n_6679));
OAI21X1 g56453(.A0 (n_4340), .A1 (n_9822), .B0 (n_5566), .Y (n_5362));
NAND2X1 g57177(.A (n_6575), .B (n_8335), .Y (n_5361));
INVX1 g57205(.A (DATA_9_6), .Y (n_5360));
NOR2X1 g57227(.A (n_1425), .B (n_5356), .Y (n_5358));
OR2X1 g57236(.A (n_5356), .B (n_5968), .Y (n_5355));
OAI21X1 g56516(.A0 (n_4288), .A1 (n_9823), .B0 (n_5566), .Y (n_5354));
OAI21X1 g56215(.A0 (n_5294), .A1 (n_4224), .B0 (n_4860), .Y (n_5353));
DFFSRX1 WX3279_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5319), .Q (WX3279), .QN ());
DFFSRX1 WX5865_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5336), .Q (WX5865), .QN ());
DFFSRX1 WX7158_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5335), .Q (WX7158), .QN ());
DFFSRX1 WX8451_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5323), .Q (WX8451), .QN ());
DFFSRX1 WX9744_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5321), .Q (WX9744), .QN ());
DFFSRX1 WX6952_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5328), .Q (), .QN (WX6952));
NOR2X1 g56337(.A (WX4410), .B (n_5712), .Y (n_5352));
NOR2X1 g56343(.A (WX4410), .B (n_5662), .Y (n_15852));
DFFSRX1 WX5701_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5316), .Q (), .QN (WX5701));
DFFSRX1 WX6994_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5304), .Q (), .QN (WX6994));
OAI21X1 g57074(.A0 (n_4616), .A1 (n_5439), .B0 (n_5314), .Y (n_5350));
OAI21X1 g57076(.A0 (n_4500), .A1 (n_5892), .B0 (n_5313), .Y (n_5348));
OAI21X1 g57077(.A0 (n_4437), .A1 (n_5841), .B0 (n_5311), .Y (n_5347));
OAI21X1 g57079(.A0 (n_4379), .A1 (n_5879), .B0 (n_5310), .Y (n_5345));
OAI21X1 g57080(.A0 (n_4343), .A1 (n_5320), .B0 (n_5309), .Y (n_5343));
OAI21X1 g57112(.A0 (n_5285), .A1 (n_4149), .B0 (n_5566), .Y (n_5342));
DFFSRX1 WX8287_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5300), .Q (), .QN (WX8287));
OAI21X1 g57206(.A0 (n_5279), .A1 (n_5709), .B0 (n_4068), .Y(DATA_9_6));
DFFSRX1 WX9580_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5297), .Q (), .QN (WX9580));
DFFSRX1 WX3115_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5293), .Q (), .QN (WX3115));
DFFSRX1 WX4574_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5318), .Q (WX4574), .QN ());
DFFSRX1 WX11037_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5305), .Q (WX11037), .QN ());
DFFSRX1 WX1986_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5307), .Q (WX1986), .QN ());
DFFSRX1 WX699_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6549), .Q (WX699), .QN ());
OAI21X1 g56344(.A0 (n_4304), .A1 (n_8541), .B0 (n_4947), .Y (n_5338));
DFFSRX1 WX4410_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5291), .Q (), .QN (WX4410));
OAI21X1 g56371(.A0 (n_4654), .A1 (n_5317), .B0 (n_5289), .Y (n_5336));
OAI21X1 g56431(.A0 (n_4115), .A1 (n_5334), .B0 (n_5282), .Y (n_5335));
NOR2X1 g57101(.A (WX4372), .B (n_5181), .Y (n_5333));
NOR2X1 g57105(.A (WX4372), .B (n_5479), .Y (n_5331));
NOR2X1 g57108(.A (WX5663), .B (n_1648), .Y (n_5330));
NOR2X1 g57109(.A (WX5663), .B (n_5662), .Y (n_6666));
NOR2X1 g57116(.A (WX6954), .B (n_5712), .Y (n_5328));
NOR2X1 g57118(.A (WX6954), .B (n_5662), .Y (n_6192));
NOR2X1 g57120(.A (WX3081), .B (n_1648), .Y (n_5325));
NOR2X1 g57121(.A (WX3081), .B (n_5811), .Y (n_6193));
DFFSRX1 WX10873_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5288), .Q (), .QN (WX10873));
DFFSRX1 WX1822_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5287), .Q (), .QN (WX1822));
OAI21X1 g56485(.A0 (n_4287), .A1 (n_5105), .B0 (n_5281), .Y (n_5323));
OAI21X1 g57203(.A0 (n_5261), .A1 (n_5889), .B0 (n_5160), .Y (n_8335));
INVX1 g57247(.A (WX533), .Y (n_5356));
OAI21X1 g56545(.A0 (n_4510), .A1 (n_5320), .B0 (n_5278), .Y (n_5321));
OAI21X1 g56248(.A0 (n_4305), .A1 (n_5535), .B0 (n_5276), .Y (n_5319));
OAI21X1 g56370(.A0 (n_4239), .A1 (n_5317), .B0 (n_5274), .Y (n_5318));
DFFSRX1 WX9700_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5272), .Q (WX9700), .QN ());
NOR2X1 g56406(.A (WX5703), .B (n_2620), .Y (n_5316));
NOR2X1 g56407(.A (WX5703), .B (n_5500), .Y (n_6691));
OAI21X1 g57098(.A0 (n_5252), .A1 (n_4380), .B0 (n_4860), .Y (n_5314));
OAI21X1 g57106(.A0 (n_5250), .A1 (n_4346), .B0 (n_5566), .Y (n_5313));
OAI21X1 g57110(.A0 (n_4501), .A1 (n_6221), .B0 (n_4860), .Y (n_5311));
OAI21X1 g57119(.A0 (n_4438), .A1 (n_6194), .B0 (n_5460), .Y (n_5310));
OAI21X1 g57122(.A0 (n_4521), .A1 (n_6667), .B0 (n_5722), .Y (n_5309));
OAI21X1 g57137(.A0 (n_4223), .A1 (n_5928), .B0 (n_5264), .Y (n_5307));
OAI21X1 g57141(.A0 (n_3813), .A1 (n_5886), .B0 (n_5263), .Y (n_5305));
NOR2X1 g56470(.A (WX6996), .B (n_1648), .Y (n_5304));
NOR2X1 g56472(.A (WX6996), .B (n_5811), .Y (n_6692));
NOR2X1 g56506(.A (WX8289), .B (n_1425), .Y (n_5300));
DFFSRX1 WX533_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5259), .Q (WX533), .QN ());
NOR2X1 g56511(.A (WX8289), .B (n_5838), .Y (n_9822));
NOR2X1 g56573(.A (WX9582), .B (n_1648), .Y (n_5297));
NOR2X1 g56575(.A (WX9582), .B (n_5822), .Y (n_9823));
NOR2X1 g56273(.A (WX3117), .B (n_5811), .Y (n_5294));
NOR2X1 g56294(.A (WX3117), .B (n_5181), .Y (n_5293));
DFFSRX1 WX8409_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5273), .Q (WX8409), .QN ());
DFFSRX1 WX4536_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5271), .Q (WX4536), .QN ());
DFFSRX1 WX5827_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5269), .Q (WX5827), .QN ());
DFFSRX1 WX7118_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5267), .Q (WX7118), .QN ());
DFFSRX1 WX3245_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5265), .Q (WX3245), .QN ());
NOR2X1 g56396(.A (WX4412), .B (n_3690), .Y (n_5291));
NOR2X1 g56401(.A (WX4412), .B (n_5427), .Y (n_8541));
OAI21X1 g56408(.A0 (n_4461), .A1 (n_6693), .B0 (n_4860), .Y (n_5289));
DFFSRX1 WX4372_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5251), .Q (), .QN (WX4372));
DFFSRX1 WX5663_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5249), .Q (), .QN (WX5663));
DFFSRX1 WX6954_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5247), .Q (), .QN (WX6954));
DFFSRX1 WX3081_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5245), .Q (), .QN (WX3081));
NOR2X1 g57159(.A (WX10875), .B (n_2620), .Y (n_5288));
NOR2X1 g57160(.A (WX1824), .B (n_2620), .Y (n_5287));
NOR2X1 g57171(.A (WX1824), .B (n_5838), .Y (n_5285));
OAI21X1 g56473(.A0 (n_4653), .A1 (n_9824), .B0 (n_5722), .Y (n_5282));
OAI21X1 g56512(.A0 (n_4114), .A1 (n_8542), .B0 (n_3183), .Y (n_5281));
MX2X1 g57265(.A (n_5257), .B (WX535), .S0 (n_6601), .Y (n_5279));
OAI21X1 g56576(.A0 (n_4286), .A1 (n_8553), .B0 (n_5460), .Y (n_5278));
OAI21X1 g56274(.A0 (n_5214), .A1 (n_4222), .B0 (n_5275), .Y (n_5276));
DFFSRX1 WX3281_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5238), .Q (WX3281), .QN ());
DFFSRX1 WX5867_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5255), .Q (WX5867), .QN ());
DFFSRX1 WX7160_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5243), .Q (WX7160), .QN ());
DFFSRX1 WX8453_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5241), .Q (WX8453), .QN ());
DFFSRX1 WX9746_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5240), .Q (WX9746), .QN ());
DFFSRX1 WX8245_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5253), .Q (), .QN (WX8245));
OAI21X1 g56402(.A0 (n_5212), .A1 (n_9413), .B0 (n_5566), .Y (n_5274));
DFFSRX1 WX5703_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5233), .Q (), .QN (WX5703));
OAI21X1 g57133(.A0 (n_4613), .A1 (n_5239), .B0 (n_5234), .Y (n_5273));
OAI21X1 g57134(.A0 (n_4552), .A1 (n_5158), .B0 (n_5232), .Y (n_5272));
OAI21X1 g57135(.A0 (n_4498), .A1 (n_5535), .B0 (n_5230), .Y (n_5271));
OAI21X1 g57136(.A0 (n_4435), .A1 (n_5493), .B0 (n_5228), .Y (n_5269));
OAI21X1 g57138(.A0 (n_4377), .A1 (n_5535), .B0 (n_5227), .Y (n_5267));
OAI21X1 g57139(.A0 (n_4339), .A1 (n_5196), .B0 (n_5226), .Y (n_5265));
OAI21X1 g57172(.A0 (n_5207), .A1 (n_4147), .B0 (n_4947), .Y (n_5264));
OAI21X1 g57174(.A0 (n_4509), .A1 (n_6682), .B0 (n_5460), .Y (n_5263));
DFFSRX1 WX6996_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5222), .Q (), .QN (WX6996));
INVX1 g57266(.A (DATA_9_5), .Y (n_5261));
NOR2X1 g57293(.A (n_5181), .B (n_5257), .Y (n_5259));
DFFSRX1 WX8289_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5219), .Q (), .QN (WX8289));
OR2X1 g57302(.A (n_5257), .B (n_5968), .Y (n_5256));
DFFSRX1 WX9582_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5217), .Q (), .QN (WX9582));
DFFSRX1 WX4576_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5236), .Q (WX4576), .QN ());
DFFSRX1 WX1988_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5225), .Q (WX1988), .QN ());
DFFSRX1 WX3117_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5237), .Q (), .QN (WX3117));
DFFSRX1 WX11039_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5224), .Q (WX11039), .QN ());
DFFSRX1 WX4412_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5213), .Q (), .QN (WX4412));
OAI21X1 g56430(.A0 (n_4215), .A1 (n_5254), .B0 (n_5211), .Y (n_5255));
NOR2X1 g57156(.A (WX8247), .B (n_5712), .Y (n_5253));
NOR2X1 g57157(.A (WX8247), .B (n_5811), .Y (n_5252));
NOR2X1 g57162(.A (WX4374), .B (n_1425), .Y (n_5251));
NOR2X1 g57165(.A (WX4374), .B (n_5662), .Y (n_5250));
NOR2X1 g57168(.A (WX5665), .B (n_5712), .Y (n_5249));
NOR2X1 g57169(.A (WX5665), .B (n_5838), .Y (n_6221));
NOR2X1 g57176(.A (WX6956), .B (n_5181), .Y (n_5247));
NOR2X1 g57178(.A (WX6956), .B (n_5427), .Y (n_6194));
NOR2X1 g57180(.A (WX3083), .B (n_5181), .Y (n_5245));
NOR2X1 g57181(.A (WX3083), .B (n_5500), .Y (n_6667));
DFFSRX1 WX10875_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5210), .Q (), .QN (WX10875));
DFFSRX1 WX1824_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5208), .Q (), .QN (WX1824));
OAI21X1 g56490(.A0 (n_4113), .A1 (n_5183), .B0 (n_5203), .Y (n_5243));
OAI21X1 g57267(.A0 (n_5187), .A1 (n_5242), .B0 (n_4066), .Y(DATA_9_5));
OAI21X1 g56544(.A0 (n_4285), .A1 (n_5320), .B0 (n_5201), .Y (n_5241));
OAI21X1 g56605(.A0 (n_4506), .A1 (n_5239), .B0 (n_5200), .Y (n_5240));
DFFSRX1 WX701_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5204), .Q (WX701), .QN ());
OAI21X1 g56307(.A0 (n_4587), .A1 (n_5085), .B0 (n_5199), .Y (n_5238));
NOR2X1 g56353(.A (WX3119), .B (n_5712), .Y (n_5237));
OAI21X1 g56429(.A0 (n_4237), .A1 (n_5235), .B0 (n_5198), .Y (n_5236));
OAI21X1 g57158(.A0 (n_5180), .A1 (n_4378), .B0 (n_6479), .Y (n_5234));
NOR2X1 g56465(.A (WX5705), .B (n_5181), .Y (n_5233));
OAI21X1 g57164(.A0 (n_4614), .A1 (n_6222), .B0 (n_5722), .Y (n_5232));
NOR2X1 g56466(.A (WX5705), .B (n_5662), .Y (n_6693));
OAI21X1 g57166(.A0 (n_4342), .A1 (n_6223), .B0 (n_5566), .Y (n_5230));
OAI21X1 g57170(.A0 (n_4499), .A1 (n_6224), .B0 (n_4860), .Y (n_5228));
OAI21X1 g57179(.A0 (n_4436), .A1 (n_6674), .B0 (n_6479), .Y (n_5227));
OAI21X1 g57182(.A0 (n_4495), .A1 (n_6225), .B0 (n_4860), .Y (n_5226));
OAI21X1 g57197(.A0 (n_4398), .A1 (n_5493), .B0 (n_5190), .Y (n_5225));
OAI21X1 g57202(.A0 (n_3811), .A1 (n_5535), .B0 (n_5189), .Y (n_5224));
NOR2X1 g56529(.A (WX6998), .B (n_5712), .Y (n_5222));
NOR2X1 g56531(.A (WX6998), .B (n_5811), .Y (n_9824));
INVX1 g57311(.A (WX535), .Y (n_5257));
NOR2X1 g56566(.A (WX8291), .B (n_2620), .Y (n_5219));
NOR2X1 g56571(.A (WX8291), .B (n_4882), .Y (n_8542));
NOR2X1 g56633(.A (WX9584), .B (n_2849), .Y (n_5217));
NOR2X1 g56635(.A (WX9584), .B (n_5427), .Y (n_8553));
DFFSRX1 WX9702_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6505), .Q (WX9702), .QN ());
DFFSRX1 WX4538_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5194), .Q (WX4538), .QN ());
DFFSRX1 WX3247_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5191), .Q (WX3247), .QN ());
DFFSRX1 WX5829_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5193), .Q (WX5829), .QN ());
DFFSRX1 WX8411_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5197), .Q (WX8411), .QN ());
DFFSRX1 WX7120_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5192), .Q (WX7120), .QN ());
NOR2X1 g56332(.A (WX3119), .B (n_5427), .Y (n_5214));
NOR2X1 g56455(.A (WX4414), .B (n_2605), .Y (n_5213));
NOR2X1 g56460(.A (WX4414), .B (n_5662), .Y (n_5212));
OAI21X1 g56467(.A0 (n_4238), .A1 (n_8543), .B0 (n_5722), .Y (n_5211));
DFFSRX1 WX8247_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5182), .Q (), .QN (WX8247));
DFFSRX1 WX4374_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5177), .Q (), .QN (WX4374));
DFFSRX1 WX5665_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5173), .Q (), .QN (WX5665));
DFFSRX1 WX6956_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5171), .Q (), .QN (WX6956));
DFFSRX1 WX3083_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5169), .Q (), .QN (WX3083));
NOR2X1 g57219(.A (WX10877), .B (n_2620), .Y (n_5210));
NOR2X1 g57220(.A (WX1826), .B (n_2620), .Y (n_5208));
NOR2X1 g57231(.A (WX1826), .B (n_5838), .Y (n_5207));
NOR2X1 g57234(.A (WX10877), .B (n_5662), .Y (n_6682));
NAND2X1 g57262(.A (n_5166), .B (n_4693), .Y (n_5204));
OAI21X1 g56532(.A0 (n_15859), .A1 (n_15860), .B0 (n_5619), .Y(n_5203));
DFFSRX1 WX535_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5162), .Q (WX535), .QN ());
OAI21X1 g56572(.A0 (n_4112), .A1 (n_8554), .B0 (n_5556), .Y (n_5201));
OAI21X1 g56636(.A0 (n_5135), .A1 (n_11595), .B0 (n_5619), .Y(n_5200));
DFFSRX1 WX3283_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5186), .Q (WX3283), .QN ());
DFFSRX1 WX5869_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5184), .Q (WX5869), .QN ());
DFFSRX1 WX7162_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5165), .Q (WX7162), .QN ());
DFFSRX1 WX8455_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5159), .Q (WX8455), .QN ());
DFFSRX1 WX9748_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5157), .Q (WX9748), .QN ());
DFFSRX1 WX9538_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5179), .Q (), .QN (WX9538));
OAI21X1 g56333(.A0 (n_5156), .A1 (n_9415), .B0 (n_5460), .Y (n_5199));
DFFSRX1 WX3119_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5154), .Q (), .QN (WX3119));
OAI21X1 g56461(.A0 (n_15861), .A1 (n_15862), .B0 (n_5722), .Y(n_5198));
DFFSRX1 WX5705_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5143), .Q (), .QN (WX5705));
OAI21X1 g57193(.A0 (n_4313), .A1 (n_5196), .B0 (n_5152), .Y (n_5197));
OAI21X1 g57195(.A0 (n_4494), .A1 (n_5334), .B0 (n_5150), .Y (n_5194));
OAI21X1 g57196(.A0 (n_4433), .A1 (n_5928), .B0 (n_5149), .Y (n_5193));
OAI21X1 g57198(.A0 (n_4375), .A1 (n_5254), .B0 (n_5148), .Y (n_5192));
OAI21X1 g57199(.A0 (n_4337), .A1 (n_5235), .B0 (n_5146), .Y (n_5191));
OAI21X1 g57232(.A0 (n_5126), .A1 (n_4145), .B0 (n_5722), .Y (n_5190));
OAI21X1 g57235(.A0 (n_4505), .A1 (n_6680), .B0 (n_4860), .Y (n_5189));
DFFSRX1 WX6998_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5141), .Q (), .QN (WX6998));
MX2X1 g57334(.A (n_5161), .B (WX537), .S0 (n_10743), .Y (n_5187));
DFFSRX1 WX8291_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5139), .Q (), .QN (WX8291));
DFFSRX1 WX9584_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5136), .Q (), .QN (WX9584));
DFFSRX1 WX4578_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5153), .Q (WX4578), .QN ());
DFFSRX1 WX11041_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5144), .Q (WX11041), .QN ());
DFFSRX1 WX1990_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5145), .Q (WX1990), .QN ());
OAI21X1 g56366(.A0 (n_4301), .A1 (n_5185), .B0 (n_5133), .Y (n_5186));
DFFSRX1 WX4414_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5132), .Q (), .QN (WX4414));
OAI21X1 g56489(.A0 (n_4662), .A1 (n_5183), .B0 (n_5129), .Y (n_5184));
NOR2X1 g57216(.A (WX8249), .B (n_5181), .Y (n_5182));
NOR2X1 g57217(.A (WX8249), .B (n_5500), .Y (n_5180));
NOR2X1 g57221(.A (WX9540), .B (n_2851), .Y (n_5179));
NOR2X1 g57222(.A (WX4376), .B (n_2851), .Y (n_5177));
NOR2X1 g57223(.A (WX9540), .B (n_5500), .Y (n_6222));
NOR2X1 g57225(.A (WX4376), .B (n_5811), .Y (n_6223));
NOR2X1 g57228(.A (WX5667), .B (n_1648), .Y (n_5173));
NOR2X1 g57229(.A (WX5667), .B (n_5811), .Y (n_6224));
NOR2X1 g57237(.A (WX6958), .B (n_5712), .Y (n_5171));
NOR2X1 g57239(.A (WX6958), .B (n_5662), .Y (n_6674));
NOR2X1 g57241(.A (WX3085), .B (n_1648), .Y (n_5169));
NOR2X1 g57242(.A (WX3085), .B (n_5811), .Y (n_6225));
DFFSRX1 WX1826_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5127), .Q (), .QN (WX1826));
DFFSRX1 WX10877_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5128), .Q (), .QN (WX10877));
NAND2X1 g57303(.A (n_5123), .B (n_6615), .Y (n_5166));
OAI21X1 g56549(.A0 (n_4111), .A1 (n_5928), .B0 (n_5122), .Y (n_5165));
INVX1 g57335(.A (DATA_9_4), .Y (n_5164));
NOR2X1 g57360(.A (n_1425), .B (n_5161), .Y (n_5162));
OR2X1 g57369(.A (n_5161), .B (n_5990), .Y (n_5160));
OAI21X1 g56604(.A0 (n_4281), .A1 (n_5158), .B0 (n_5121), .Y (n_5159));
OAI21X1 g56664(.A0 (n_4265), .A1 (n_5490), .B0 (n_5119), .Y (n_5157));
NOR2X1 g56391(.A (WX3121), .B (n_5427), .Y (n_5156));
NOR2X1 g56412(.A (WX3121), .B (n_3188), .Y (n_5154));
OAI21X1 g56488(.A0 (n_4235), .A1 (n_5825), .B0 (n_5111), .Y (n_5153));
OAI21X1 g57218(.A0 (n_4376), .A1 (n_6227), .B0 (n_4860), .Y (n_5152));
OAI21X1 g57226(.A0 (n_4338), .A1 (n_6195), .B0 (n_5619), .Y (n_5150));
OAI21X1 g57230(.A0 (n_4497), .A1 (n_6226), .B0 (n_5566), .Y (n_5149));
OAI21X1 g57240(.A0 (n_4434), .A1 (n_6228), .B0 (n_4947), .Y (n_5148));
OAI21X1 g57243(.A0 (n_4487), .A1 (n_6675), .B0 (n_3183), .Y (n_5146));
OAI21X1 g57259(.A0 (n_4213), .A1 (n_5254), .B0 (n_5110), .Y (n_5145));
OAI21X1 g57263(.A0 (n_3810), .A1 (n_5320), .B0 (n_5109), .Y (n_5144));
NOR2X1 g56524(.A (WX5707), .B (n_2620), .Y (n_5143));
NOR2X1 g56525(.A (WX5707), .B (n_5838), .Y (n_8543));
OAI21X1 g57336(.A0 (n_5089), .A1 (n_6091), .B0 (n_4062), .Y(DATA_9_4));
NOR2X1 g56589(.A (WX7000), .B (n_5712), .Y (n_5141));
NOR2X1 g56591(.A (WX7000), .B (n_5500), .Y (n_15860));
DFFSRX1 WX5831_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5113), .Q (WX5831), .QN ());
NOR2X1 g56626(.A (WX8293), .B (n_5181), .Y (n_5139));
NOR2X1 g56631(.A (WX8293), .B (n_5479), .Y (n_8554));
NOR2X1 g56692(.A (WX9586), .B (n_1425), .Y (n_5136));
NOR2X1 g56694(.A (WX9586), .B (n_5662), .Y (n_5135));
DFFSRX1 WX3249_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5118), .Q (WX3249), .QN ());
DFFSRX1 WX8413_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5117), .Q (WX8413), .QN ());
DFFSRX1 WX9704_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5116), .Q (WX9704), .QN ());
DFFSRX1 WX4540_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5115), .Q (WX4540), .QN ());
DFFSRX1 WX7122_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5112), .Q (WX7122), .QN ());
DFFSRX1 WX703_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5107), .Q (WX703), .QN ());
OAI21X1 g56392(.A0 (n_5084), .A1 (n_11626), .B0 (n_5722), .Y(n_5133));
DFFSRX1 WX8249_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5104), .Q (), .QN (WX8249));
DFFSRX1 WX9540_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5102), .Q (), .QN (WX9540));
DFFSRX1 WX4376_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5100), .Q (), .QN (WX4376));
DFFSRX1 WX5667_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5097), .Q (), .QN (WX5667));
DFFSRX1 WX6958_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5095), .Q (), .QN (WX6958));
DFFSRX1 WX3085_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5092), .Q (), .QN (WX3085));
NOR2X1 g56514(.A (WX4416), .B (n_1425), .Y (n_5132));
NOR2X1 g56519(.A (WX4416), .B (n_5500), .Y (n_15862));
OAI21X1 g56526(.A0 (n_4236), .A1 (n_12492), .B0 (n_7087), .Y(n_5129));
NOR2X1 g57285(.A (WX10879), .B (n_1648), .Y (n_5128));
NOR2X1 g57286(.A (WX1828), .B (n_3188), .Y (n_5127));
NOR2X1 g57297(.A (WX1828), .B (n_4882), .Y (n_5126));
NOR2X1 g57299(.A (WX10879), .B (n_5427), .Y (n_6680));
OAI21X1 g57333(.A0 (n_5069), .A1 (n_5889), .B0 (n_4961), .Y (n_5123));
OAI21X1 g56565(.A0 (n_5064), .A1 (n_4661), .B0 (n_5556), .Y (n_5122));
INVX1 g57382(.A (WX537), .Y (n_5161));
OAI21X1 g56632(.A0 (n_5060), .A1 (n_10713), .B0 (n_5556), .Y(n_5121));
OAI21X1 g56695(.A0 (n_4280), .A1 (n_12493), .B0 (n_5619), .Y(n_5119));
DFFSRX1 WX3285_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5106), .Q (WX3285), .QN ());
DFFSRX1 WX5871_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5090), .Q (WX5871), .QN ());
DFFSRX1 WX7164_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5088), .Q (WX7164), .QN ());
DFFSRX1 WX8457_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5087), .Q (WX8457), .QN ());
DFFSRX1 WX9750_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5086), .Q (WX9750), .QN ());
DFFSRX1 WX3121_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5083), .Q (), .QN (WX3121));
OAI21X1 g57254(.A0 (n_4647), .A1 (n_5158), .B0 (n_5082), .Y (n_5118));
OAI21X1 g57255(.A0 (n_4611), .A1 (n_5235), .B0 (n_5081), .Y (n_5117));
OAI21X1 g57256(.A0 (n_4548), .A1 (n_5239), .B0 (n_5080), .Y (n_5116));
OAI21X1 g57257(.A0 (n_4492), .A1 (n_5439), .B0 (n_5079), .Y (n_5115));
OAI21X1 g57258(.A0 (n_4431), .A1 (n_5879), .B0 (n_5078), .Y (n_5113));
OAI21X1 g57260(.A0 (n_4132), .A1 (n_5879), .B0 (n_5076), .Y (n_5112));
OAI21X1 g56520(.A0 (n_4578), .A1 (n_6694), .B0 (n_7087), .Y (n_5111));
OAI21X1 g57298(.A0 (n_5053), .A1 (n_4143), .B0 (n_5460), .Y (n_5110));
OAI21X1 g57300(.A0 (n_4264), .A1 (n_7507), .B0 (n_5460), .Y (n_5109));
DFFSRX1 WX5707_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5071), .Q (), .QN (WX5707));
NAND2X2 g57326(.A (n_5072), .B (n_4692), .Y (n_5107));
DFFSRX1 WX537_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5067), .Q (WX537), .QN ());
DFFSRX1 WX7000_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5063), .Q (), .QN (WX7000));
DFFSRX1 WX8293_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5062), .Q (), .QN (WX8293));
DFFSRX1 WX9586_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5059), .Q (), .QN (WX9586));
DFFSRX1 WX4580_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5075), .Q (WX4580), .QN ());
DFFSRX1 WX11043_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5073), .Q (WX11043), .QN ());
DFFSRX1 WX1992_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5074), .Q (WX1992), .QN ());
OAI21X1 g56425(.A0 (n_4580), .A1 (n_5105), .B0 (n_5056), .Y (n_5106));
NOR2X1 g57282(.A (WX8251), .B (n_5712), .Y (n_5104));
NOR2X1 g57283(.A (WX8251), .B (n_5811), .Y (n_6227));
NOR2X1 g57287(.A (WX9542), .B (n_1425), .Y (n_5102));
NOR2X1 g57288(.A (WX4378), .B (n_5181), .Y (n_5100));
NOR2X1 g57291(.A (WX4378), .B (n_4882), .Y (n_6195));
NOR2X1 g57294(.A (WX5669), .B (n_5712), .Y (n_5097));
NOR2X1 g57295(.A (WX5669), .B (n_4882), .Y (n_6226));
NOR2X1 g57301(.A (WX6960), .B (n_5712), .Y (n_5095));
DFFSRX1 WX4416_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5050), .Q (), .QN (WX4416));
NOR2X1 g57304(.A (WX6960), .B (n_5822), .Y (n_6228));
NOR2X1 g57305(.A (WX3087), .B (n_1648), .Y (n_5092));
NOR2X1 g57307(.A (WX3087), .B (n_5427), .Y (n_6675));
DFFSRX1 WX10879_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5055), .Q (), .QN (WX10879));
DFFSRX1 WX1828_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5054), .Q (), .QN (WX1828));
OAI21X1 g56548(.A0 (n_4211), .A1 (n_5649), .B0 (n_5047), .Y (n_5090));
MX2X1 g57400(.A (n_5066), .B (WX539), .S0 (n_4061), .Y (n_5089));
OAI21X1 g56602(.A0 (n_4326), .A1 (n_5841), .B0 (n_5046), .Y (n_5088));
OAI21X1 g56663(.A0 (n_4565), .A1 (n_5576), .B0 (n_5045), .Y (n_5087));
OAI21X1 g56722(.A0 (n_4263), .A1 (n_5085), .B0 (n_5043), .Y (n_5086));
NOR2X1 g56450(.A (WX3123), .B (n_5427), .Y (n_5084));
NOR2X1 g56471(.A (WX3123), .B (n_5712), .Y (n_5083));
OAI21X1 g57281(.A0 (n_5028), .A1 (n_4252), .B0 (n_5566), .Y (n_5082));
OAI21X1 g57284(.A0 (n_4374), .A1 (n_6197), .B0 (n_5460), .Y (n_5081));
OAI21X1 g57290(.A0 (n_5022), .A1 (n_4312), .B0 (n_4947), .Y (n_5080));
OAI21X1 g57292(.A0 (n_4336), .A1 (n_6229), .B0 (n_3183), .Y (n_5079));
OAI21X1 g57296(.A0 (n_4493), .A1 (n_6196), .B0 (n_4860), .Y (n_5078));
OAI21X1 g57306(.A0 (n_4432), .A1 (n_6672), .B0 (n_4947), .Y (n_5076));
OAI21X1 g56546(.A0 (n_4233), .A1 (n_5235), .B0 (n_5034), .Y (n_5075));
OAI21X1 g57324(.A0 (n_4394), .A1 (n_5892), .B0 (n_5036), .Y (n_5074));
OAI21X1 g57330(.A0 (n_3818), .A1 (n_5439), .B0 (n_5035), .Y (n_5073));
NAND2X1 g57371(.A (n_6615), .B (n_8320), .Y (n_5072));
NOR2X1 g56584(.A (WX5709), .B (n_5181), .Y (n_5071));
NOR2X1 g56585(.A (WX5709), .B (n_5052), .Y (n_12492));
INVX1 g57402(.A (DATA_9_3), .Y (n_5069));
NOR2X1 g57450(.A (n_5181), .B (n_5066), .Y (n_5067));
OR2X1 g57457(.A (n_5066), .B (n_3828), .Y (n_5065));
NOR2X1 g56624(.A (WX7002), .B (n_5500), .Y (n_5064));
NOR2X1 g56649(.A (WX7002), .B (n_1425), .Y (n_5063));
NOR2X1 g56685(.A (WX8295), .B (n_5181), .Y (n_5062));
NOR2X1 g56690(.A (WX8295), .B (n_5662), .Y (n_5060));
NOR2X1 g56750(.A (WX9588), .B (n_5712), .Y (n_5059));
NOR2X1 g56752(.A (WX9588), .B (n_5427), .Y (n_12493));
DFFSRX1 WX5833_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5038), .Q (WX5833), .QN ());
DFFSRX1 WX3251_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5042), .Q (WX3251), .QN ());
DFFSRX1 WX8415_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5041), .Q (WX8415), .QN ());
DFFSRX1 WX9706_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5040), .Q (WX9706), .QN ());
DFFSRX1 WX4542_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5039), .Q (WX4542), .QN ());
DFFSRX1 WX7124_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5037), .Q (WX7124), .QN ());
OAI21X1 g56451(.A0 (n_15863), .A1 (n_15864), .B0 (n_5566), .Y(n_5056));
DFFSRX1 WX8251_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5027), .Q (), .QN (WX8251));
DFFSRX1 WX9542_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5025), .Q (), .QN (WX9542));
DFFSRX1 WX4378_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5024), .Q (), .QN (WX4378));
DFFSRX1 WX5669_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5020), .Q (), .QN (WX5669));
DFFSRX1 WX6960_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5017), .Q (), .QN (WX6960));
DFFSRX1 WX3087_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5016), .Q (), .QN (WX3087));
NOR2X1 g57350(.A (WX10881), .B (n_5181), .Y (n_5055));
NOR2X1 g57351(.A (WX1830), .B (n_2620), .Y (n_5054));
NOR2X1 g57364(.A (WX1830), .B (n_5052), .Y (n_5053));
NOR2X1 g57367(.A (WX10881), .B (n_5811), .Y (n_7507));
NOR2X1 g56574(.A (WX4418), .B (n_3188), .Y (n_5050));
NOR2X1 g56578(.A (WX4418), .B (n_5822), .Y (n_6694));
OAI21X1 g56586(.A0 (n_4992), .A1 (n_10717), .B0 (n_6497), .Y(n_5047));
OAI21X1 g57403(.A0 (n_4991), .A1 (n_5965), .B0 (n_4060), .Y(DATA_9_3));
OAI21X1 g56625(.A0 (n_4210), .A1 (n_8544), .B0 (n_4947), .Y (n_5046));
OAI21X1 g56691(.A0 (n_4985), .A1 (n_4325), .B0 (n_5566), .Y (n_5045));
OAI21X1 g56753(.A0 (n_4564), .A1 (n_6695), .B0 (n_5706), .Y (n_5043));
DFFSRX1 WX3287_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5030), .Q (WX3287), .QN ());
DFFSRX1 WX5873_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5012), .Q (WX5873), .QN ());
DFFSRX1 WX7166_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5011), .Q (WX7166), .QN ());
DFFSRX1 WX8459_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5010), .Q (WX8459), .QN ());
DFFSRX1 WX9752_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5009), .Q (WX9752), .QN ());
DFFSRX1 WX705_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_6621), .Q (WX705), .QN ());
DFFSRX1 WX3123_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_5007), .Q (), .QN (WX3123));
OAI21X1 g57318(.A0 (n_4642), .A1 (n_5879), .B0 (n_5005), .Y (n_5042));
OAI21X1 g57319(.A0 (n_4609), .A1 (n_5474), .B0 (n_5004), .Y (n_5041));
OAI21X1 g57321(.A0 (n_4546), .A1 (n_5841), .B0 (n_5003), .Y (n_5040));
OAI21X1 g57322(.A0 (n_4490), .A1 (n_5105), .B0 (n_5001), .Y (n_5039));
OAI21X1 g57323(.A0 (n_4429), .A1 (n_5493), .B0 (n_4999), .Y (n_5038));
OAI21X1 g57325(.A0 (n_4130), .A1 (n_5183), .B0 (n_4998), .Y (n_5037));
OAI21X1 g57365(.A0 (n_4973), .A1 (n_4141), .B0 (n_5460), .Y (n_5036));
OAI21X1 g57370(.A0 (n_4262), .A1 (n_7508), .B0 (n_4860), .Y (n_5035));
OAI21X1 g56579(.A0 (n_15865), .A1 (n_15866), .B0 (n_5556), .Y(n_5034));
OAI21X1 g57397(.A0 (n_4966), .A1 (n_5889), .B0 (n_4873), .Y (n_8320));
DFFSRX1 WX5709_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4994), .Q (), .QN (WX5709));
INVX1 g57468(.A (WX539), .Y (n_5066));
DFFSRX1 WX7002_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4988), .Q (), .QN (WX7002));
DFFSRX1 WX8295_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4986), .Q (), .QN (WX8295));
DFFSRX1 WX9588_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4984), .Q (), .QN (WX9588));
DFFSRX1 WX4582_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4995), .Q (WX4582), .QN ());
DFFSRX1 WX11045_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4996), .Q (WX11045), .QN ());
DFFSRX1 WX1994_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4997), .Q (WX1994), .QN ());
OAI21X1 g56484(.A0 (n_4297), .A1 (n_5928), .B0 (n_4979), .Y (n_5030));
NOR2X1 g57345(.A (WX3089), .B (n_5822), .Y (n_5028));
NOR2X1 g57347(.A (WX8253), .B (n_5712), .Y (n_5027));
NOR2X1 g57348(.A (WX8253), .B (n_5811), .Y (n_6197));
NOR2X1 g57354(.A (WX9544), .B (n_1425), .Y (n_5025));
NOR2X1 g57355(.A (WX4380), .B (n_3188), .Y (n_5024));
NOR2X1 g57356(.A (WX9544), .B (n_5500), .Y (n_5022));
NOR2X1 g57358(.A (WX4380), .B (n_5052), .Y (n_6229));
NOR2X1 g57361(.A (WX5671), .B (n_2620), .Y (n_5020));
NOR2X1 g57362(.A (WX5671), .B (n_5052), .Y (n_6196));
NOR2X1 g57368(.A (WX6962), .B (n_5712), .Y (n_5017));
NOR2X1 g57374(.A (WX3089), .B (n_2849), .Y (n_5016));
NOR2X1 g57375(.A (WX6962), .B (n_5500), .Y (n_6672));
DFFSRX1 WX10881_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4976), .Q (), .QN (WX10881));
DFFSRX1 WX1830_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4974), .Q (), .QN (WX1830));
DFFSRX1 WX4418_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4970), .Q (), .QN (WX4418));
OAI21X1 g56608(.A0 (n_4392), .A1 (n_5886), .B0 (n_4968), .Y (n_5012));
DFFSRX1 WX539_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4964), .Q (WX539), .QN ());
OAI21X1 g56661(.A0 (n_4324), .A1 (n_5830), .B0 (n_4962), .Y (n_5011));
OAI21X1 g56721(.A0 (n_4563), .A1 (n_5085), .B0 (n_4959), .Y (n_5010));
OAI21X1 g56782(.A0 (n_4504), .A1 (n_4803), .B0 (n_4958), .Y (n_5009));
DFFSRX1 WX649_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4960), .Q (WX649), .QN ());
DFFSRX1 WX647_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4956), .Q (WX647), .QN ());
DFFSRX1 WX645_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4980), .Q (WX645), .QN ());
DFFSRX1 WX707_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4978), .Q (WX707), .QN ());
NOR2X1 g56509(.A (WX3125), .B (n_5662), .Y (n_15864));
NOR2X1 g56530(.A (WX3125), .B (n_5712), .Y (n_5007));
OAI21X1 g57346(.A0 (n_4939), .A1 (n_4250), .B0 (n_4947), .Y (n_5005));
OAI21X1 g57349(.A0 (n_4936), .A1 (n_4131), .B0 (n_5460), .Y (n_5004));
OAI21X1 g57357(.A0 (n_4610), .A1 (n_6231), .B0 (n_4860), .Y (n_5003));
OAI21X1 g57359(.A0 (n_4646), .A1 (n_6198), .B0 (n_4947), .Y (n_5001));
OAI21X1 g57363(.A0 (n_4491), .A1 (n_6230), .B0 (n_4860), .Y (n_4999));
OAI21X1 g57376(.A0 (n_4924), .A1 (n_4430), .B0 (n_4947), .Y (n_4998));
OAI21X1 g57393(.A0 (n_4205), .A1 (n_5105), .B0 (n_4949), .Y (n_4997));
OAI21X1 g57396(.A0 (n_3809), .A1 (n_5418), .B0 (n_4948), .Y (n_4996));
OAI21X1 g56606(.A0 (n_4458), .A1 (n_5239), .B0 (n_4946), .Y (n_4995));
NOR2X1 g56643(.A (WX5711), .B (n_5181), .Y (n_4994));
NOR2X1 g56645(.A (WX5711), .B (n_5500), .Y (n_4992));
MX2X1 g57508(.A (n_4963), .B (WX541), .S0 (n_6613), .Y (n_4991));
NOR2X1 g56683(.A (WX7004), .B (n_4882), .Y (n_8544));
NOR2X1 g56708(.A (WX7004), .B (n_2620), .Y (n_4988));
DFFSRX1 WX7126_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4950), .Q (WX7126), .QN ());
NOR2X1 g56744(.A (WX8297), .B (n_3690), .Y (n_4986));
NOR2X1 g56748(.A (WX8297), .B (n_5427), .Y (n_4985));
NOR2X1 g56808(.A (WX9590), .B (n_3188), .Y (n_4984));
NOR2X1 g56811(.A (WX9590), .B (n_5662), .Y (n_6695));
DFFSRX1 WX8417_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4954), .Q (WX8417), .QN ());
DFFSRX1 WX9708_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4953), .Q (WX9708), .QN ());
DFFSRX1 WX3253_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4955), .Q (WX3253), .QN ());
DFFSRX1 WX5835_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4951), .Q (WX5835), .QN ());
DFFSRX1 WX4544_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4952), .Q (WX4544), .QN ());
DFFSRX1 WX3289_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4942), .Q (WX3289), .QN ());
NAND2X1 g57200(.A (n_4944), .B (n_4745), .Y (n_4980));
OAI21X1 g56510(.A0 (n_4204), .A1 (n_12494), .B0 (n_5722), .Y(n_4979));
NAND2X2 g57328(.A (n_4941), .B (n_4690), .Y (n_4978));
DFFSRX1 WX8253_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4938), .Q (), .QN (WX8253));
DFFSRX1 WX9544_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4935), .Q (), .QN (WX9544));
DFFSRX1 WX4380_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4934), .Q (), .QN (WX4380));
DFFSRX1 WX5671_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4930), .Q (), .QN (WX5671));
DFFSRX1 WX6962_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4927), .Q (), .QN (WX6962));
DFFSRX1 WX3089_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4925), .Q (), .QN (WX3089));
NOR2X1 g57439(.A (WX10883), .B (n_5712), .Y (n_4976));
NOR2X1 g57440(.A (WX1832), .B (n_5712), .Y (n_4974));
NOR2X1 g57454(.A (WX1832), .B (n_5662), .Y (n_4973));
NOR2X1 g57458(.A (WX10883), .B (n_5479), .Y (n_7508));
NOR2X1 g56634(.A (WX4420), .B (n_5712), .Y (n_4970));
NOR2X1 g56637(.A (WX4420), .B (n_5479), .Y (n_15866));
OAI21X1 g56646(.A0 (n_4905), .A1 (n_4232), .B0 (n_4947), .Y (n_4968));
INVX1 g57510(.A (DATA_9_2), .Y (n_4966));
NOR2X1 g57544(.A (n_2849), .B (n_4963), .Y (n_4964));
OAI21X1 g56684(.A0 (n_4904), .A1 (n_10719), .B0 (n_5566), .Y(n_4962));
OR2X1 g57583(.A (n_4963), .B (n_5968), .Y (n_4961));
NAND2X2 g55783(.A (n_4943), .B (n_4728), .Y (n_4960));
OAI21X1 g56749(.A0 (n_4323), .A1 (n_8545), .B0 (n_5619), .Y (n_4959));
OAI21X1 g56812(.A0 (n_15867), .A1 (n_15868), .B0 (n_4860), .Y(n_4958));
DFFSRX1 WX5875_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4923), .Q (WX5875), .QN ());
DFFSRX1 WX7168_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4922), .Q (WX7168), .QN ());
DFFSRX1 WX8461_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4921), .Q (WX8461), .QN ());
DFFSRX1 WX9754_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4920), .Q (WX9754), .QN ());
NAND2X2 g55780(.A (n_4945), .B (n_4729), .Y (n_4956));
DFFSRX1 WX3125_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4918), .Q (), .QN (WX3125));
OAI21X1 g57387(.A0 (n_4636), .A1 (n_5841), .B0 (n_4917), .Y (n_4955));
OAI21X1 g57388(.A0 (n_4606), .A1 (n_5549), .B0 (n_4916), .Y (n_4954));
OAI21X1 g57390(.A0 (n_4544), .A1 (n_5415), .B0 (n_4915), .Y (n_4953));
OAI21X1 g57391(.A0 (n_4486), .A1 (n_5415), .B0 (n_4913), .Y (n_4952));
OAI21X1 g57392(.A0 (n_4427), .A1 (n_5439), .B0 (n_4912), .Y (n_4951));
OAI21X1 g57395(.A0 (n_4128), .A1 (n_5415), .B0 (n_4911), .Y (n_4950));
OAI21X1 g57455(.A0 (n_4887), .A1 (n_4139), .B0 (n_5460), .Y (n_4949));
OAI21X1 g57459(.A0 (n_4503), .A1 (n_6681), .B0 (n_4947), .Y (n_4948));
OAI21X1 g56638(.A0 (n_4883), .A1 (n_4570), .B0 (n_5460), .Y (n_4946));
OAI21X1 g57511(.A0 (n_4876), .A1 (n_5709), .B0 (n_4053), .Y(DATA_9_2));
DFFSRX1 WX5711_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4906), .Q (), .QN (WX5711));
DFFSRX1 WX7004_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4903), .Q (), .QN (WX7004));
DFFSRX1 WX8297_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4902), .Q (), .QN (WX8297));
DFFSRX1 WX4584_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4907), .Q (WX4584), .QN ());
DFFSRX1 WX11047_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4908), .Q (WX11047), .QN ());
DFFSRX1 WX1996_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4909), .Q (WX1996), .QN ());
DFFSRX1 WX9590_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4899), .Q (), .QN (WX9590));
NAND2X1 g55782(.A (n_6555), .B (n_8336), .Y (n_4945));
NAND2X1 g57233(.A (n_6583), .B (n_8337), .Y (n_4944));
NAND2X1 g55794(.A (n_4888), .B (n_6555), .Y (n_4943));
OAI21X1 g56543(.A0 (n_4571), .A1 (n_5600), .B0 (n_4893), .Y (n_4942));
NAND2X1 g57373(.A (n_6615), .B (n_8322), .Y (n_4941));
NOR2X1 g57434(.A (WX3091), .B (n_5500), .Y (n_4939));
NOR2X1 g57436(.A (WX8255), .B (n_5712), .Y (n_4938));
NOR2X1 g57437(.A (WX8255), .B (n_5500), .Y (n_4936));
NOR2X1 g57443(.A (WX9546), .B (n_3188), .Y (n_4935));
NOR2X1 g57444(.A (WX4382), .B (n_2851), .Y (n_4934));
NOR2X1 g57445(.A (WX9546), .B (n_4882), .Y (n_6231));
NOR2X1 g57447(.A (WX4382), .B (n_4882), .Y (n_6198));
NOR2X1 g57451(.A (WX5673), .B (n_2851), .Y (n_4930));
NOR2X1 g57452(.A (WX5673), .B (n_5479), .Y (n_6230));
NOR2X1 g57456(.A (WX6964), .B (n_1425), .Y (n_4927));
NOR2X1 g57460(.A (WX3091), .B (n_3188), .Y (n_4925));
NOR2X1 g57461(.A (WX6964), .B (n_5822), .Y (n_4924));
DFFSRX1 WX10883_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4891), .Q (), .QN (WX10883));
DFFSRX1 WX1832_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4890), .Q (), .QN (WX1832));
DFFSRX1 WX4420_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4884), .Q (), .QN (WX4420));
OAI21X1 g56667(.A0 (n_4209), .A1 (n_5468), .B0 (n_4881), .Y (n_4923));
INVX1 g57605(.A (WX541), .Y (n_4963));
OAI21X1 g56720(.A0 (n_4645), .A1 (n_5535), .B0 (n_4880), .Y (n_4922));
OAI21X1 g56780(.A0 (n_4279), .A1 (n_5439), .B0 (n_4879), .Y (n_4921));
OAI21X1 g56841(.A0 (n_4261), .A1 (n_5845), .B0 (n_4877), .Y (n_4920));
NOR2X1 g56569(.A (WX3127), .B (n_5811), .Y (n_12494));
NOR2X1 g56590(.A (WX3127), .B (n_1425), .Y (n_4918));
OAI21X1 g57435(.A0 (n_4473), .A1 (n_6232), .B0 (n_5556), .Y (n_4917));
OAI21X1 g57438(.A0 (n_4853), .A1 (n_4129), .B0 (n_5556), .Y (n_4916));
OAI21X1 g57446(.A0 (n_4607), .A1 (n_6199), .B0 (n_5619), .Y (n_4915));
OAI21X1 g57448(.A0 (n_4641), .A1 (n_6200), .B0 (n_5619), .Y (n_4913));
OAI21X1 g57453(.A0 (n_4489), .A1 (n_6676), .B0 (n_4860), .Y (n_4912));
OAI21X1 g57462(.A0 (n_4842), .A1 (n_4428), .B0 (n_5460), .Y (n_4911));
OAI21X1 g57496(.A0 (n_4203), .A1 (n_6050), .B0 (n_4861), .Y (n_4909));
OAI21X1 g57503(.A0 (n_3808), .A1 (n_5549), .B0 (n_4859), .Y (n_4908));
OAI21X1 g56665(.A0 (n_4456), .A1 (n_5598), .B0 (n_4858), .Y (n_4907));
DFFSRX1 WX541_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4875), .Q (WX541), .QN ());
NOR2X1 g56701(.A (WX5713), .B (n_1648), .Y (n_4906));
NOR2X1 g56704(.A (WX5713), .B (n_5479), .Y (n_4905));
NOR2X1 g56742(.A (WX7006), .B (n_5662), .Y (n_4904));
NOR2X1 g56766(.A (WX7006), .B (n_5181), .Y (n_4903));
NOR2X1 g56803(.A (WX8299), .B (n_1425), .Y (n_4902));
NOR2X1 g56806(.A (WX8299), .B (n_5479), .Y (n_8545));
DFFSRX1 WX3255_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4871), .Q (WX3255), .QN ());
DFFSRX1 WX8419_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4870), .Q (WX8419), .QN ());
DFFSRX1 WX9710_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4869), .Q (WX9710), .QN ());
DFFSRX1 WX4546_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4867), .Q (WX4546), .QN ());
DFFSRX1 WX5837_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4865), .Q (WX5837), .QN ());
DFFSRX1 WX7128_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4864), .Q (WX7128), .QN ());
NOR2X1 g56867(.A (WX9592), .B (n_2620), .Y (n_4899));
NOR2X1 g56871(.A (WX9592), .B (n_5479), .Y (n_15868));
OAI21X1 g55784(.A0 (n_4790), .A1 (n_5889), .B0 (n_3653), .Y (n_8336));
OAI21X1 g57261(.A0 (n_4827), .A1 (n_5889), .B0 (n_3600), .Y (n_8337));
OAI21X1 g56570(.A0 (n_4819), .A1 (n_11600), .B0 (n_5722), .Y(n_4893));
OAI21X1 g57399(.A0 (n_4801), .A1 (n_5889), .B0 (n_3692), .Y (n_8322));
DFFSRX1 WX8255_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4854), .Q (), .QN (WX8255));
DFFSRX1 WX9546_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4852), .Q (), .QN (WX9546));
DFFSRX1 WX4382_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4851), .Q (), .QN (WX4382));
DFFSRX1 WX5673_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4848), .Q (), .QN (WX5673));
DFFSRX1 WX6964_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4845), .Q (), .QN (WX6964));
DFFSRX1 WX3091_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4844), .Q (), .QN (WX3091));
NOR2X1 g57524(.A (WX10885), .B (n_5712), .Y (n_4891));
NOR2X1 g57526(.A (WX1834), .B (n_3188), .Y (n_4890));
OAI21X1 g55804(.A0 (n_4832), .A1 (n_5889), .B0 (n_3686), .Y (n_4888));
NOR2X1 g57551(.A (WX1834), .B (n_4882), .Y (n_4887));
NOR2X1 g57588(.A (WX10885), .B (n_5838), .Y (n_6681));
NOR2X1 g56693(.A (WX4422), .B (n_3690), .Y (n_4884));
NOR2X1 g56696(.A (WX4422), .B (n_4882), .Y (n_4883));
OAI21X1 g56705(.A0 (n_4786), .A1 (n_4457), .B0 (n_4860), .Y (n_4881));
OAI21X1 g56743(.A0 (n_4208), .A1 (n_9438), .B0 (n_5275), .Y (n_4880));
OAI21X1 g56807(.A0 (n_4775), .A1 (n_4643), .B0 (n_5722), .Y (n_4879));
DFFSRX1 WX3291_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4857), .Q (WX3291), .QN ());
DFFSRX1 WX5877_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4841), .Q (WX5877), .QN ());
DFFSRX1 WX7170_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4840), .Q (WX7170), .QN ());
DFFSRX1 WX8463_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4839), .Q (WX8463), .QN ());
DFFSRX1 WX9756_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4838), .Q (WX9756), .QN ());
OAI21X1 g56872(.A0 (n_4835), .A1 (n_11602), .B0 (n_6497), .Y(n_4877));
MX2X1 g57867(.A (n_4874), .B (WX543), .S0 (n_4052), .Y (n_4876));
NOR2X1 g58169(.A (n_1425), .B (n_4874), .Y (n_4875));
OR2X1 g58174(.A (n_4874), .B (n_5990), .Y (n_4873));
DFFSRX1 WX1938_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4828), .Q (WX1938), .QN ());
DFFSRX1 WX9716_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4816), .Q (WX9716), .QN ());
DFFSRX1 WX8425_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4820), .Q (WX8425), .QN ());
DFFSRX1 WX3261_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4823), .Q (WX3261), .QN ());
DFFSRX1 WX3127_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4802), .Q (), .QN (WX3127));
OAI21X1 g57476(.A0 (n_4633), .A1 (n_5317), .B0 (n_4799), .Y (n_4871));
OAI21X1 g57480(.A0 (n_4604), .A1 (n_5317), .B0 (n_4797), .Y (n_4870));
OAI21X1 g57484(.A0 (n_4542), .A1 (n_4868), .B0 (n_4796), .Y (n_4869));
OAI21X1 g57488(.A0 (n_4255), .A1 (n_4866), .B0 (n_4795), .Y (n_4867));
OAI21X1 g57492(.A0 (n_4423), .A1 (n_5185), .B0 (n_4794), .Y (n_4865));
OAI21X1 g57499(.A0 (n_4373), .A1 (n_5482), .B0 (n_4793), .Y (n_4864));
INVX1 g57512(.A (DATA_9_1), .Y (n_4863));
OAI21X1 g57552(.A0 (n_4765), .A1 (n_4137), .B0 (n_4860), .Y (n_4861));
OAI21X1 g57589(.A0 (n_4260), .A1 (n_7509), .B0 (n_5722), .Y (n_4859));
OAI21X1 g56697(.A0 (n_4758), .A1 (n_4568), .B0 (n_4860), .Y (n_4858));
DFFSRX1 WX5713_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4788), .Q (), .QN (WX5713));
DFFSRX1 WX7006_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4781), .Q (), .QN (WX7006));
DFFSRX1 WX3293_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4798), .Q (WX3293), .QN ());
DFFSRX1 WX4586_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4792), .Q (WX4586), .QN ());
DFFSRX1 WX3231_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4791), .Q (WX3231), .QN ());
DFFSRX1 WX4524_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4785), .Q (WX4524), .QN ());
DFFSRX1 WX5879_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4784), .Q (WX5879), .QN ());
DFFSRX1 WX3233_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4783), .Q (WX3233), .QN ());
DFFSRX1 WX7172_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4780), .Q (WX7172), .QN ());
DFFSRX1 WX4526_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4779), .Q (WX4526), .QN ());
DFFSRX1 WX5817_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4778), .Q (WX5817), .QN ());
DFFSRX1 WX8465_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4774), .Q (WX8465), .QN ());
DFFSRX1 WX5819_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4773), .Q (WX5819), .QN ());
DFFSRX1 WX7110_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4772), .Q (WX7110), .QN ());
DFFSRX1 WX8403_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4834), .Q (WX8403), .QN ());
DFFSRX1 WX7112_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4833), .Q (WX7112), .QN ());
DFFSRX1 WX8405_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4830), .Q (WX8405), .QN ());
DFFSRX1 WX9698_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4829), .Q (WX9698), .QN ());
DFFSRX1 WX11049_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4804), .Q (WX11049), .QN ());
DFFSRX1 WX3259_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4824), .Q (WX3259), .QN ());
DFFSRX1 WX3257_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4825), .Q (WX3257), .QN ());
DFFSRX1 WX8421_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4822), .Q (WX8421), .QN ());
DFFSRX1 WX8423_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4821), .Q (WX8423), .QN ());
DFFSRX1 WX9714_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4817), .Q (WX9714), .QN ());
DFFSRX1 WX9712_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4818), .Q (WX9712), .QN ());
DFFSRX1 WX4550_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4814), .Q (WX4550), .QN ());
DFFSRX1 WX4548_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4815), .Q (WX4548), .QN ());
DFFSRX1 WX5841_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4811), .Q (WX5841), .QN ());
DFFSRX1 WX5839_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4812), .Q (WX5839), .QN ());
DFFSRX1 WX1998_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4809), .Q (WX1998), .QN ());
DFFSRX1 WX2000_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4808), .Q (WX2000), .QN ());
DFFSRX1 WX7130_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4807), .Q (WX7130), .QN ());
DFFSRX1 WX7132_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4806), .Q (WX7132), .QN ());
DFFSRX1 WX7134_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4805), .Q (WX7134), .QN ());
DFFSRX1 WX8299_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4777), .Q (), .QN (WX8299));
DFFSRX1 WX4552_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4813), .Q (WX4552), .QN ());
DFFSRX1 WX5843_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4810), .Q (WX5843), .QN ());
DFFSRX1 WX9592_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4837), .Q (), .QN (WX9592));
DFFSRX1 WX11051_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4760), .Q (WX11051), .QN ());
OAI21X1 g56603(.A0 (n_4569), .A1 (n_5158), .B0 (n_4761), .Y (n_4857));
OAI21X1 g57513(.A0 (n_4679), .A1 (n_5965), .B0 (n_4051), .Y(DATA_9_1));
NOR2X1 g57516(.A (WX3093), .B (n_5500), .Y (n_6232));
NOR2X1 g57521(.A (WX8257), .B (n_1425), .Y (n_4854));
NOR2X1 g57522(.A (WX8257), .B (n_5500), .Y (n_4853));
NOR2X1 g57529(.A (WX9548), .B (n_1648), .Y (n_4852));
NOR2X1 g57530(.A (WX4384), .B (n_5712), .Y (n_4851));
NOR2X1 g57531(.A (WX9548), .B (n_5500), .Y (n_6199));
NOR2X1 g57536(.A (WX4384), .B (n_5838), .Y (n_6200));
NOR2X1 g57545(.A (WX5675), .B (n_3690), .Y (n_4848));
NOR2X1 g57546(.A (WX5675), .B (n_4882), .Y (n_6676));
NOR2X1 g57580(.A (WX6966), .B (n_3690), .Y (n_4845));
NOR2X1 g57590(.A (WX3093), .B (n_1648), .Y (n_4844));
NOR2X1 g57591(.A (WX6966), .B (n_4670), .Y (n_4842));
DFFSRX1 WX1834_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4768), .Q (), .QN (WX1834));
DFFSRX1 WX10885_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4769), .Q (), .QN (WX10885));
DFFSRX1 WX4422_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4759), .Q (), .QN (WX4422));
OAI21X1 g56725(.A0 (n_4207), .A1 (n_5439), .B0 (n_4756), .Y (n_4841));
OAI21X1 g56779(.A0 (n_4640), .A1 (n_5729), .B0 (n_4755), .Y (n_4840));
DFFSRX1 WX10991_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4762), .Q (WX10991), .QN ());
DFFSRX1 WX1940_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4757), .Q (WX1940), .QN ());
DFFSRX1 WX9758_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4770), .Q (WX9758), .QN ());
OAI21X1 g56839(.A0 (n_4560), .A1 (n_5085), .B0 (n_4754), .Y (n_4839));
DFFSRX1 WX9696_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4766), .Q (WX9696), .QN ());
OAI21X1 g56899(.A0 (n_4259), .A1 (n_5334), .B0 (n_4771), .Y (n_4838));
NOR2X1 g56926(.A (WX9594), .B (n_1425), .Y (n_4837));
NOR2X1 g56929(.A (WX9594), .B (n_5427), .Y (n_4835));
DFFSRX1 WX10989_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4746), .Q (WX10989), .QN ());
OAI21X1 g56956(.A0 (n_4319), .A1 (n_6050), .B0 (n_4750), .Y (n_4834));
OAI21X1 g56961(.A0 (n_4383), .A1 (n_4868), .B0 (n_4749), .Y (n_4833));
INVX1 g55845(.A (DATA_9_29), .Y (n_4832));
OAI21X1 g57015(.A0 (n_4618), .A1 (n_4866), .B0 (n_4748), .Y (n_4830));
INVX1 g58206(.A (WX543), .Y (n_4874));
OAI21X1 g57075(.A0 (n_4275), .A1 (n_5183), .B0 (n_4747), .Y (n_4829));
OAI21X1 g57320(.A0 (n_4596), .A1 (n_5918), .B0 (n_4652), .Y (n_4828));
INVX1 g57331(.A (DATA_9_31), .Y (n_4827));
OAI21X1 g57477(.A0 (n_4631), .A1 (n_5928), .B0 (n_4651), .Y (n_4825));
OAI21X1 g57478(.A0 (n_4629), .A1 (n_5841), .B0 (n_4744), .Y (n_4824));
OAI21X1 g57479(.A0 (n_4624), .A1 (n_5439), .B0 (n_4743), .Y (n_4823));
OAI21X1 g57481(.A0 (n_4601), .A1 (n_4866), .B0 (n_4742), .Y (n_4822));
OAI21X1 g57482(.A0 (n_4598), .A1 (n_5474), .B0 (n_4741), .Y (n_4821));
OAI21X1 g57483(.A0 (n_4594), .A1 (n_5418), .B0 (n_4740), .Y (n_4820));
NOR2X1 g56629(.A (WX3129), .B (n_4882), .Y (n_4819));
OAI21X1 g57485(.A0 (n_4538), .A1 (n_5892), .B0 (n_4739), .Y (n_4818));
OAI21X1 g57486(.A0 (n_4626), .A1 (n_5490), .B0 (n_4738), .Y (n_4817));
OAI21X1 g57487(.A0 (n_4536), .A1 (n_4868), .B0 (n_4737), .Y (n_4816));
OAI21X1 g57489(.A0 (n_4484), .A1 (n_5535), .B0 (n_4736), .Y (n_4815));
OAI21X1 g57490(.A0 (n_4482), .A1 (n_5415), .B0 (n_4735), .Y (n_4814));
OAI21X1 g57491(.A0 (n_4480), .A1 (n_5482), .B0 (n_4734), .Y (n_4813));
OAI21X1 g57493(.A0 (n_4421), .A1 (n_5196), .B0 (n_4650), .Y (n_4812));
OAI21X1 g57494(.A0 (n_4416), .A1 (n_5493), .B0 (n_4733), .Y (n_4811));
OAI21X1 g57495(.A0 (n_4414), .A1 (n_5185), .B0 (n_4731), .Y (n_4810));
OAI21X1 g57497(.A0 (n_4201), .A1 (n_5576), .B0 (n_4730), .Y (n_4809));
OAI21X1 g57498(.A0 (n_4387), .A1 (n_5882), .B0 (n_4649), .Y (n_4808));
OAI21X1 g57500(.A0 (n_4371), .A1 (n_5598), .B0 (n_4689), .Y (n_4807));
OAI21X1 g57501(.A0 (n_4369), .A1 (n_5493), .B0 (n_4687), .Y (n_4806));
OAI21X1 g57502(.A0 (n_4365), .A1 (n_5882), .B0 (n_4686), .Y (n_4805));
OAI21X1 g57504(.A0 (n_3807), .A1 (n_4803), .B0 (n_4688), .Y (n_4804));
NOR2X1 g56650(.A (WX3129), .B (n_1425), .Y (n_4802));
INVX1 g57514(.A (DATA_9_0), .Y (n_4801));
OAI21X1 g57517(.A0 (n_4677), .A1 (n_4463), .B0 (n_5460), .Y (n_4799));
OAI21X1 g56662(.A0 (n_4567), .A1 (n_5235), .B0 (n_4696), .Y (n_4798));
OAI21X1 g57523(.A0 (n_4674), .A1 (n_4127), .B0 (n_5460), .Y (n_4797));
OAI21X1 g57532(.A0 (n_4605), .A1 (n_6660), .B0 (n_5566), .Y (n_4796));
OAI21X1 g57538(.A0 (n_4671), .A1 (n_4634), .B0 (n_5566), .Y (n_4795));
OAI21X1 g57547(.A0 (n_4485), .A1 (n_6201), .B0 (n_4947), .Y (n_4794));
OAI21X1 g57592(.A0 (n_4426), .A1 (n_6668), .B0 (n_4947), .Y (n_4793));
OAI21X1 g56723(.A0 (n_4454), .A1 (n_5729), .B0 (n_4685), .Y (n_4792));
OAI21X1 g56726(.A0 (n_4125), .A1 (n_5439), .B0 (n_4684), .Y (n_4791));
INVX1 g55805(.A (DATA_9_30), .Y (n_4790));
NOR2X1 g56759(.A (WX5715), .B (n_1425), .Y (n_4788));
NOR2X1 g56762(.A (WX5715), .B (n_5427), .Y (n_4786));
OAI21X1 g56781(.A0 (n_4540), .A1 (n_4803), .B0 (n_4419), .Y (n_4785));
OAI21X1 g56784(.A0 (n_4390), .A1 (n_5750), .B0 (n_4683), .Y (n_4784));
OAI21X1 g56785(.A0 (n_4367), .A1 (n_5750), .B0 (n_4388), .Y (n_4783));
NOR2X1 g56801(.A (WX7008), .B (n_5427), .Y (n_9438));
NOR2X1 g56824(.A (WX7008), .B (n_2851), .Y (n_4781));
OAI21X1 g56838(.A0 (n_4638), .A1 (n_5535), .B0 (n_4682), .Y (n_4780));
OAI21X1 g56840(.A0 (n_4528), .A1 (n_5535), .B0 (n_4681), .Y (n_4779));
OAI21X1 g56842(.A0 (n_4446), .A1 (n_4803), .B0 (n_4680), .Y (n_4778));
NOR2X1 g56862(.A (WX8301), .B (n_5712), .Y (n_4777));
NOR2X1 g56865(.A (WX8301), .B (n_5479), .Y (n_4775));
OAI21X1 g56897(.A0 (n_4277), .A1 (n_5393), .B0 (n_4753), .Y (n_4774));
OAI21X1 g56900(.A0 (n_4444), .A1 (n_5535), .B0 (n_4752), .Y (n_4773));
OAI21X1 g56902(.A0 (n_4385), .A1 (n_5468), .B0 (n_4751), .Y (n_4772));
OAI21X1 g56930(.A0 (n_4332), .A1 (n_4559), .B0 (n_4947), .Y (n_4771));
OAI21X1 g56958(.A0 (n_4257), .A1 (n_5196), .B0 (n_4678), .Y (n_4770));
OAI21X1 g55846(.A0 (n_4178), .A1 (n_5843), .B0 (n_4037), .Y(DATA_9_29));
NOR2X1 g58163(.A (WX10887), .B (n_5712), .Y (n_4769));
NOR2X1 g58164(.A (WX1836), .B (n_1648), .Y (n_4768));
OAI21X1 g57016(.A0 (n_4088), .A1 (n_5439), .B0 (n_4660), .Y (n_4766));
NOR2X1 g58172(.A (WX1836), .B (n_4882), .Y (n_4765));
NOR2X1 g58176(.A (WX10887), .B (n_6438), .Y (n_7509));
DFFSRX1 WX543_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4657), .Q (WX543), .QN ());
OAI21X1 g57332(.A0 (n_4328), .A1 (n_5242), .B0 (n_4086), .Y(DATA_9_31));
OAI21X1 g55803(.A0 (n_3842), .A1 (n_5183), .B0 (n_4658), .Y (n_4762));
OAI21X1 g56630(.A0 (n_4327), .A1 (n_10721), .B0 (n_5556), .Y(n_4761));
OAI21X1 g57505(.A0 (n_3806), .A1 (n_4803), .B0 (n_4648), .Y (n_4760));
OAI21X1 g57515(.A0 (n_4109), .A1 (n_6091), .B0 (n_4047), .Y(DATA_9_0));
DFFSRX1 WX8257_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4676), .Q (), .QN (WX8257));
DFFSRX1 WX9548_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4673), .Q (), .QN (WX9548));
DFFSRX1 WX4384_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4672), .Q (), .QN (WX4384));
DFFSRX1 WX5675_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4669), .Q (), .QN (WX5675));
DFFSRX1 WX6966_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4667), .Q (), .QN (WX6966));
DFFSRX1 WX3093_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4665), .Q (), .QN (WX3093));
OAI21X1 g55806(.A0 (n_4334), .A1 (n_5242), .B0 (n_4031), .Y(DATA_9_30));
NOR2X1 g56751(.A (WX4424), .B (n_5712), .Y (n_4759));
NOR2X1 g56754(.A (WX4424), .B (n_5838), .Y (n_4758));
OAI21X1 g55796(.A0 (n_4295), .A1 (n_5183), .B0 (n_4659), .Y (n_4757));
OAI21X1 g56763(.A0 (n_4455), .A1 (n_6684), .B0 (n_5722), .Y (n_4756));
OAI21X1 g56802(.A0 (n_4126), .A1 (n_11604), .B0 (n_5275), .Y(n_4755));
OAI21X1 g56866(.A0 (n_4335), .A1 (n_4639), .B0 (n_5722), .Y (n_4754));
OAI21X1 g56924(.A0 (n_3845), .A1 (n_9419), .B0 (n_6497), .Y (n_4753));
OAI21X1 g56934(.A0 (n_4527), .A1 (n_6202), .B0 (n_5460), .Y (n_4752));
OAI21X1 g56942(.A0 (n_6886), .A1 (n_6213), .B0 (n_4947), .Y (n_4751));
DFFSRX1 WX9594_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4333), .Q (), .QN (WX9594));
OAI21X1 g56979(.A0 (n_4384), .A1 (n_6183), .B0 (n_4947), .Y (n_4750));
OAI21X1 g57001(.A0 (n_3639), .A1 (n_6451), .B0 (n_5566), .Y (n_4749));
OAI21X1 g57039(.A0 (n_4382), .A1 (n_6670), .B0 (n_5460), .Y (n_4748));
OAI21X1 g57104(.A0 (n_4617), .A1 (n_6203), .B0 (n_4860), .Y (n_4747));
OAI21X1 g57329(.A0 (n_3843), .A1 (n_5105), .B0 (n_4331), .Y (n_4746));
OR2X1 g57366(.A (n_4330), .B (n_4697), .Y (n_4745));
OAI21X1 g57519(.A0 (n_3447), .A1 (n_4459), .B0 (n_4947), .Y (n_4744));
DFFSRX1 WX3129_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4320), .Q (), .QN (WX3129));
OAI21X1 g57520(.A0 (n_3433), .A1 (n_4451), .B0 (n_5619), .Y (n_4743));
OAI21X1 g57525(.A0 (n_4372), .A1 (n_6662), .B0 (n_5460), .Y (n_4742));
OAI21X1 g57527(.A0 (n_4370), .A1 (n_6663), .B0 (n_5460), .Y (n_4741));
OAI21X1 g57528(.A0 (n_3601), .A1 (n_4368), .B0 (n_5556), .Y (n_4740));
OAI21X1 g57533(.A0 (n_3850), .A1 (n_4602), .B0 (n_4860), .Y (n_4739));
OAI21X1 g57534(.A0 (n_4599), .A1 (n_6204), .B0 (n_3183), .Y (n_4738));
OAI21X1 g57535(.A0 (n_4597), .A1 (n_6661), .B0 (n_4860), .Y (n_4737));
OAI21X1 g57539(.A0 (n_3857), .A1 (n_6632), .B0 (n_5460), .Y (n_4736));
OAI21X1 g57540(.A0 (n_4630), .A1 (n_6205), .B0 (n_5722), .Y (n_4735));
OAI21X1 g57542(.A0 (n_3434), .A1 (n_4627), .B0 (n_5566), .Y (n_4734));
OAI21X1 g57549(.A0 (n_4483), .A1 (n_6206), .B0 (n_6479), .Y (n_4733));
OAI21X1 g57550(.A0 (n_4481), .A1 (n_6208), .B0 (n_4860), .Y (n_4731));
OAI21X1 g57553(.A0 (n_4090), .A1 (n_4135), .B0 (n_5722), .Y (n_4730));
OR2X1 g57554(.A (n_4199), .B (n_4697), .Y (n_4729));
OR2X1 g57555(.A (n_4197), .B (n_4697), .Y (n_4728));
OR2X1 g57556(.A (n_4194), .B (n_4697), .Y (n_4727));
OR2X1 g57557(.A (n_4192), .B (n_4697), .Y (n_4725));
OR2X1 g57558(.A (n_4190), .B (n_4697), .Y (n_4723));
OR2X1 g57559(.A (n_4187), .B (n_4697), .Y (n_4722));
OR2X1 g57560(.A (n_4185), .B (n_4697), .Y (n_4721));
OR2X1 g57561(.A (n_4182), .B (n_4697), .Y (n_4720));
OR2X1 g57563(.A (n_4180), .B (n_4697), .Y (n_4719));
OR2X1 g57564(.A (n_4177), .B (n_4697), .Y (n_4717));
OR2X1 g57565(.A (n_4175), .B (n_4697), .Y (n_4716));
OR2X1 g57566(.A (n_4173), .B (n_4697), .Y (n_4715));
OR2X1 g57567(.A (n_4171), .B (n_4697), .Y (n_4714));
OR2X1 g57568(.A (n_4169), .B (n_4697), .Y (n_15853));
OR2X1 g57569(.A (n_4167), .B (n_4697), .Y (n_4711));
OR2X1 g57572(.A (n_4161), .B (n_4697), .Y (n_4706));
OR2X1 g57573(.A (n_4159), .B (n_4697), .Y (n_4704));
OR2X1 g57575(.A (n_4155), .B (n_4697), .Y (n_4702));
OR2X1 g57579(.A (n_4146), .B (n_4697), .Y (n_4698));
OAI21X1 g56689(.A0 (n_3698), .A1 (n_4386), .B0 (n_5566), .Y (n_4696));
OR2X1 g57581(.A (n_4144), .B (n_4697), .Y (n_4695));
OR2X1 g57584(.A (n_4140), .B (n_4697), .Y (n_4693));
OR2X1 g57585(.A (n_4138), .B (n_4697), .Y (n_4692));
OR2X1 g57587(.A (n_4134), .B (n_4697), .Y (n_4690));
OAI21X1 g57593(.A0 (n_4422), .A1 (n_6207), .B0 (n_5460), .Y (n_4689));
OAI21X1 g57594(.A0 (n_4258), .A1 (n_7510), .B0 (n_5706), .Y (n_4688));
OAI21X1 g57595(.A0 (n_4420), .A1 (n_6677), .B0 (n_4947), .Y (n_4687));
OAI21X1 g57596(.A0 (n_4415), .A1 (n_6664), .B0 (n_5619), .Y (n_4686));
OAI21X1 g56755(.A0 (n_4083), .A1 (n_4566), .B0 (n_5566), .Y (n_4685));
OAI21X1 g56768(.A0 (n_4595), .A1 (n_6182), .B0 (n_4860), .Y (n_4684));
DFFSRX1 WX5715_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4221), .Q (), .QN (WX5715));
DFFSRX1 WX7008_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4108), .Q (), .QN (WX7008));
OAI21X1 g56821(.A0 (n_3689), .A1 (n_10723), .B0 (n_4860), .Y(n_4683));
OAI21X1 g56861(.A0 (n_3688), .A1 (n_4389), .B0 (n_4860), .Y (n_4682));
OAI21X1 g56870(.A0 (n_4366), .A1 (n_6669), .B0 (n_7087), .Y (n_4681));
OAI21X1 g56876(.A0 (n_4539), .A1 (n_6212), .B0 (n_5722), .Y (n_4680));
MX2X1 g57868(.A (n_4656), .B (WX545), .S0 (n_4050), .Y (n_4679));
DFFSRX1 WX8301_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4107), .Q (), .QN (WX8301));
OAI21X1 g56988(.A0 (n_4276), .A1 (n_8546), .B0 (n_4860), .Y (n_4678));
NOR2X1 g58159(.A (WX3095), .B (n_5662), .Y (n_4677));
NOR2X1 g58160(.A (WX8259), .B (n_1648), .Y (n_4676));
NOR2X1 g58161(.A (WX9550), .B (n_6438), .Y (n_6660));
NOR2X1 g58162(.A (WX8259), .B (n_4882), .Y (n_4674));
NOR2X1 g58165(.A (WX9550), .B (n_2851), .Y (n_4673));
NOR2X1 g58166(.A (WX4386), .B (n_2620), .Y (n_4672));
NOR2X1 g58168(.A (WX4386), .B (n_4670), .Y (n_4671));
NOR2X1 g58170(.A (WX5677), .B (n_1648), .Y (n_4669));
NOR2X1 g58171(.A (WX5677), .B (n_4670), .Y (n_6201));
NOR2X1 g58173(.A (WX6968), .B (n_1648), .Y (n_4667));
NOR2X1 g58175(.A (WX3095), .B (n_3690), .Y (n_4665));
NOR2X1 g58177(.A (WX6968), .B (n_6438), .Y (n_6668));
DFFSRX1 WX1836_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4093), .Q (), .QN (WX1836));
DFFSRX1 WX10887_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4092), .Q (), .QN (WX10887));
AOI21X1 g57785(.A0 (_2210_), .A1 (n_4608), .B0 (n_4661), .Y (n_4662));
OAI21X1 g57044(.A0 (n_3439), .A1 (n_4318), .B0 (n_6479), .Y (n_4660));
OAI21X1 g55817(.A0 (n_3437), .A1 (n_4198), .B0 (n_7087), .Y (n_4659));
OAI21X1 g55819(.A0 (n_3436), .A1 (n_4274), .B0 (n_6479), .Y (n_4658));
NOR2X1 g58609(.A (n_5181), .B (n_4656), .Y (n_4657));
OR2X1 g58614(.A (n_4656), .B (n_5990), .Y (n_4655));
AOI21X1 g57783(.A0 (_2212_), .A1 (n_4468), .B0 (n_4653), .Y (n_4654));
OAI21X1 g57353(.A0 (n_3435), .A1 (n_4329), .B0 (n_4860), .Y (n_4652));
OAI21X1 g57518(.A0 (n_3864), .A1 (n_4240), .B0 (n_4947), .Y (n_4651));
OAI21X1 g57548(.A0 (n_3855), .A1 (n_4254), .B0 (n_5722), .Y (n_4650));
OAI21X1 g57562(.A0 (n_3648), .A1 (n_4133), .B0 (n_4860), .Y (n_4649));
OAI21X1 g57597(.A0 (n_4256), .A1 (n_7511), .B0 (n_4947), .Y (n_4648));
AOI21X1 g57611(.A0 (_2163_), .A1 (n_4644), .B0 (n_4646), .Y (n_4647));
AOI21X1 g57613(.A0 (_2239_), .A1 (n_4644), .B0 (n_4643), .Y (n_4645));
AOI21X1 g57614(.A0 (_2162_), .A1 (n_4644), .B0 (n_4641), .Y (n_4642));
AOI21X1 g57615(.A0 (_2238_), .A1 (n_4562), .B0 (n_4639), .Y (n_4640));
AOI21X1 g57616(.A0 (_2237_), .A1 (n_4628), .B0 (n_9418), .Y (n_4638));
AOI21X1 g57617(.A0 (_2161_), .A1 (n_4562), .B0 (n_4634), .Y (n_4636));
AOI21X1 g57618(.A0 (_2160_), .A1 (n_4644), .B0 (n_6632), .Y (n_4633));
AOI21X1 g57619(.A0 (_2159_), .A1 (n_4644), .B0 (n_4630), .Y (n_4631));
AOI21X1 g57620(.A0 (_2158_), .A1 (n_4628), .B0 (n_4627), .Y (n_4629));
AOI21X1 g57621(.A0 (_2323_), .A1 (n_4628), .B0 (n_4625), .Y (n_4626));
AOI21X1 g57622(.A0 (_2157_), .A1 (n_4628), .B0 (n_4623), .Y (n_4624));
AOI21X1 g57623(.A0 (_2156_), .A1 (n_4562), .B0 (n_9404), .Y (n_4622));
AOI21X1 g57625(.A0 (_2154_), .A1 (n_4615), .B0 (n_9410), .Y (n_4620));
AOI21X1 g57627(.A0 (_2299_), .A1 (n_4603), .B0 (n_4617), .Y (n_4618));
AOI21X1 g57629(.A0 (_2298_), .A1 (n_4615), .B0 (n_4614), .Y (n_4616));
AOI21X1 g57630(.A0 (_2297_), .A1 (n_4615), .B0 (n_6508), .Y (n_4613));
AOI21X1 g57633(.A0 (_2295_), .A1 (n_4615), .B0 (n_4610), .Y (n_4611));
AOI21X1 g57635(.A0 (_2294_), .A1 (n_4608), .B0 (n_4607), .Y (n_4609));
AOI21X1 g57636(.A0 (_2293_), .A1 (n_4600), .B0 (n_4605), .Y (n_4606));
AOI21X1 g57638(.A0 (_2292_), .A1 (n_4603), .B0 (n_4602), .Y (n_4604));
AOI21X1 g57640(.A0 (_2291_), .A1 (n_4600), .B0 (n_4599), .Y (n_4601));
AOI21X1 g57641(.A0 (_2290_), .A1 (n_4593), .B0 (n_4597), .Y (n_4598));
AOI21X1 g57642(.A0 (_2140_), .A1 (n_4586), .B0 (n_4595), .Y (n_4596));
AOI21X1 g57644(.A0 (_2289_), .A1 (n_4593), .B0 (n_4592), .Y (n_4594));
AOI21X1 g57645(.A0 (_2288_), .A1 (n_4593), .B0 (n_4590), .Y (n_4591));
AOI21X1 g57646(.A0 (_2287_), .A1 (n_4615), .B0 (n_4588), .Y (n_4589));
AOI21X1 g57647(.A0 (_2147_), .A1 (n_4586), .B0 (n_9412), .Y (n_4587));
AOI21X1 g57650(.A0 (_2285_), .A1 (n_4600), .B0 (n_4583), .Y (n_4584));
AOI21X1 g57651(.A0 (_2284_), .A1 (n_4579), .B0 (n_4581), .Y (n_4582));
AOI21X1 g57652(.A0 (_2145_), .A1 (n_4579), .B0 (n_4578), .Y (n_4580));
AOI21X1 g57653(.A0 (_2283_), .A1 (n_4579), .B0 (n_9408), .Y (n_4577));
AOI21X1 g57654(.A0 (_2282_), .A1 (n_4615), .B0 (n_4574), .Y (n_4575));
AOI21X1 g57657(.A0 (_2280_), .A1 (n_4600), .B0 (n_4572), .Y (n_4573));
AOI21X1 g57660(.A0 (_2143_), .A1 (n_4579), .B0 (n_4570), .Y (n_4571));
AOI21X1 g57663(.A0 (_2142_), .A1 (n_4579), .B0 (n_4568), .Y (n_4569));
AOI21X1 g57667(.A0 (_2141_), .A1 (n_4603), .B0 (n_4566), .Y (n_4567));
AOI21X1 g57669(.A0 (_2273_), .A1 (n_4562), .B0 (n_4564), .Y (n_4565));
AOI21X1 g57670(.A0 (_2272_), .A1 (n_4562), .B0 (n_9416), .Y (n_4563));
AOI21X1 g57672(.A0 (_2270_), .A1 (n_4586), .B0 (n_4559), .Y (n_4560));
AOI21X1 g57673(.A0 (_2137_), .A1 (n_4579), .B0 (n_4557), .Y (n_4558));
AOI21X1 g57675(.A0 (_2136_), .A1 (n_4579), .B0 (n_4555), .Y (n_4556));
AOI21X1 g57676(.A0 (_2135_), .A1 (n_4579), .B0 (n_4553), .Y (n_4554));
AOI21X1 g57678(.A0 (_2330_), .A1 (n_4562), .B0 (n_4551), .Y (n_4552));
AOI21X1 g57680(.A0 (_2328_), .A1 (n_4593), .B0 (n_4547), .Y (n_4548));
AOI21X1 g57681(.A0 (_2327_), .A1 (n_4593), .B0 (n_4545), .Y (n_4546));
AOI21X1 g57682(.A0 (_2326_), .A1 (n_4593), .B0 (n_4543), .Y (n_4544));
AOI21X1 g57683(.A0 (_2325_), .A1 (n_4593), .B0 (n_4541), .Y (n_4542));
AOI21X1 g57684(.A0 (_2204_), .A1 (n_4586), .B0 (n_4539), .Y (n_4540));
AOI21X1 g57685(.A0 (_2324_), .A1 (n_4562), .B0 (n_4537), .Y (n_4538));
AOI21X1 g57686(.A0 (_2322_), .A1 (n_4562), .B0 (n_4535), .Y (n_4536));
AOI21X1 g57687(.A0 (_2321_), .A1 (n_4608), .B0 (n_4533), .Y (n_4534));
AOI21X1 g57688(.A0 (_2320_), .A1 (n_4608), .B0 (n_4531), .Y (n_4532));
AOI21X1 g57689(.A0 (_2319_), .A1 (n_4600), .B0 (n_4529), .Y (n_4530));
AOI21X1 g57691(.A0 (_2203_), .A1 (n_4608), .B0 (n_4527), .Y (n_4528));
AOI21X1 g57692(.A0 (_2317_), .A1 (n_4608), .B0 (n_4525), .Y (n_4526));
AOI21X1 g57694(.A0 (_2315_), .A1 (n_4562), .B0 (n_4523), .Y (n_4524));
AOI21X1 g57696(.A0 (_2134_), .A1 (n_4608), .B0 (n_4521), .Y (n_4522));
AOI21X1 g57698(.A0 (_2202_), .A1 (n_4600), .B0 (n_4519), .Y (n_4520));
AOI21X1 g57699(.A0 (_2312_), .A1 (n_4600), .B0 (n_4517), .Y (n_4518));
AOI21X1 g57700(.A0 (_2311_), .A1 (n_4600), .B0 (n_4515), .Y (n_4516));
AOI21X1 g57701(.A0 (_2310_), .A1 (n_4562), .B0 (n_4513), .Y (n_4514));
AOI21X1 g57702(.A0 (_2309_), .A1 (n_4562), .B0 (n_6488), .Y (n_4512));
AOI21X1 g57703(.A0 (_2308_), .A1 (n_4608), .B0 (n_4509), .Y (n_4510));
AOI21X1 g57704(.A0 (_2201_), .A1 (n_4608), .B0 (n_4507), .Y (n_4508));
AOI21X1 g57705(.A0 (_2307_), .A1 (n_4608), .B0 (n_4505), .Y (n_4506));
AOI21X1 g57708(.A0 (_2304_), .A1 (n_4628), .B0 (n_4503), .Y (n_4504));
AOI21X1 g57711(.A0 (_2200_), .A1 (n_4644), .B0 (n_4501), .Y (n_4502));
DFFSRX1 WX4424_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_4084), .Q (), .QN (WX4424));
AOI21X1 g57713(.A0 (_2199_), .A1 (n_4644), .B0 (n_4499), .Y (n_4500));
AOI21X1 g57714(.A0 (_2198_), .A1 (n_4562), .B0 (n_4497), .Y (n_4498));
AOI21X1 g57715(.A0 (_2133_), .A1 (n_4562), .B0 (n_4495), .Y (n_4496));
AOI21X1 g57716(.A0 (_2197_), .A1 (n_4628), .B0 (n_4493), .Y (n_4494));
AOI21X1 g57717(.A0 (_2196_), .A1 (n_4628), .B0 (n_4491), .Y (n_4492));
AOI21X1 g57718(.A0 (_2195_), .A1 (n_4644), .B0 (n_4489), .Y (n_4490));
AOI21X1 g57719(.A0 (_2132_), .A1 (n_4644), .B0 (n_4487), .Y (n_4488));
AOI21X1 g57720(.A0 (_2194_), .A1 (n_4562), .B0 (n_4485), .Y (n_4486));
AOI21X1 g57722(.A0 (_2192_), .A1 (n_4562), .B0 (n_4483), .Y (n_4484));
AOI21X1 g57723(.A0 (_2191_), .A1 (n_4644), .B0 (n_4481), .Y (n_4482));
AOI21X1 g57725(.A0 (_2190_), .A1 (n_4644), .B0 (n_4479), .Y (n_4480));
AOI21X1 g57726(.A0 (_2189_), .A1 (n_4644), .B0 (n_4477), .Y (n_4478));
AOI21X1 g57727(.A0 (_2188_), .A1 (n_4562), .B0 (n_9420), .Y (n_4476));
AOI21X1 g57732(.A0 (_2129_), .A1 (n_4471), .B0 (n_4473), .Y (n_4474));
AOI21X1 g57733(.A0 (_2184_), .A1 (n_4471), .B0 (n_9426), .Y (n_4472));
AOI21X1 g57735(.A0 (_2182_), .A1 (n_4468), .B0 (n_4467), .Y (n_4469));
AOI21X1 g57736(.A0 (_2181_), .A1 (n_4562), .B0 (n_4465), .Y (n_4466));
AOI21X1 g57737(.A0 (_2128_), .A1 (n_4603), .B0 (n_4463), .Y (n_4464));
AOI21X1 g57738(.A0 (_2180_), .A1 (n_4603), .B0 (n_4461), .Y (n_4462));
AOI21X1 g57744(.A0 (_2126_), .A1 (n_4468), .B0 (n_4459), .Y (n_4460));
AOI21X1 g57745(.A0 (_2175_), .A1 (n_4593), .B0 (n_4457), .Y (n_4458));
AOI21X1 g57746(.A0 (_2174_), .A1 (n_4593), .B0 (n_4455), .Y (n_4456));
AOI21X1 g57747(.A0 (_2173_), .A1 (n_4471), .B0 (n_10722), .Y(n_4454));
AOI21X1 g57748(.A0 (_2125_), .A1 (n_4471), .B0 (n_4451), .Y (n_4452));
AOI21X1 g57750(.A0 (_2123_), .A1 (n_4471), .B0 (n_4449), .Y (n_4450));
AOI21X1 g57751(.A0 (_2122_), .A1 (n_4586), .B0 (n_4447), .Y (n_4448));
AOI21X1 g57752(.A0 (_2236_), .A1 (n_4586), .B0 (n_6885), .Y (n_4446));
AOI21X1 g57753(.A0 (_2235_), .A1 (n_4586), .B0 (n_6451), .Y (n_4444));
AOI21X1 g57755(.A0 (_2234_), .A1 (n_4439), .B0 (n_4441), .Y (n_4442));
AOI21X1 g57756(.A0 (_2233_), .A1 (n_4439), .B0 (n_4438), .Y (n_4440));
AOI21X1 g57757(.A0 (_2232_), .A1 (n_4439), .B0 (n_4436), .Y (n_4437));
AOI21X1 g57759(.A0 (_2231_), .A1 (n_4586), .B0 (n_4434), .Y (n_4435));
AOI21X1 g57760(.A0 (_2230_), .A1 (n_4586), .B0 (n_4432), .Y (n_4433));
AOI21X1 g57761(.A0 (_2229_), .A1 (n_4586), .B0 (n_4430), .Y (n_4431));
AOI21X1 g57762(.A0 (_2228_), .A1 (n_4586), .B0 (n_4428), .Y (n_4429));
AOI21X1 g57763(.A0 (_2227_), .A1 (n_4603), .B0 (n_4426), .Y (n_4427));
AOI21X1 g57764(.A0 (_2119_), .A1 (n_4603), .B0 (n_4424), .Y (n_4425));
AOI21X1 g57765(.A0 (_2226_), .A1 (n_4586), .B0 (n_4422), .Y (n_4423));
AOI21X1 g57766(.A0 (_2225_), .A1 (n_4586), .B0 (n_4420), .Y (n_4421));
OAI21X1 g56810(.A0 (n_3642), .A1 (n_4124), .B0 (n_4860), .Y (n_4419));
AOI21X1 g57767(.A0 (_2118_), .A1 (n_4562), .B0 (n_4417), .Y (n_4418));
AOI21X1 g57768(.A0 (_2224_), .A1 (n_4562), .B0 (n_4415), .Y (n_4416));
AOI21X1 g57769(.A0 (_2223_), .A1 (n_4603), .B0 (n_4413), .Y (n_4414));
AOI21X1 g57770(.A0 (_2222_), .A1 (n_4439), .B0 (n_4411), .Y (n_4412));
AOI21X1 g57771(.A0 (_2221_), .A1 (n_4603), .B0 (n_4409), .Y (n_4410));
AOI21X1 g57772(.A0 (_2220_), .A1 (n_4439), .B0 (n_9422), .Y (n_4408));
AOI21X1 g57774(.A0 (_2219_), .A1 (n_4468), .B0 (n_4405), .Y (n_4406));
AOI21X1 g57775(.A0 (_2218_), .A1 (n_4471), .B0 (n_4403), .Y (n_4404));
AOI21X1 g57777(.A0 (_2217_), .A1 (n_4439), .B0 (n_4401), .Y (n_4402));
AOI21X1 g57778(.A0 (_2216_), .A1 (n_4439), .B0 (n_4399), .Y (n_4400));
AOI21X1 g57781(.A0 (_2115_), .A1 (n_4439), .B0 (n_9414), .Y (n_4398));
AOI21X1 g57782(.A0 (_2213_), .A1 (n_4562), .B0 (n_4395), .Y (n_4396));
AOI21X1 g57788(.A0 (_2113_), .A1 (n_4468), .B0 (n_10714), .Y(n_4394));
AOI21X1 g57789(.A0 (_2208_), .A1 (n_4468), .B0 (n_10718), .Y(n_4392));
AOI21X1 g57792(.A0 (_2205_), .A1 (n_4600), .B0 (n_4389), .Y (n_4390));
OAI21X1 g56827(.A0 (n_3443), .A1 (n_4294), .B0 (n_4860), .Y (n_4388));
AOI21X1 g57800(.A0 (_2109_), .A1 (n_4471), .B0 (n_4386), .Y (n_4387));
AOI21X1 g57828(.A0 (_2268_), .A1 (n_4586), .B0 (n_4384), .Y (n_4385));
AOI21X1 g57829(.A0 (_2267_), .A1 (n_4603), .B0 (n_4382), .Y (n_4383));
AOI21X1 g57830(.A0 (_2266_), .A1 (n_4471), .B0 (n_4380), .Y (n_4381));
AOI21X1 g57831(.A0 (_2265_), .A1 (n_4468), .B0 (n_4378), .Y (n_4379));
AOI21X1 g57832(.A0 (_2264_), .A1 (n_4603), .B0 (n_4376), .Y (n_4377));
AOI21X1 g57833(.A0 (_2263_), .A1 (n_4468), .B0 (n_4374), .Y (n_4375));
AOI21X1 g57837(.A0 (_2259_), .A1 (n_4603), .B0 (n_4372), .Y (n_4373));
AOI21X1 g57839(.A0 (_2258_), .A1 (n_4644), .B0 (n_4370), .Y (n_4371));
AOI21X1 g57840(.A0 (_2257_), .A1 (n_4628), .B0 (n_4368), .Y (n_4369));
AOI21X1 g57841(.A0 (_2171_), .A1 (n_4628), .B0 (n_4366), .Y (n_4367));
AOI21X1 g57842(.A0 (_2256_), .A1 (n_4628), .B0 (n_4364), .Y (n_4365));
AOI21X1 g57843(.A0 (_2255_), .A1 (n_4562), .B0 (n_4362), .Y (n_4363));
AOI21X1 g57844(.A0 (_2254_), .A1 (n_4628), .B0 (n_4360), .Y (n_4361));
AOI21X1 g57845(.A0 (_2170_), .A1 (n_4593), .B0 (n_4358), .Y (n_4359));
AOI21X1 g57846(.A0 (_2253_), .A1 (n_4593), .B0 (n_4356), .Y (n_4357));
AOI21X1 g57847(.A0 (_2169_), .A1 (n_4579), .B0 (n_4354), .Y (n_4355));
AOI21X1 g57849(.A0 (_2251_), .A1 (n_4593), .B0 (n_9406), .Y (n_4353));
AOI21X1 g57850(.A0 (_2168_), .A1 (n_4615), .B0 (n_4350), .Y (n_4351));
AOI21X1 g57852(.A0 (_2249_), .A1 (n_4615), .B0 (n_4348), .Y (n_4349));
AOI21X1 g57853(.A0 (_2167_), .A1 (n_4615), .B0 (n_4346), .Y (n_4347));
AOI21X1 g57855(.A0 (_2247_), .A1 (n_4468), .B0 (n_9428), .Y (n_4345));
AOI21X1 g57856(.A0 (_2166_), .A1 (n_4468), .B0 (n_4342), .Y (n_4343));
AOI21X1 g57858(.A0 (_2245_), .A1 (n_4468), .B0 (n_4340), .Y (n_4341));
AOI21X1 g57859(.A0 (_2165_), .A1 (n_4628), .B0 (n_4338), .Y (n_4339));
AOI21X1 g57862(.A0 (_2164_), .A1 (n_4628), .B0 (n_4336), .Y (n_4337));
NOR2X1 g56923(.A (WX8303), .B (n_5479), .Y (n_4335));
MX2X1 g55844(.A (n_2888), .B (WX487), .S0 (n_10747), .Y (n_4334));
NOR2X1 g56984(.A (WX9596), .B (n_1425), .Y (n_4333));
NOR2X1 g56987(.A (WX9596), .B (n_5479), .Y (n_4332));
OAI21X1 g57352(.A0 (n_3431), .A1 (n_4087), .B0 (n_4860), .Y (n_4331));
AOI21X1 g57394(.A0 (_2108_), .A1 (n_4184), .B0 (n_4329), .Y (n_4330));
MX2X1 g57401(.A (n_3599), .B (WX485), .S0 (n_9433), .Y (n_4328));
NOR2X1 g56688(.A (WX3131), .B (n_4670), .Y (n_4327));
AOI21X1 g57610(.A0 (_2241_), .A1 (n_4644), .B0 (n_4325), .Y (n_4326));
AOI21X1 g57612(.A0 (_2240_), .A1 (n_4644), .B0 (n_4323), .Y (n_4324));
AOI21X1 g57624(.A0 (_2155_), .A1 (n_4615), .B0 (n_11605), .Y(n_4322));
NOR2X1 g56709(.A (WX3131), .B (n_3690), .Y (n_4320));
AOI21X1 g57626(.A0 (_2300_), .A1 (n_4562), .B0 (n_4318), .Y (n_4319));
AOI21X1 g57628(.A0 (_2153_), .A1 (n_4615), .B0 (n_4316), .Y (n_4317));
AOI21X1 g57631(.A0 (_2152_), .A1 (n_4603), .B0 (n_4314), .Y (n_4315));
AOI21X1 g57632(.A0 (_2296_), .A1 (n_4615), .B0 (n_4312), .Y (n_4313));
AOI21X1 g57634(.A0 (_2151_), .A1 (n_4615), .B0 (n_4310), .Y (n_4311));
AOI21X1 g57637(.A0 (_2150_), .A1 (n_4600), .B0 (n_4308), .Y (n_4309));
AOI21X1 g57639(.A0 (_2149_), .A1 (n_4600), .B0 (n_11619), .Y(n_4307));
AOI21X1 g57643(.A0 (_2148_), .A1 (n_4593), .B0 (n_4304), .Y (n_4305));
AOI21X1 g57648(.A0 (_2286_), .A1 (n_4615), .B0 (n_4302), .Y (n_4303));
AOI21X1 g57649(.A0 (_2146_), .A1 (n_4600), .B0 (n_11623), .Y(n_4301));
AOI21X1 g57655(.A0 (_2281_), .A1 (n_4615), .B0 (n_4298), .Y (n_4299));
AOI21X1 g57656(.A0 (_2144_), .A1 (n_4600), .B0 (n_11597), .Y(n_4297));
AOI21X1 g57658(.A0 (_2139_), .A1 (n_4579), .B0 (n_4294), .Y (n_4295));
AOI21X1 g57659(.A0 (_2279_), .A1 (n_4579), .B0 (n_4292), .Y (n_4293));
AOI21X1 g57661(.A0 (_2278_), .A1 (n_4579), .B0 (n_4290), .Y (n_4291));
AOI21X1 g57662(.A0 (_2277_), .A1 (n_4579), .B0 (n_4288), .Y (n_4289));
AOI21X1 g57664(.A0 (_2276_), .A1 (n_4579), .B0 (n_4286), .Y (n_4287));
AOI21X1 g57665(.A0 (_2275_), .A1 (n_4579), .B0 (n_11596), .Y(n_4285));
AOI21X1 g57666(.A0 (_2138_), .A1 (n_4603), .B0 (n_4282), .Y (n_4283));
AOI21X1 g57668(.A0 (_2274_), .A1 (n_4603), .B0 (n_4280), .Y (n_4281));
AOI21X1 g57671(.A0 (_2271_), .A1 (n_4586), .B0 (n_11601), .Y(n_4279));
AOI21X1 g57674(.A0 (_2269_), .A1 (n_4579), .B0 (n_4276), .Y (n_4277));
AOI21X1 g57677(.A0 (_2331_), .A1 (n_4562), .B0 (n_4274), .Y (n_4275));
AOI21X1 g57690(.A0 (_2318_), .A1 (n_4600), .B0 (n_4272), .Y (n_4273));
AOI21X1 g57693(.A0 (_2316_), .A1 (n_4562), .B0 (n_7084), .Y (n_4271));
AOI21X1 g57695(.A0 (_2314_), .A1 (n_4608), .B0 (n_6469), .Y (n_4269));
AOI21X1 g57697(.A0 (_2313_), .A1 (n_4600), .B0 (n_4266), .Y (n_4267));
AOI21X1 g57706(.A0 (_2306_), .A1 (n_4608), .B0 (n_4264), .Y (n_4265));
AOI21X1 g57707(.A0 (_2305_), .A1 (n_4628), .B0 (n_4262), .Y (n_4263));
AOI21X1 g57709(.A0 (_2303_), .A1 (n_4562), .B0 (n_4260), .Y (n_4261));
AOI21X1 g57710(.A0 (_2302_), .A1 (n_4562), .B0 (n_4258), .Y (n_4259));
AOI21X1 g57712(.A0 (_2301_), .A1 (n_4593), .B0 (n_4256), .Y (n_4257));
AOI21X1 g57721(.A0 (_2193_), .A1 (n_4562), .B0 (n_4254), .Y (n_4255));
AOI21X1 g57724(.A0 (_2131_), .A1 (n_4644), .B0 (n_4252), .Y (n_4253));
AOI21X1 g57728(.A0 (_2130_), .A1 (n_4562), .B0 (n_4250), .Y (n_4251));
AOI21X1 g57729(.A0 (_2187_), .A1 (n_4468), .B0 (n_4248), .Y (n_4249));
AOI21X1 g57730(.A0 (_2186_), .A1 (n_4608), .B0 (n_11607), .Y(n_4247));
AOI21X1 g57731(.A0 (_2185_), .A1 (n_4608), .B0 (n_4244), .Y (n_4245));
AOI21X1 g57734(.A0 (_2183_), .A1 (n_4468), .B0 (n_11615), .Y(n_4243));
AOI21X1 g57739(.A0 (_2127_), .A1 (n_4471), .B0 (n_4240), .Y (n_4241));
AOI21X1 g57740(.A0 (_2179_), .A1 (n_4471), .B0 (n_4238), .Y (n_4239));
AOI21X1 g57741(.A0 (_2178_), .A1 (n_4439), .B0 (n_4236), .Y (n_4237));
AOI21X1 g57742(.A0 (_2177_), .A1 (n_4439), .B0 (n_10716), .Y(n_4235));
AOI21X1 g57743(.A0 (_2176_), .A1 (n_4593), .B0 (n_4232), .Y (n_4233));
AOI21X1 g57749(.A0 (_2124_), .A1 (n_4471), .B0 (n_4230), .Y (n_4231));
AOI21X1 g57754(.A0 (_2121_), .A1 (n_4439), .B0 (n_4228), .Y (n_4229));
AOI21X1 g57758(.A0 (_2120_), .A1 (n_4439), .B0 (n_11611), .Y(n_4227));
AOI21X1 g57773(.A0 (_2117_), .A1 (n_4439), .B0 (n_4224), .Y (n_4225));
AOI21X1 g57776(.A0 (_2116_), .A1 (n_4439), .B0 (n_4222), .Y (n_4223));
NOR2X1 g56817(.A (WX5717), .B (n_2620), .Y (n_4221));
AOI21X1 g57779(.A0 (_2215_), .A1 (n_4439), .B0 (n_4219), .Y (n_4220));
AOI21X1 g57780(.A0 (_2214_), .A1 (n_4439), .B0 (n_11617), .Y(n_4218));
NOR2X1 g56820(.A (WX5717), .B (n_5052), .Y (n_6684));
AOI21X1 g57784(.A0 (_2211_), .A1 (n_4468), .B0 (n_11621), .Y(n_4215));
AOI21X1 g57786(.A0 (_2114_), .A1 (n_4468), .B0 (n_11625), .Y(n_4213));
AOI21X1 g57787(.A0 (_2209_), .A1 (n_4608), .B0 (n_4210), .Y (n_4211));
AOI21X1 g57790(.A0 (_2207_), .A1 (n_4562), .B0 (n_4208), .Y (n_4209));
AOI21X1 g57791(.A0 (_2206_), .A1 (n_4600), .B0 (n_11603), .Y(n_4207));
AOI21X1 g57793(.A0 (_2112_), .A1 (n_4471), .B0 (n_4204), .Y (n_4205));
AOI21X1 g57794(.A0 (_2111_), .A1 (n_4471), .B0 (n_11599), .Y(n_4203));
AOI21X1 g57795(.A0 (_2110_), .A1 (n_4471), .B0 (n_10720), .Y(n_4201));
AOI21X1 g57796(.A0 (_2107_), .A1 (n_3831), .B0 (n_4198), .Y (n_4199));
AOI21X1 g57797(.A0 (_2106_), .A1 (n_3831), .B0 (n_4195), .Y (n_4197));
AOI21X1 g57798(.A0 (_2105_), .A1 (n_3831), .B0 (n_4193), .Y (n_4194));
AOI21X1 g57799(.A0 (_2104_), .A1 (n_5828), .B0 (n_4191), .Y (n_4192));
AOI21X1 g57801(.A0 (_2103_), .A1 (n_5828), .B0 (n_4188), .Y (n_4190));
AOI21X1 g57802(.A0 (_2102_), .A1 (n_3831), .B0 (n_4186), .Y (n_4187));
AOI21X1 g57803(.A0 (_2101_), .A1 (n_4184), .B0 (n_4183), .Y (n_4185));
AOI21X1 g57804(.A0 (_2100_), .A1 (n_5828), .B0 (n_4181), .Y (n_4182));
AOI21X1 g57805(.A0 (_2099_), .A1 (n_4184), .B0 (n_4179), .Y (n_4180));
MX2X1 g55904(.A (n_3685), .B (WX489), .S0 (n_7082), .Y (n_4178));
AOI21X1 g57806(.A0 (_2098_), .A1 (n_4184), .B0 (n_4176), .Y (n_4177));
AOI21X1 g57807(.A0 (_2097_), .A1 (n_4150), .B0 (n_4174), .Y (n_4175));
AOI21X1 g57808(.A0 (_2096_), .A1 (n_4184), .B0 (n_4172), .Y (n_4173));
AOI21X1 g57809(.A0 (_2095_), .A1 (n_4184), .B0 (n_4170), .Y (n_4171));
AOI21X1 g57810(.A0 (_2094_), .A1 (n_5828), .B0 (n_4168), .Y (n_4169));
AOI21X1 g57811(.A0 (_2093_), .A1 (n_4184), .B0 (n_4166), .Y (n_4167));
AOI21X1 g57812(.A0 (_2092_), .A1 (n_5828), .B0 (n_4164), .Y (n_4165));
AOI21X1 g57813(.A0 (_2091_), .A1 (n_5828), .B0 (n_4162), .Y (n_4163));
AOI21X1 g57814(.A0 (_2090_), .A1 (n_4184), .B0 (n_4160), .Y (n_4161));
AOI21X1 g57815(.A0 (_2089_), .A1 (n_5828), .B0 (n_4158), .Y (n_4159));
AOI21X1 g57816(.A0 (_2088_), .A1 (n_4184), .B0 (n_4156), .Y (n_4157));
AOI21X1 g57817(.A0 (_2087_), .A1 (n_4184), .B0 (n_4154), .Y (n_4155));
AOI21X1 g57818(.A0 (_2086_), .A1 (n_5828), .B0 (n_4152), .Y (n_4153));
AOI21X1 g57819(.A0 (_2085_), .A1 (n_4150), .B0 (n_4149), .Y (n_4151));
AOI21X1 g57820(.A0 (_2084_), .A1 (n_5828), .B0 (n_4147), .Y (n_4148));
AOI21X1 g57821(.A0 (_2083_), .A1 (n_3831), .B0 (n_4145), .Y (n_4146));
AOI21X1 g57822(.A0 (_2082_), .A1 (n_5828), .B0 (n_4143), .Y (n_4144));
AOI21X1 g57823(.A0 (_2081_), .A1 (n_5828), .B0 (n_4141), .Y (n_4142));
AOI21X1 g57824(.A0 (_2080_), .A1 (n_4184), .B0 (n_4139), .Y (n_4140));
AOI21X1 g57825(.A0 (_2079_), .A1 (n_4184), .B0 (n_4137), .Y (n_4138));
AOI21X1 g57826(.A0 (_2078_), .A1 (n_4150), .B0 (n_4135), .Y (n_4136));
AOI21X1 g57827(.A0 (_2077_), .A1 (n_5828), .B0 (n_4133), .Y (n_4134));
AOI21X1 g57834(.A0 (_2262_), .A1 (n_4608), .B0 (n_4131), .Y (n_4132));
AOI21X1 g57835(.A0 (_2261_), .A1 (n_4471), .B0 (n_4129), .Y (n_4130));
AOI21X1 g57836(.A0 (_2260_), .A1 (n_4471), .B0 (n_4127), .Y (n_4128));
NOR2X1 g56860(.A (WX7010), .B (n_5479), .Y (n_4126));
AOI21X1 g57838(.A0 (_2172_), .A1 (n_4562), .B0 (n_4124), .Y (n_4125));
AOI21X1 g57848(.A0 (_2252_), .A1 (n_4593), .B0 (n_4122), .Y (n_4123));
AOI21X1 g57851(.A0 (_2250_), .A1 (n_4603), .B0 (n_11609), .Y(n_4121));
AOI21X1 g57854(.A0 (_2248_), .A1 (n_4615), .B0 (n_11613), .Y(n_4119));
AOI21X1 g57857(.A0 (_2246_), .A1 (n_4468), .B0 (n_4116), .Y (n_4117));
AOI21X1 g57860(.A0 (_2244_), .A1 (n_4628), .B0 (n_4114), .Y (n_4115));
AOI21X1 g57861(.A0 (_2243_), .A1 (n_4628), .B0 (n_4112), .Y (n_4113));
AOI21X1 g57863(.A0 (_2242_), .A1 (n_4562), .B0 (n_10712), .Y(n_4111));
MX2X1 g57869(.A (n_3695), .B (WX547), .S0 (n_9437), .Y (n_4109));
NOR2X1 g56883(.A (WX7010), .B (n_2851), .Y (n_4108));
NOR2X1 g56920(.A (WX8303), .B (n_1648), .Y (n_4107));
AND2X1 g57963(.A (n_3980), .B (n_4106), .Y (n_4566));
AND2X1 g57965(.A (n_3979), .B (n_4106), .Y (n_4564));
AND2X1 g57969(.A (n_3977), .B (n_4105), .Y (n_4559));
AND2X1 g57970(.A (n_3976), .B (n_4105), .Y (n_4557));
AND2X1 g57972(.A (n_3975), .B (n_4101), .Y (n_4551));
AND2X1 g57975(.A (n_3974), .B (n_4103), .Y (n_4549));
AND2X1 g57976(.A (n_3973), .B (n_4104), .Y (n_4555));
AND2X1 g57977(.A (n_3972), .B (n_4105), .Y (n_4553));
AND2X1 g57978(.A (n_3971), .B (n_4106), .Y (n_4539));
AND2X1 g57980(.A (n_3970), .B (n_4104), .Y (n_4547));
AND2X1 g57981(.A (n_3969), .B (n_4105), .Y (n_4527));
AND2X1 g57982(.A (n_3968), .B (n_4106), .Y (n_4521));
AND2X1 g57983(.A (n_3967), .B (n_4103), .Y (n_4519));
AND2X1 g57984(.A (n_3966), .B (n_4096), .Y (n_4507));
AND2X1 g57986(.A (n_3965), .B (n_4104), .Y (n_4501));
AND2X1 g57987(.A (n_3964), .B (n_4104), .Y (n_4545));
AND2X1 g57988(.A (n_3963), .B (n_4104), .Y (n_4499));
AND2X1 g57990(.A (n_3962), .B (n_4106), .Y (n_4497));
AND2X1 g57991(.A (n_3961), .B (n_4100), .Y (n_4495));
AND2X1 g57992(.A (n_3960), .B (n_4103), .Y (n_4493));
AND2X1 g57993(.A (n_3959), .B (n_4096), .Y (n_4491));
AND2X1 g57995(.A (n_3957), .B (n_6452), .Y (n_4543));
AND2X1 g57996(.A (n_3958), .B (n_4101), .Y (n_4489));
AND2X1 g57997(.A (n_3956), .B (n_4101), .Y (n_4487));
AND2X1 g57998(.A (n_3955), .B (n_4100), .Y (n_4485));
AND2X1 g58001(.A (n_3954), .B (n_6633), .Y (n_4483));
AND2X1 g58002(.A (n_3953), .B (n_4099), .Y (n_4541));
AND2X1 g58003(.A (n_3952), .B (n_4099), .Y (n_4481));
AND2X1 g58005(.A (n_3951), .B (n_4096), .Y (n_4479));
AND2X1 g58007(.A (n_4099), .B (n_7281), .Y (n_4477));
AND2X1 g58011(.A (n_3948), .B (n_6452), .Y (n_4537));
AND2X1 g58015(.A (n_3947), .B (n_4101), .Y (n_4473));
AND2X1 g58018(.A (n_3945), .B (n_4099), .Y (n_4625));
AND2X1 g58020(.A (n_3944), .B (n_6452), .Y (n_4467));
AND2X1 g58021(.A (n_3943), .B (n_4099), .Y (n_4465));
AND2X1 g58022(.A (n_3942), .B (n_4106), .Y (n_4463));
AND2X1 g58023(.A (n_3941), .B (n_4104), .Y (n_4461));
AND2X1 g58027(.A (n_3940), .B (n_4106), .Y (n_4535));
AND2X1 g58031(.A (n_3939), .B (n_6633), .Y (n_4459));
AND2X1 g58032(.A (n_3938), .B (n_6452), .Y (n_4457));
AND2X1 g58033(.A (n_3937), .B (n_4099), .Y (n_4533));
AND2X1 g58035(.A (n_3936), .B (n_4096), .Y (n_4455));
AND2X1 g58038(.A (n_3934), .B (n_4106), .Y (n_4451));
AND2X1 g58039(.A (n_3933), .B (n_4095), .Y (n_4531));
AND2X1 g58042(.A (n_3932), .B (n_4099), .Y (n_4529));
AND2X1 g58044(.A (n_4103), .B (n_8340), .Y (n_4449));
AND2X1 g58047(.A (n_3930), .B (n_6452), .Y (n_4447));
AND2X1 g58051(.A (n_3927), .B (n_4100), .Y (n_4441));
AND2X1 g58052(.A (n_3926), .B (n_4100), .Y (n_4438));
AND2X1 g58053(.A (n_3925), .B (n_4096), .Y (n_4525));
AND2X1 g58055(.A (n_3924), .B (n_4100), .Y (n_4436));
AND2X1 g58057(.A (n_3923), .B (n_4096), .Y (n_4434));
AND2X1 g58058(.A (n_3922), .B (n_4100), .Y (n_4432));
AND2X1 g58060(.A (n_3921), .B (n_4100), .Y (n_4430));
AND2X1 g58062(.A (n_3920), .B (n_4096), .Y (n_4428));
AND2X1 g58064(.A (n_3919), .B (n_6452), .Y (n_4426));
AND2X1 g58065(.A (n_6633), .B (n_8346), .Y (n_4424));
AND2X1 g58066(.A (n_3917), .B (n_4105), .Y (n_4422));
AND2X1 g58067(.A (n_3916), .B (n_6633), .Y (n_4420));
AND2X1 g58068(.A (n_3915), .B (n_4105), .Y (n_4523));
AND2X1 g58069(.A (n_3913), .B (n_4095), .Y (n_4417));
AND2X1 g58070(.A (n_3914), .B (n_4099), .Y (n_4415));
AND2X1 g58072(.A (n_3912), .B (n_4095), .Y (n_4413));
AND2X1 g58073(.A (n_3911), .B (n_4104), .Y (n_4411));
AND2X1 g58075(.A (n_3910), .B (n_6633), .Y (n_4409));
AND2X1 g58079(.A (n_3908), .B (n_4104), .Y (n_4405));
AND2X1 g58080(.A (n_4095), .B (n_8341), .Y (n_4403));
AND2X1 g58082(.A (n_3906), .B (n_4095), .Y (n_4401));
AND2X1 g58085(.A (n_4100), .B (n_8344), .Y (n_4399));
AND2X1 g58089(.A (n_3903), .B (n_6452), .Y (n_4395));
AND2X1 g58091(.A (n_3901), .B (n_4100), .Y (n_4517));
AND2X1 g58092(.A (n_6633), .B (n_8349), .Y (n_4653));
AND2X1 g58095(.A (n_3900), .B (n_4101), .Y (n_4661));
AND2X1 g58098(.A (n_3898), .B (n_4017), .Y (n_4515));
AND2X1 g58104(.A (n_4105), .B (n_9403), .Y (n_4389));
AND2X1 g58106(.A (n_3895), .B (n_6633), .Y (n_4513));
AND2X1 g58113(.A (n_3893), .B (n_4104), .Y (n_4509));
AND2X1 g58114(.A (n_3892), .B (n_4104), .Y (n_4386));
AND2X1 g58116(.A (n_3891), .B (n_4101), .Y (n_4505));
AND2X1 g58119(.A (n_3890), .B (n_6633), .Y (n_4384));
AND2X1 g58120(.A (n_3889), .B (n_4103), .Y (n_4382));
AND2X1 g58121(.A (n_3888), .B (n_4094), .Y (n_4380));
AND2X1 g58122(.A (n_3887), .B (n_4094), .Y (n_4503));
AND2X1 g58123(.A (n_3886), .B (n_6452), .Y (n_4378));
AND2X1 g58124(.A (n_3885), .B (n_4096), .Y (n_4376));
AND2X1 g58125(.A (n_3884), .B (n_6633), .Y (n_4374));
AND2X1 g58130(.A (n_3883), .B (n_4096), .Y (n_4372));
AND2X1 g58132(.A (n_3882), .B (n_4095), .Y (n_4370));
AND2X1 g58134(.A (n_3881), .B (n_4096), .Y (n_4368));
AND2X1 g58135(.A (n_3880), .B (n_4096), .Y (n_4366));
AND2X1 g58136(.A (n_3879), .B (n_4095), .Y (n_4364));
AND2X1 g58137(.A (n_3878), .B (n_4095), .Y (n_4362));
AND2X1 g58138(.A (n_3877), .B (n_4095), .Y (n_4360));
AND2X1 g58139(.A (n_3876), .B (n_4096), .Y (n_4358));
AND2X1 g58140(.A (n_3875), .B (n_4096), .Y (n_4356));
AND2X1 g58142(.A (n_3874), .B (n_6452), .Y (n_4354));
AND2X1 g58145(.A (n_3872), .B (n_4094), .Y (n_4350));
AND2X1 g58147(.A (n_3871), .B (n_4094), .Y (n_4348));
AND2X1 g58149(.A (n_3870), .B (n_6452), .Y (n_4346));
AND2X1 g58151(.A (n_3868), .B (n_4096), .Y (n_4342));
AND2X1 g58153(.A (n_4101), .B (n_8347), .Y (n_4340));
AND2X1 g58154(.A (n_4096), .B (n_7282), .Y (n_4338));
AND2X1 g58157(.A (n_3865), .B (n_6633), .Y (n_4336));
DFFSRX1 WX8259_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3863), .Q (), .QN (WX8259));
DFFSRX1 WX9550_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3860), .Q (), .QN (WX9550));
DFFSRX1 WX4386_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3859), .Q (), .QN (WX4386));
DFFSRX1 WX5677_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3856), .Q (), .QN (WX5677));
DFFSRX1 WX6968_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3854), .Q (), .QN (WX6968));
DFFSRX1 WX3095_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3853), .Q (), .QN (WX3095));
NOR2X1 g58604(.A (WX1838), .B (n_2620), .Y (n_4093));
NOR2X1 g58605(.A (WX10889), .B (n_1425), .Y (n_4092));
NOR2X1 g58612(.A (WX1838), .B (n_5479), .Y (n_4090));
NOR2X1 g58618(.A (WX10889), .B (n_5662), .Y (n_7510));
INVX1 g58812(.A (WX545), .Y (n_4656));
AOI21X1 g57389(.A0 (_2332_), .A1 (n_4562), .B0 (n_4087), .Y (n_4088));
NAND2X1 g57449(.A (n_9433), .B (n_4015), .Y (n_4086));
NOR2X1 g56809(.A (WX4426), .B (n_1425), .Y (n_4084));
NOR2X1 g56813(.A (WX4426), .B (n_5479), .Y (n_4083));
NAND2X1 g57874(.A (n_6645), .B (n_4078), .Y (n_4082));
NAND2X1 g57875(.A (n_4079), .B (n_4078), .Y (n_4080));
NAND2X1 g57876(.A (n_4076), .B (n_4078), .Y (n_4077));
NAND2X1 g57877(.A (n_10731), .B (n_4015), .Y (n_4075));
NAND2X1 g57878(.A (n_4071), .B (n_4078), .Y (n_4072));
NAND2X1 g57879(.A (n_4069), .B (n_4078), .Y (n_4070));
NAND2X1 g57880(.A (n_6601), .B (n_4078), .Y (n_4068));
NAND2X1 g57881(.A (n_10743), .B (n_4058), .Y (n_4066));
NAND2X1 g57882(.A (n_7074), .B (n_4078), .Y (n_4064));
NAND2X1 g57883(.A (n_4061), .B (n_4078), .Y (n_4062));
NAND2X1 g57884(.A (n_6613), .B (n_4058), .Y (n_4060));
NAND2X1 g57885(.A (n_9800), .B (n_4058), .Y (n_4057));
NAND2X1 g57886(.A (n_10727), .B (n_4015), .Y (n_4055));
NAND2X1 g57887(.A (n_4052), .B (n_4078), .Y (n_4053));
NAND2X1 g57888(.A (n_4050), .B (n_4078), .Y (n_4051));
NAND2X1 g57889(.A (n_7078), .B (n_4015), .Y (n_4049));
NAND2X1 g57890(.A (n_9437), .B (n_4015), .Y (n_4047));
NAND2X1 g57891(.A (n_4044), .B (n_3173), .Y (n_4045));
NAND2X1 g57892(.A (n_7062), .B (n_4078), .Y (n_4043));
NAND2X1 g57893(.A (n_4040), .B (n_4015), .Y (n_4041));
NAND2X1 g57894(.A (n_4038), .B (n_4078), .Y (n_4039));
NAND2X1 g57895(.A (n_7082), .B (n_4078), .Y (n_4037));
NAND2X1 g57896(.A (n_6573), .B (n_4058), .Y (n_4035));
NAND2X1 g57897(.A (n_7070), .B (n_4078), .Y (n_4033));
NAND2X1 g57898(.A (n_10747), .B (n_4015), .Y (n_4031));
NAND2X1 g57899(.A (n_10735), .B (n_4058), .Y (n_4029));
NAND2X1 g57900(.A (n_4026), .B (n_4058), .Y (n_4027));
NAND2X1 g57901(.A (n_6553), .B (n_4058), .Y (n_4025));
NAND2X1 g57902(.A (n_7066), .B (n_4078), .Y (n_4023));
NAND2X1 g57903(.A (n_10739), .B (n_4078), .Y (n_4021));
NAND2X1 g57904(.A (n_4018), .B (n_4058), .Y (n_4019));
AND2X1 g57906(.A (n_4014), .B (n_4094), .Y (n_4646));
AND2X1 g57908(.A (n_4013), .B (n_4104), .Y (n_4643));
AND2X1 g57909(.A (n_4012), .B (n_4095), .Y (n_4641));
AND2X1 g57910(.A (n_4011), .B (n_4104), .Y (n_4639));
AND2X1 g57912(.A (n_4009), .B (n_4103), .Y (n_4634));
AND2X1 g57914(.A (n_4007), .B (n_4106), .Y (n_4630));
AND2X1 g57915(.A (n_4006), .B (n_4096), .Y (n_4627));
AND2X1 g57916(.A (n_4005), .B (n_4096), .Y (n_4623));
AND2X1 g57921(.A (n_4002), .B (n_6633), .Y (n_4617));
AND2X1 g57923(.A (n_4001), .B (n_4096), .Y (n_4614));
AND2X1 g57927(.A (n_3999), .B (n_4101), .Y (n_4610));
AND2X1 g57929(.A (n_3998), .B (n_4017), .Y (n_4607));
AND2X1 g57930(.A (n_3997), .B (n_4017), .Y (n_4605));
AND2X1 g57932(.A (n_3996), .B (n_4017), .Y (n_4602));
AND2X1 g57934(.A (n_3995), .B (n_4017), .Y (n_4599));
AND2X1 g57935(.A (n_3994), .B (n_4017), .Y (n_4597));
AND2X1 g57936(.A (n_3992), .B (n_4017), .Y (n_4595));
AND2X1 g57938(.A (n_3993), .B (n_4017), .Y (n_4592));
AND2X1 g57939(.A (n_3991), .B (n_4017), .Y (n_4590));
AND2X1 g57940(.A (n_3990), .B (n_4017), .Y (n_4588));
AND2X1 g57944(.A (n_3988), .B (n_4105), .Y (n_4583));
AND2X1 g57945(.A (n_3987), .B (n_4099), .Y (n_4581));
AND2X1 g57946(.A (n_3985), .B (n_4105), .Y (n_4578));
AND2X1 g57949(.A (n_3984), .B (n_4094), .Y (n_4574));
AND2X1 g57952(.A (n_4106), .B (n_8345), .Y (n_4572));
AND2X1 g57955(.A (n_3982), .B (n_4105), .Y (n_4570));
AND2X1 g57959(.A (n_3981), .B (n_6452), .Y (n_4568));
AND2X1 g57964(.A (n_4106), .B (n_9401), .Y (n_4280));
AND2X1 g57966(.A (n_3778), .B (n_4058), .Y (n_4195));
AND2X1 g57971(.A (n_3776), .B (n_4094), .Y (n_4276));
AND2X1 g57973(.A (n_3775), .B (n_4016), .Y (n_4193));
AND2X1 g57974(.A (n_3774), .B (n_4016), .Y (n_4191));
AND2X1 g57979(.A (n_3773), .B (n_4015), .Y (n_4188));
AND2X1 g57985(.A (n_3772), .B (n_4016), .Y (n_4186));
AND2X1 g57989(.A (n_3771), .B (n_4058), .Y (n_4183));
AND2X1 g57994(.A (n_3770), .B (n_4016), .Y (n_4181));
AND2X1 g57999(.A (n_3769), .B (n_6633), .Y (n_4254));
AND2X1 g58000(.A (n_3768), .B (n_4016), .Y (n_4179));
AND2X1 g58004(.A (n_3767), .B (n_4104), .Y (n_4252));
AND2X1 g58006(.A (n_3766), .B (n_4015), .Y (n_4176));
AND2X1 g58009(.A (n_3765), .B (n_4103), .Y (n_4250));
AND2X1 g58010(.A (n_3764), .B (n_6452), .Y (n_4248));
AND2X1 g58013(.A (n_3762), .B (n_4016), .Y (n_4174));
AND2X1 g58014(.A (n_3761), .B (n_4104), .Y (n_4244));
AND2X1 g58019(.A (n_3759), .B (n_4058), .Y (n_4172));
DFFSRX1 WX8303_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3846), .Q (), .QN (WX8303));
AND2X1 g58024(.A (n_3757), .B (n_4095), .Y (n_4240));
AND2X1 g58025(.A (n_3758), .B (n_4094), .Y (n_4238));
AND2X1 g58026(.A (n_4103), .B (n_9400), .Y (n_4236));
AND2X1 g58028(.A (n_3755), .B (n_4016), .Y (n_4170));
AND2X1 g58030(.A (n_3753), .B (n_4096), .Y (n_4232));
AND2X1 g58034(.A (n_3752), .B (n_4016), .Y (n_4168));
AND2X1 g58037(.A (n_3751), .B (n_4015), .Y (n_4166));
AND2X1 g58040(.A (n_3750), .B (n_4096), .Y (n_4230));
AND2X1 g58041(.A (n_3749), .B (n_4016), .Y (n_4164));
AND2X1 g58043(.A (n_3748), .B (n_4016), .Y (n_4162));
AND2X1 g58045(.A (n_3747), .B (n_4058), .Y (n_4160));
AND2X1 g58046(.A (n_3746), .B (n_4103), .Y (n_4272));
AND2X1 g58050(.A (n_4100), .B (n_8342), .Y (n_4228));
AND2X1 g58054(.A (n_3744), .B (n_4015), .Y (n_4158));
AND2X1 g58059(.A (n_3742), .B (n_4015), .Y (n_4156));
AND2X1 g58063(.A (n_3740), .B (n_4015), .Y (n_4154));
AND2X1 g58071(.A (n_3739), .B (n_4016), .Y (n_4152));
AND2X1 g58074(.A (n_3738), .B (n_4058), .Y (n_4149));
AND2X1 g58078(.A (n_3736), .B (n_4096), .Y (n_4224));
AND2X1 g58081(.A (n_3735), .B (n_4099), .Y (n_4222));
AND2X1 g58083(.A (n_3733), .B (n_4100), .Y (n_4266));
AND2X1 g58084(.A (n_3734), .B (n_4016), .Y (n_4147));
AND2X1 g58086(.A (n_3732), .B (n_4096), .Y (n_4219));
AND2X1 g58087(.A (n_3731), .B (n_4016), .Y (n_4145));
AND2X1 g58093(.A (n_3729), .B (n_4016), .Y (n_4143));
AND2X1 g58097(.A (n_3726), .B (n_4106), .Y (n_4210));
AND2X1 g58101(.A (n_4099), .B (n_8338), .Y (n_4208));
AND2X1 g58102(.A (n_3724), .B (n_4058), .Y (n_4141));
AND2X1 g58105(.A (n_3722), .B (n_4058), .Y (n_4139));
AND2X1 g58107(.A (n_4103), .B (n_9402), .Y (n_4204));
AND2X1 g58110(.A (n_3719), .B (n_4016), .Y (n_4137));
AND2X1 g58111(.A (n_3718), .B (n_4015), .Y (n_4135));
AND2X1 g58115(.A (n_3716), .B (n_4016), .Y (n_4133));
AND2X1 g58117(.A (n_3715), .B (n_4101), .Y (n_4264));
AND2X1 g58118(.A (n_3714), .B (n_4100), .Y (n_4262));
AND2X1 g58126(.A (n_3713), .B (n_4106), .Y (n_4131));
AND2X1 g58127(.A (n_3712), .B (n_4103), .Y (n_4260));
AND2X1 g58128(.A (n_3711), .B (n_4096), .Y (n_4129));
AND2X1 g58129(.A (n_3710), .B (n_4095), .Y (n_4127));
AND2X1 g58131(.A (n_3709), .B (n_4096), .Y (n_4124));
AND2X1 g58133(.A (n_3708), .B (n_4095), .Y (n_4258));
AND2X1 g58141(.A (n_3707), .B (n_4096), .Y (n_4256));
AND2X1 g58143(.A (n_4101), .B (n_8339), .Y (n_4122));
AND2X1 g58152(.A (n_3703), .B (n_4096), .Y (n_4116));
AND2X1 g58155(.A (n_3702), .B (n_4096), .Y (n_4114));
AND2X1 g58156(.A (n_3701), .B (n_4101), .Y (n_4112));
DFFSRX1 WX9596_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3800), .Q (), .QN (WX9596));
DFFSRX1 WX545_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3696), .Q (WX545), .QN ());
NOR2X1 g57441(.A (n_3699), .B (n_3269), .Y (n_4329));
DFFSRX1 WX3131_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3694), .Q (), .QN (WX3131));
DFFSRX1 WX5717_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3691), .Q (), .QN (WX5717));
DFFSRX1 WX7010_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3848), .Q (), .QN (WX7010));
AND2X1 g57905(.A (n_3805), .B (n_4103), .Y (n_4325));
AND2X1 g57907(.A (n_3804), .B (n_4103), .Y (n_4323));
AND2X1 g57920(.A (n_3802), .B (n_4096), .Y (n_4318));
AND2X1 g57922(.A (n_3801), .B (n_4096), .Y (n_4316));
AND2X1 g57925(.A (n_3799), .B (n_4101), .Y (n_4314));
AND2X1 g57926(.A (n_3798), .B (n_4101), .Y (n_4312));
AND2X1 g57928(.A (n_3796), .B (n_4096), .Y (n_4310));
AND2X1 g57931(.A (n_3795), .B (n_4017), .Y (n_4308));
AND2X1 g57937(.A (n_3793), .B (n_4105), .Y (n_4304));
AND2X1 g57942(.A (n_3792), .B (n_4017), .Y (n_4302));
AND2X1 g57948(.A (n_3790), .B (n_4058), .Y (n_4198));
AND2X1 g57950(.A (n_4099), .B (n_8343), .Y (n_4298));
AND2X1 g57953(.A (n_3787), .B (n_4104), .Y (n_4294));
AND2X1 g57954(.A (n_3786), .B (n_4105), .Y (n_4292));
AND2X1 g57956(.A (n_3785), .B (n_4094), .Y (n_4290));
AND2X1 g57957(.A (n_4094), .B (n_8348), .Y (n_4288));
AND2X1 g57958(.A (n_3783), .B (n_4106), .Y (n_4274));
AND2X1 g57960(.A (n_3782), .B (n_4094), .Y (n_4286));
AND2X1 g57961(.A (n_3781), .B (n_4105), .Y (n_4282));
XOR2X1 g58226(.A (n_812), .B (n_3596), .Y (n_4014));
XOR2X1 g58228(.A (n_811), .B (n_3595), .Y (n_4013));
XOR2X1 g58229(.A (n_810), .B (n_3594), .Y (n_4012));
XOR2X1 g58230(.A (n_507), .B (n_3593), .Y (n_4011));
XOR2X1 g58231(.A (n_809), .B (n_3592), .Y (n_8323));
XOR2X1 g58232(.A (n_770), .B (n_3591), .Y (n_4009));
XOR2X1 g58234(.A (n_508), .B (n_3589), .Y (n_4007));
XOR2X1 g58235(.A (n_807), .B (n_3588), .Y (n_4006));
XOR2X1 g58236(.A (n_803), .B (n_3587), .Y (n_4005));
XOR2X1 g58237(.A (n_806), .B (n_3586), .Y (n_8314));
XOR2X1 g58239(.A (n_515), .B (n_3585), .Y (n_8317));
XOR2X1 g58241(.A (n_801), .B (n_3584), .Y (n_4002));
XOR2X1 g58243(.A (n_799), .B (n_3583), .Y (n_4001));
XOR2X1 g58244(.A (n_798), .B (n_3582), .Y (n_4000));
XOR2X1 g58247(.A (n_794), .B (n_3581), .Y (n_3999));
XOR2X1 g58249(.A (n_791), .B (n_3580), .Y (n_3998));
XOR2X1 g58250(.A (n_619), .B (n_3579), .Y (n_3997));
XOR2X1 g58252(.A (n_790), .B (n_3578), .Y (n_3996));
XOR2X1 g58253(.A (n_623), .B (n_3577), .Y (n_3995));
XOR2X1 g58255(.A (n_643), .B (n_3576), .Y (n_3994));
XOR2X1 g58256(.A (n_670), .B (n_3575), .Y (n_3993));
XOR2X1 g58257(.A (n_787), .B (n_3574), .Y (n_3992));
XOR2X1 g58259(.A (n_789), .B (n_3573), .Y (n_3991));
XOR2X1 g58260(.A (n_786), .B (n_3572), .Y (n_3990));
XOR2X1 g58261(.A (n_785), .B (n_3571), .Y (n_8318));
XOR2X1 g58263(.A (n_757), .B (n_3570), .Y (n_3988));
XOR2X1 g58265(.A (n_783), .B (n_3569), .Y (n_3987));
XOR2X1 g58266(.A (n_793), .B (n_3568), .Y (n_8316));
XOR2X1 g58267(.A (n_781), .B (n_3567), .Y (n_3985));
XOR2X1 g58269(.A (n_780), .B (n_3566), .Y (n_3984));
XOR2X1 g58272(.A (n_778), .B (n_3565), .Y (n_8345));
XOR2X1 g58275(.A (n_637), .B (n_3564), .Y (n_3982));
XOR2X1 g58278(.A (n_688), .B (n_3492), .Y (n_3981));
XOR2X1 g58283(.A (n_802), .B (n_3538), .Y (n_3980));
XOR2X1 g58285(.A (n_755), .B (n_3563), .Y (n_3979));
XOR2X1 g58287(.A (n_768), .B (n_3562), .Y (n_8321));
XOR2X1 g58289(.A (n_765), .B (n_3561), .Y (n_3977));
XOR2X1 g58290(.A (n_503), .B (n_3560), .Y (n_3976));
XOR2X1 g58292(.A (n_530), .B (n_3559), .Y (n_3975));
XOR2X1 g58295(.A (n_723), .B (n_3558), .Y (n_3974));
XOR2X1 g58296(.A (n_762), .B (n_3557), .Y (n_3973));
XOR2X1 g58297(.A (n_758), .B (n_3556), .Y (n_3972));
XOR2X1 g58298(.A (n_756), .B (n_3501), .Y (n_3971));
XOR2X1 g58300(.A (n_750), .B (n_3555), .Y (n_3970));
XOR2X1 g58301(.A (n_752), .B (n_3554), .Y (n_3969));
XOR2X1 g58302(.A (n_748), .B (n_3552), .Y (n_3968));
XOR2X1 g58303(.A (n_749), .B (n_3553), .Y (n_3967));
XOR2X1 g58304(.A (n_746), .B (n_3550), .Y (n_3966));
XOR2X1 g58306(.A (n_671), .B (n_3549), .Y (n_3965));
XOR2X1 g58307(.A (n_650), .B (n_3547), .Y (n_3964));
XOR2X1 g58308(.A (n_782), .B (n_3548), .Y (n_3963));
XOR2X1 g58310(.A (n_702), .B (n_3546), .Y (n_3962));
XOR2X1 g58311(.A (n_742), .B (n_3545), .Y (n_3961));
XOR2X1 g58312(.A (n_743), .B (n_3544), .Y (n_3960));
XOR2X1 g58313(.A (n_715), .B (n_3543), .Y (n_3959));
XOR2X1 g58315(.A (n_531), .B (n_3542), .Y (n_3958));
XOR2X1 g58316(.A (n_700), .B (n_3541), .Y (n_3957));
XOR2X1 g58317(.A (n_706), .B (n_3539), .Y (n_3956));
XOR2X1 g58318(.A (n_741), .B (n_3540), .Y (n_3955));
XOR2X1 g58321(.A (n_535), .B (n_3537), .Y (n_3954));
XOR2X1 g58322(.A (n_766), .B (n_3535), .Y (n_3953));
XOR2X1 g58323(.A (n_731), .B (n_3536), .Y (n_3952));
XOR2X1 g58325(.A (n_737), .B (n_3475), .Y (n_3951));
XOR2X1 g58327(.A (n_647), .B (n_3534), .Y (n_7281));
XOR2X1 g58328(.A (n_759), .B (n_3533), .Y (n_8324));
XOR2X1 g58331(.A (n_730), .B (n_3532), .Y (n_3948));
XOR2X1 g58335(.A (n_727), .B (n_3531), .Y (n_3947));
XOR2X1 g58336(.A (n_720), .B (n_3597), .Y (n_8326));
XOR2X1 g58338(.A (n_722), .B (n_3551), .Y (n_3945));
XOR2X1 g58340(.A (n_526), .B (n_3530), .Y (n_3944));
XOR2X1 g58341(.A (n_725), .B (n_3529), .Y (n_3943));
XOR2X1 g58342(.A (n_602), .B (n_6425), .Y (n_3942));
XOR2X1 g58343(.A (n_740), .B (n_3474), .Y (n_3941));
XOR2X1 g58346(.A (n_504), .B (n_3527), .Y (n_3940));
XOR2X1 g58351(.A (n_788), .B (n_3526), .Y (n_3939));
XOR2X1 g58352(.A (n_721), .B (n_3525), .Y (n_3938));
XOR2X1 g58353(.A (n_519), .B (n_3523), .Y (n_3937));
XOR2X1 g58355(.A (n_760), .B (n_3524), .Y (n_3936));
XOR2X1 g58356(.A (n_625), .B (n_3522), .Y (n_8355));
XOR2X1 g58358(.A (n_734), .B (n_3521), .Y (n_3934));
XOR2X1 g58359(.A (n_719), .B (n_3520), .Y (n_3933));
XOR2X1 g58362(.A (n_714), .B (n_3519), .Y (n_3932));
XOR2X1 g58364(.A (n_713), .B (n_3518), .Y (n_8340));
XOR2X1 g58367(.A (n_709), .B (n_3517), .Y (n_3930));
XOR2X1 g58368(.A (n_711), .B (n_3516), .Y (n_6884));
XOR2X1 g58371(.A (n_708), .B (n_3514), .Y (n_3927));
XOR2X1 g58372(.A (n_705), .B (n_3513), .Y (n_3926));
XOR2X1 g58373(.A (n_701), .B (n_3512), .Y (n_3925));
XOR2X1 g58375(.A (n_703), .B (n_3511), .Y (n_3924));
XOR2X1 g58377(.A (n_763), .B (n_3510), .Y (n_3923));
XOR2X1 g58378(.A (n_698), .B (n_3509), .Y (n_3922));
XOR2X1 g58380(.A (n_696), .B (n_3508), .Y (n_3921));
XOR2X1 g58382(.A (n_695), .B (n_3507), .Y (n_3920));
XOR2X1 g58384(.A (n_690), .B (n_3506), .Y (n_3919));
XOR2X1 g58385(.A (n_689), .B (n_3504), .Y (n_8346));
XOR2X1 g58386(.A (n_491), .B (n_3505), .Y (n_3917));
XOR2X1 g58387(.A (n_492), .B (n_3503), .Y (n_3916));
XOR2X1 g58388(.A (n_685), .B (n_3498), .Y (n_3915));
XOR2X1 g58389(.A (n_686), .B (n_3500), .Y (n_3914));
XOR2X1 g58390(.A (n_495), .B (n_3502), .Y (n_3913));
XOR2X1 g58391(.A (n_684), .B (n_3499), .Y (n_3912));
XOR2X1 g58393(.A (n_681), .B (n_3497), .Y (n_3911));
XOR2X1 g58395(.A (n_496), .B (n_3496), .Y (n_3910));
XOR2X1 g58397(.A (n_678), .B (n_3495), .Y (n_8325));
XOR2X1 g58399(.A (n_675), .B (n_3494), .Y (n_3908));
XOR2X1 g58400(.A (n_497), .B (n_3493), .Y (n_8341));
XOR2X1 g58402(.A (n_672), .B (n_3491), .Y (n_3906));
XOR2X1 g58405(.A (n_669), .B (n_3490), .Y (n_8344));
XOR2X1 g58409(.A (n_662), .B (n_3488), .Y (n_8319));
XOR2X1 g58410(.A (n_728), .B (n_3489), .Y (n_3903));
XOR2X1 g58411(.A (n_661), .B (n_3487), .Y (n_8349));
XOR2X1 g58412(.A (n_659), .B (n_3486), .Y (n_3901));
XOR2X1 g58415(.A (n_657), .B (n_3485), .Y (n_3900));
XOR2X1 g58418(.A (n_654), .B (n_3484), .Y (n_8353));
XOR2X1 g58419(.A (n_651), .B (n_3483), .Y (n_3898));
XOR2X1 g58420(.A (n_653), .B (n_3482), .Y (n_8351));
XOR2X1 g58424(.A (n_645), .B (n_3481), .Y (n_9403));
XOR2X1 g58426(.A (n_641), .B (n_3480), .Y (n_3895));
XOR2X1 g58429(.A (n_500), .B (n_3479), .Y (n_3894));
XOR2X1 g58433(.A (n_501), .B (n_3478), .Y (n_3893));
XOR2X1 g58434(.A (n_638), .B (n_3477), .Y (n_3892));
XOR2X1 g58436(.A (n_636), .B (n_3476), .Y (n_3891));
XOR2X1 g58439(.A (n_630), .B (n_7485), .Y (n_3890));
XOR2X1 g58440(.A (n_735), .B (n_3472), .Y (n_3889));
XOR2X1 g58441(.A (n_629), .B (n_3471), .Y (n_3888));
XOR2X1 g58442(.A (n_626), .B (n_3469), .Y (n_3887));
XOR2X1 g58443(.A (n_764), .B (n_3470), .Y (n_3886));
XOR2X1 g58444(.A (n_627), .B (n_3468), .Y (n_3885));
XOR2X1 g58445(.A (n_808), .B (n_3467), .Y (n_3884));
XOR2X1 g58450(.A (n_617), .B (n_3466), .Y (n_3883));
XOR2X1 g58451(.A (n_616), .B (n_3465), .Y (n_3882));
XOR2X1 g58453(.A (n_506), .B (n_3464), .Y (n_3881));
XOR2X1 g58455(.A (n_509), .B (n_3462), .Y (n_3880));
XOR2X1 g58456(.A (n_614), .B (n_3463), .Y (n_3879));
XOR2X1 g58457(.A (n_612), .B (n_3461), .Y (n_3878));
XOR2X1 g58458(.A (n_510), .B (n_3460), .Y (n_3877));
XOR2X1 g58459(.A (n_610), .B (n_3459), .Y (n_3876));
XOR2X1 g58460(.A (n_609), .B (n_3458), .Y (n_3875));
XOR2X1 g58462(.A (n_607), .B (n_3457), .Y (n_3874));
XOR2X1 g58464(.A (n_514), .B (n_3456), .Y (n_8315));
XOR2X1 g58465(.A (n_604), .B (n_3455), .Y (n_3872));
XOR2X1 g58467(.A (n_516), .B (n_3454), .Y (n_3871));
XOR2X1 g58469(.A (n_634), .B (n_3453), .Y (n_3870));
XOR2X1 g58470(.A (n_603), .B (n_3452), .Y (n_8327));
XOR2X1 g58471(.A (n_601), .B (n_3451), .Y (n_3868));
XOR2X1 g58473(.A (n_600), .B (n_3450), .Y (n_8347));
XOR2X1 g58474(.A (n_683), .B (n_3449), .Y (n_7282));
XOR2X1 g58478(.A (n_815), .B (n_3598), .Y (n_3865));
NAND2X1 g58480(.A (n_3682), .B (n_3633), .Y (n_4079));
NAND2X1 g58481(.A (n_3681), .B (n_3632), .Y (n_4076));
NAND2X2 g58483(.A (n_3678), .B (n_3628), .Y (n_4071));
NAND2X2 g58485(.A (n_3676), .B (n_3621), .Y (n_4069));
NAND2X1 g58488(.A (n_3679), .B (n_3626), .Y (n_4061));
NAND2X2 g58492(.A (n_3670), .B (n_3622), .Y (n_4052));
NAND2X1 g58493(.A (n_3669), .B (n_3620), .Y (n_4050));
NAND2X2 g58496(.A (n_3666), .B (n_3616), .Y (n_4044));
NAND2X2 g58498(.A (n_3664), .B (n_3612), .Y (n_4040));
NAND2X1 g58499(.A (n_3663), .B (n_3614), .Y (n_4038));
NAND2X1 g58505(.A (n_3658), .B (n_3609), .Y (n_4026));
NAND2X1 g58509(.A (n_3684), .B (n_3637), .Y (n_4018));
NOR2X1 g58599(.A (WX3097), .B (n_3218), .Y (n_3864));
NOR2X1 g58601(.A (WX8261), .B (n_5181), .Y (n_3863));
NOR2X1 g58603(.A (WX8261), .B (n_5838), .Y (n_6662));
NOR2X1 g58606(.A (WX9552), .B (n_2851), .Y (n_3860));
NOR2X1 g58607(.A (WX4388), .B (n_1425), .Y (n_3859));
NOR2X1 g58608(.A (WX4388), .B (n_5838), .Y (n_3857));
NOR2X1 g58610(.A (WX5679), .B (n_5712), .Y (n_3856));
NOR2X1 g58611(.A (WX5679), .B (n_5838), .Y (n_3855));
NOR2X1 g58613(.A (WX6970), .B (n_5712), .Y (n_3854));
NOR2X1 g58616(.A (WX3097), .B (n_5712), .Y (n_3853));
NOR2X1 g58617(.A (WX6970), .B (n_5662), .Y (n_6207));
NOR2X1 g58619(.A (WX9552), .B (n_5479), .Y (n_3850));
DFFSRX1 WX1838_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3647), .Q (), .QN (WX1838));
DFFSRX1 WX10889_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3650), .Q (), .QN (WX10889));
NOR2X1 g57442(.A (n_3652), .B (n_4150), .Y (n_4087));
DFFSRX1 WX4426_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3643), .Q (), .QN (WX4426));
NOR2X1 g56941(.A (WX7012), .B (n_1425), .Y (n_3848));
NOR2X1 g56978(.A (WX8305), .B (n_1425), .Y (n_3846));
NOR2X1 g56982(.A (WX8305), .B (n_5479), .Y (n_3845));
AOI22X1 g60674(.A0 (DATA_0_19), .A1 (n_3828), .B0 (_2352_), .B1(n_5873), .Y (n_3844));
AOI22X1 g60675(.A0 (DATA_0_31), .A1 (n_5968), .B0 (_2364_), .B1(n_3831), .Y (n_3843));
AOI22X1 g60676(.A0 (DATA_0_30), .A1 (n_5968), .B0 (_2363_), .B1(n_3840), .Y (n_3842));
AOI22X1 g60677(.A0 (DATA_0_29), .A1 (n_4670), .B0 (_2362_), .B1(n_3840), .Y (n_3841));
AOI22X1 g60678(.A0 (DATA_0_27), .A1 (n_3828), .B0 (_2360_), .B1(n_3840), .Y (n_3839));
AOI22X1 g60679(.A0 (DATA_0_26), .A1 (n_3828), .B0 (_2359_), .B1(n_3835), .Y (n_3837));
AOI22X1 g60680(.A0 (DATA_0_24), .A1 (n_4882), .B0 (_2357_), .B1(n_3835), .Y (n_3836));
AOI22X1 g60681(.A0 (DATA_0_28), .A1 (n_3828), .B0 (_2361_), .B1(n_3831), .Y (n_3834));
AOI22X1 g60682(.A0 (DATA_0_21), .A1 (n_5968), .B0 (_2354_), .B1(n_3831), .Y (n_3833));
AOI22X1 g60683(.A0 (DATA_0_22), .A1 (n_4670), .B0 (_2355_), .B1(n_3831), .Y (n_3830));
AOI22X1 g60684(.A0 (DATA_0_17), .A1 (n_3828), .B0 (_2350_), .B1(n_3835), .Y (n_3829));
AOI22X1 g60685(.A0 (DATA_0_23), .A1 (n_4670), .B0 (_2356_), .B1(n_3835), .Y (n_3827));
AOI22X1 g60686(.A0 (DATA_0_16), .A1 (n_4882), .B0 (_2349_), .B1(n_3835), .Y (n_3826));
AOI22X1 g60688(.A0 (DATA_0_14), .A1 (n_4882), .B0 (_2347_), .B1(n_3835), .Y (n_3824));
AOI22X1 g60690(.A0 (DATA_0_25), .A1 (n_4670), .B0 (_2358_), .B1(n_3835), .Y (n_3822));
AOI22X1 g60691(.A0 (DATA_0_12), .A1 (n_5968), .B0 (_2345_), .B1(n_3840), .Y (n_3821));
AOI22X1 g60692(.A0 (DATA_0_20), .A1 (n_5968), .B0 (_2353_), .B1(n_3840), .Y (n_3819));
AOI22X1 g60693(.A0 (DATA_0_4), .A1 (n_3828), .B0 (_2337_), .B1(n_3840), .Y (n_3818));
AOI22X1 g60694(.A0 (DATA_0_11), .A1 (n_5968), .B0 (_2344_), .B1(n_3840), .Y (n_3817));
AOI22X1 g60695(.A0 (DATA_0_10), .A1 (n_5968), .B0 (_2343_), .B1(n_3840), .Y (n_3816));
AOI22X1 g60696(.A0 (DATA_0_9), .A1 (n_5968), .B0 (_2342_), .B1(n_3840), .Y (n_3815));
AOI22X1 g60698(.A0 (DATA_0_7), .A1 (n_5968), .B0 (_2340_), .B1(n_5873), .Y (n_3813));
AOI22X1 g60699(.A0 (DATA_0_18), .A1 (n_3828), .B0 (_2351_), .B1(n_5873), .Y (n_3812));
AOI22X1 g60700(.A0 (DATA_0_6), .A1 (n_3828), .B0 (_2339_), .B1(n_3840), .Y (n_3811));
AOI22X1 g60701(.A0 (DATA_0_5), .A1 (n_3828), .B0 (_2338_), .B1(n_3840), .Y (n_3810));
AOI22X1 g60702(.A0 (DATA_0_3), .A1 (n_3828), .B0 (_2336_), .B1(n_3835), .Y (n_3809));
AOI22X1 g60703(.A0 (DATA_0_2), .A1 (n_5968), .B0 (_2335_), .B1(n_3835), .Y (n_3808));
AOI22X1 g60704(.A0 (DATA_0_1), .A1 (n_5968), .B0 (_2334_), .B1(n_3840), .Y (n_3807));
AOI22X1 g60705(.A0 (DATA_0_0), .A1 (n_3828), .B0 (_2333_), .B1(n_3835), .Y (n_3806));
XOR2X1 g58225(.A (n_538), .B (n_3409), .Y (n_3805));
XOR2X1 g58227(.A (n_814), .B (n_3408), .Y (n_3804));
XOR2X1 g58238(.A (n_805), .B (n_3403), .Y (n_9389));
XOR2X1 g58240(.A (n_804), .B (n_3402), .Y (n_3802));
XOR2X1 g58242(.A (n_800), .B (n_3401), .Y (n_3801));
NOR2X1 g57043(.A (WX9598), .B (n_5181), .Y (n_3800));
XOR2X1 g58245(.A (n_796), .B (n_3400), .Y (n_3799));
XOR2X1 g58246(.A (n_795), .B (n_3399), .Y (n_3798));
NOR2X1 g57046(.A (WX9598), .B (n_5838), .Y (n_8546));
XOR2X1 g58248(.A (n_792), .B (n_3398), .Y (n_3796));
XOR2X1 g58251(.A (n_736), .B (n_3397), .Y (n_3795));
XOR2X1 g58254(.A (n_521), .B (n_3394), .Y (n_9396));
XOR2X1 g58258(.A (n_522), .B (n_3393), .Y (n_3793));
XOR2X1 g58262(.A (n_784), .B (n_3390), .Y (n_3792));
XOR2X1 g58264(.A (n_773), .B (n_3389), .Y (n_9398));
XOR2X1 g58268(.A (n_813), .B (n_3388), .Y (n_3790));
XOR2X1 g58270(.A (n_744), .B (n_3387), .Y (n_8343));
XOR2X1 g58271(.A (n_779), .B (n_3386), .Y (n_9385));
XOR2X1 g58273(.A (n_525), .B (n_3385), .Y (n_3787));
XOR2X1 g58274(.A (n_631), .B (n_3257), .Y (n_3786));
XOR2X1 g58276(.A (n_777), .B (n_3384), .Y (n_3785));
XOR2X1 g58277(.A (n_674), .B (n_3379), .Y (n_8348));
XOR2X1 g58279(.A (n_772), .B (n_3378), .Y (n_3783));
XOR2X1 g58280(.A (n_527), .B (n_3376), .Y (n_3782));
XOR2X1 g58281(.A (n_775), .B (n_3375), .Y (n_3781));
XOR2X1 g58282(.A (n_776), .B (n_3374), .Y (n_9384));
XOR2X1 g58284(.A (n_774), .B (n_3373), .Y (n_9401));
XOR2X1 g58286(.A (n_767), .B (n_3372), .Y (n_3778));
XOR2X1 g58288(.A (n_529), .B (n_3371), .Y (n_9387));
XOR2X1 g58291(.A (n_599), .B (n_3370), .Y (n_3776));
XOR2X1 g58293(.A (n_691), .B (n_3369), .Y (n_3775));
XOR2X1 g58294(.A (n_754), .B (n_3366), .Y (n_3774));
XOR2X1 g58299(.A (n_753), .B (n_3363), .Y (n_3773));
XOR2X1 g58305(.A (n_745), .B (n_3360), .Y (n_3772));
XOR2X1 g58309(.A (n_532), .B (n_3359), .Y (n_3771));
XOR2X1 g58314(.A (n_628), .B (n_3356), .Y (n_3770));
XOR2X1 g58319(.A (n_739), .B (n_3352), .Y (n_3769));
XOR2X1 g58320(.A (n_667), .B (n_3349), .Y (n_3768));
XOR2X1 g58324(.A (n_738), .B (n_3348), .Y (n_3767));
XOR2X1 g58326(.A (n_632), .B (n_3377), .Y (n_3766));
XOR2X1 g58329(.A (n_733), .B (n_3345), .Y (n_3765));
XOR2X1 g58330(.A (n_633), .B (n_3344), .Y (n_3764));
XOR2X1 g58332(.A (n_732), .B (n_3343), .Y (n_9390));
XOR2X1 g58333(.A (n_747), .B (n_3342), .Y (n_3762));
XOR2X1 g58334(.A (n_729), .B (n_3341), .Y (n_3761));
XOR2X1 g58337(.A (n_518), .B (n_3340), .Y (n_9394));
XOR2X1 g58339(.A (n_726), .B (n_3339), .Y (n_3759));
XOR2X1 g58344(.A (n_536), .B (n_3336), .Y (n_3758));
XOR2X1 g58345(.A (n_724), .B (n_3335), .Y (n_3757));
XOR2X1 g58347(.A (n_505), .B (n_3353), .Y (n_9400));
XOR2X1 g58348(.A (n_537), .B (n_3334), .Y (n_3755));
XOR2X1 g58349(.A (n_797), .B (n_3333), .Y (n_8352));
XOR2X1 g58350(.A (n_751), .B (n_3330), .Y (n_3753));
XOR2X1 g58354(.A (n_622), .B (n_3327), .Y (n_3752));
XOR2X1 g58357(.A (n_761), .B (n_3324), .Y (n_3751));
XOR2X1 g58360(.A (n_611), .B (n_3323), .Y (n_3750));
XOR2X1 g58361(.A (n_718), .B (n_3272), .Y (n_3749));
XOR2X1 g58363(.A (n_717), .B (n_3322), .Y (n_3748));
XOR2X1 g58365(.A (n_712), .B (n_3319), .Y (n_3747));
XOR2X1 g58366(.A (n_710), .B (n_3318), .Y (n_3746));
XOR2X1 g58370(.A (n_707), .B (n_3315), .Y (n_8342));
XOR2X1 g58374(.A (n_704), .B (n_3314), .Y (n_3744));
XOR2X1 g58376(.A (n_699), .B (n_3313), .Y (n_9392));
XOR2X1 g58379(.A (n_697), .B (n_3312), .Y (n_3742));
XOR2X1 g58381(.A (n_693), .B (n_3311), .Y (n_3741));
XOR2X1 g58383(.A (n_692), .B (n_3310), .Y (n_3740));
XOR2X1 g58392(.A (n_682), .B (n_3305), .Y (n_3739));
XOR2X1 g58394(.A (n_680), .B (n_3304), .Y (n_3738));
XOR2X1 g58396(.A (n_677), .B (n_3303), .Y (n_3737));
XOR2X1 g58398(.A (n_676), .B (n_3302), .Y (n_3736));
XOR2X1 g58401(.A (n_673), .B (n_3301), .Y (n_3735));
XOR2X1 g58403(.A (n_668), .B (n_3300), .Y (n_3734));
XOR2X1 g58404(.A (n_665), .B (n_3299), .Y (n_3733));
XOR2X1 g58406(.A (n_666), .B (n_6515), .Y (n_3732));
XOR2X1 g58407(.A (n_664), .B (n_3297), .Y (n_3731));
XOR2X1 g58408(.A (n_663), .B (n_3296), .Y (n_9395));
XOR2X1 g58413(.A (n_658), .B (n_3293), .Y (n_3729));
XOR2X1 g58414(.A (n_660), .B (n_3292), .Y (n_9397));
XOR2X1 g58416(.A (n_655), .B (n_3291), .Y (n_9399));
XOR2X1 g58417(.A (n_499), .B (n_3290), .Y (n_3726));
XOR2X1 g58421(.A (n_652), .B (n_3287), .Y (n_8338));
XOR2X1 g58422(.A (n_648), .B (n_3286), .Y (n_3724));
XOR2X1 g58423(.A (n_649), .B (n_3285), .Y (n_9388));
XOR2X1 g58425(.A (n_644), .B (n_3282), .Y (n_3722));
XOR2X1 g58427(.A (n_642), .B (n_3281), .Y (n_9402));
XOR2X1 g58428(.A (n_687), .B (n_3280), .Y (n_9386));
XOR2X1 g58430(.A (n_656), .B (n_3278), .Y (n_3719));
XOR2X1 g58431(.A (n_640), .B (n_3276), .Y (n_3718));
XOR2X1 g58432(.A (n_639), .B (n_3273), .Y (n_8354));
XOR2X1 g58435(.A (n_502), .B (n_3268), .Y (n_3716));
XOR2X1 g58437(.A (n_635), .B (n_3265), .Y (n_3715));
XOR2X1 g58438(.A (n_716), .B (n_3260), .Y (n_3714));
XOR2X1 g58446(.A (n_831), .B (n_3256), .Y (n_3713));
XOR2X1 g58447(.A (n_618), .B (n_3254), .Y (n_3712));
XOR2X1 g58448(.A (n_621), .B (n_3255), .Y (n_3711));
XOR2X1 g58449(.A (n_620), .B (n_3253), .Y (n_3710));
XOR2X1 g58452(.A (n_615), .B (n_3250), .Y (n_3709));
XOR2X1 g58454(.A (n_613), .B (n_3249), .Y (n_3708));
XOR2X1 g58461(.A (n_606), .B (n_3244), .Y (n_3707));
XOR2X1 g58463(.A (n_608), .B (n_3243), .Y (n_8339));
XOR2X1 g58466(.A (n_605), .B (n_3242), .Y (n_9391));
XOR2X1 g58468(.A (n_624), .B (n_3241), .Y (n_9393));
XOR2X1 g58472(.A (n_646), .B (n_3240), .Y (n_3703));
XOR2X1 g58475(.A (n_679), .B (n_3239), .Y (n_3702));
XOR2X1 g58476(.A (n_598), .B (n_3238), .Y (n_3701));
XOR2X1 g58477(.A (n_816), .B (n_3237), .Y (n_8350));
XOR2X1 g57506(.A (n_850), .B (n_3414), .Y (n_3699));
NOR2X1 g56747(.A (WX3133), .B (n_5662), .Y (n_3698));
NOR2X1 g59506(.A (n_1425), .B (n_3695), .Y (n_3696));
NOR2X1 g56767(.A (WX3133), .B (n_1648), .Y (n_3694));
OR2X1 g59514(.A (n_3695), .B (n_5990), .Y (n_3692));
DFFSRX1 _2081__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3606), .Q (_2081_), .QN ());
DFFSRX1 _2088__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3605), .Q (_2088_), .QN ());
DFFSRX1 _2093__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3604), .Q (_2093_), .QN ());
NOR2X1 g56875(.A (WX5719), .B (n_3690), .Y (n_3691));
NOR2X1 g56880(.A (WX5719), .B (n_5427), .Y (n_3689));
NOR2X1 g56919(.A (WX7012), .B (n_5500), .Y (n_3688));
NOR2X1 g57097(.A (WX8245), .B (n_5662), .Y (n_6670));
OR2X1 g55937(.A (n_3685), .B (n_4882), .Y (n_3686));
NAND2X1 g58510(.A (n_3411), .B (n_2512), .Y (n_3684));
NAND2X1 g58514(.A (n_3405), .B (n_2454), .Y (n_3682));
NAND2X1 g58518(.A (n_3396), .B (n_2499), .Y (n_3681));
NAND2X1 g58520(.A (n_3362), .B (n_2473), .Y (n_3679));
NAND2X2 g58522(.A (n_3383), .B (n_2495), .Y (n_3678));
NAND2X2 g58526(.A (n_3365), .B (n_2447), .Y (n_3676));
NAND2X2 g58539(.A (n_3347), .B (n_2467), .Y (n_3670));
NAND2X1 g58541(.A (n_3338), .B (n_2469), .Y (n_3669));
NAND2X2 g58549(.A (n_3321), .B (n_2459), .Y (n_3666));
NAND2X2 g58552(.A (n_3309), .B (n_2438), .Y (n_3664));
NAND2X1 g58553(.A (n_3307), .B (n_2444), .Y (n_3663));
NAND2X1 g58564(.A (n_3262), .B (n_2423), .Y (n_3658));
DFFSRX1 WX8261_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3236), .Q (), .QN (WX8261));
DFFSRX1 WX9552_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3235), .Q (), .QN (WX9552));
DFFSRX1 WX4388_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3234), .Q (), .QN (WX4388));
DFFSRX1 WX5679_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3233), .Q (), .QN (WX5679));
DFFSRX1 WX6970_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3231), .Q (), .QN (WX6970));
DFFSRX1 WX3097_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3230), .Q (), .QN (WX3097));
OR2X1 g55877(.A (n_2888), .B (n_3828), .Y (n_3653));
XOR2X1 g57507(.A (n_849), .B (n_3178), .Y (n_3652));
NOR2X1 g59503(.A (WX10891), .B (n_1648), .Y (n_3650));
NOR2X1 g59510(.A (WX4390), .B (n_5479), .Y (n_6205));
NOR2X1 g59511(.A (WX1840), .B (n_5479), .Y (n_3648));
NOR2X1 g59515(.A (WX1840), .B (n_1425), .Y (n_3647));
NOR2X1 g59517(.A (WX6972), .B (n_5662), .Y (n_6677));
NOR2X1 g59518(.A (WX10891), .B (n_5662), .Y (n_7511));
NOR2X1 g56868(.A (WX4364), .B (n_2605), .Y (n_3643));
AND2X1 g56869(.A (WX4364), .B (n_5873), .Y (n_3642));
NOR2X1 g56927(.A (WX4366), .B (n_5427), .Y (n_6669));
DFFSRX1 WX7012_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3219), .Q (), .QN (WX7012));
INVX1 g60387(.A (WX547), .Y (n_3695));
NOR2X1 g56991(.A (WX5659), .B (n_5838), .Y (n_6202));
DFFSRX1 WX8305_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3217), .Q (), .QN (WX8305));
NOR2X1 g57059(.A (WX6952), .B (n_5838), .Y (n_3639));
DFFSRX1 _2152__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3210), .Q (_2152_), .QN ());
DFFSRX1 WX9598_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3216), .Q (), .QN (WX9598));
DFFSRX1 _2189__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3204), .Q (_2189_), .QN ());
NOR2X1 g57163(.A (WX9538), .B (n_5811), .Y (n_6203));
NAND2X1 g58512(.A (n_3410), .B (n_2511), .Y (n_3637));
NAND2X1 g58517(.A (n_3404), .B (n_2453), .Y (n_3633));
NAND2X1 g58521(.A (n_3395), .B (n_2498), .Y (n_3632));
NAND2X1 g58530(.A (n_3382), .B (n_2494), .Y (n_3628));
NAND2X1 g58532(.A (n_3361), .B (n_2472), .Y (n_3626));
NAND2X1 g58540(.A (n_3346), .B (n_2466), .Y (n_3622));
NAND2X1 g58543(.A (n_3364), .B (n_2446), .Y (n_3621));
NAND2X1 g58544(.A (n_3337), .B (n_2468), .Y (n_3620));
NAND2X1 g58551(.A (n_3320), .B (n_2458), .Y (n_3616));
NAND2X1 g58555(.A (n_3306), .B (n_2443), .Y (n_3614));
NAND2X1 g58561(.A (n_3308), .B (n_2437), .Y (n_3612));
NAND2X1 g58567(.A (n_3261), .B (n_2422), .Y (n_3609));
NOR2X1 g58572(.A (n_3181), .B (n_3690), .Y (n_3606));
NOR2X1 g58573(.A (n_3180), .B (n_5712), .Y (n_3605));
NOR2X1 g58574(.A (n_3179), .B (n_1648), .Y (n_3604));
AND2X1 g61727(.A (WX9556), .B (n_5873), .Y (n_6661));
AND2X1 g62334(.A (WX8265), .B (n_5873), .Y (n_3601));
OR2X1 g62530(.A (n_3599), .B (n_5990), .Y (n_3600));
XOR2X1 g58924(.A (WX4604), .B (n_3157), .Y (n_3598));
XOR2X1 g58927(.A (WX5921), .B (n_2930), .Y (n_3597));
XOR2X1 g58930(.A (WX4606), .B (n_3055), .Y (n_3596));
XOR2X1 g58931(.A (WX8525), .B (n_3155), .Y (n_3595));
XOR2X1 g58932(.A (WX4608), .B (n_3153), .Y (n_3594));
XOR2X1 g58933(.A (WX8527), .B (n_3154), .Y (n_3593));
XOR2X1 g58934(.A (WX8529), .B (n_3152), .Y (n_3592));
XOR2X1 g58935(.A (WX4610), .B (n_3151), .Y (n_3591));
XOR2X1 g58939(.A (WX4614), .B (n_3147), .Y (n_3589));
XOR2X1 g58940(.A (WX4616), .B (n_3145), .Y (n_3588));
XOR2X1 g58941(.A (WX4618), .B (n_3156), .Y (n_3587));
XOR2X1 g58944(.A (WX4620), .B (n_3142), .Y (n_3586));
XOR2X1 g58946(.A (WX4624), .B (n_3139), .Y (n_3585));
XOR2X1 g58948(.A (WX9762), .B (n_3138), .Y (n_3584));
XOR2X1 g58950(.A (WX9764), .B (n_3135), .Y (n_3583));
XOR2X1 g58951(.A (WX9766), .B (n_3134), .Y (n_3582));
XOR2X1 g58954(.A (WX9770), .B (n_3131), .Y (n_3581));
XOR2X1 g58956(.A (WX9772), .B (n_3127), .Y (n_3580));
XOR2X1 g58957(.A (WX9774), .B (n_3096), .Y (n_3579));
XOR2X1 g58959(.A (WX9776), .B (n_3125), .Y (n_3578));
XOR2X1 g58962(.A (WX9778), .B (n_2943), .Y (n_3577));
XOR2X1 g58964(.A (WX9780), .B (n_2972), .Y (n_3576));
XOR2X1 g58965(.A (WX9782), .B (n_3001), .Y (n_3575));
XOR2X1 g58967(.A (WX3295), .B (n_3123), .Y (n_3574));
XOR2X1 g58968(.A (WX9784), .B (n_3017), .Y (n_3573));
XOR2X1 g58969(.A (WX9786), .B (n_3121), .Y (n_3572));
XOR2X1 g58972(.A (WX4638), .B (n_3057), .Y (n_3571));
XOR2X1 g58974(.A (WX9790), .B (n_3118), .Y (n_3570));
XOR2X1 g58976(.A (WX9792), .B (n_3117), .Y (n_3569));
XOR2X1 g58977(.A (WX9794), .B (n_3126), .Y (n_3568));
XOR2X1 g58978(.A (WX4642), .B (n_3116), .Y (n_3567));
XOR2X1 g58980(.A (WX9796), .B (n_2954), .Y (n_3566));
XOR2X1 g58983(.A (WX9800), .B (n_2936), .Y (n_3565));
XOR2X1 g58985(.A (WX4646), .B (n_3113), .Y (n_3564));
XOR2X1 g58998(.A (WX9814), .B (n_3107), .Y (n_3563));
DFFSRX1 _2113__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3215), .Q (_2113_), .QN ());
XOR2X1 g59000(.A (WX9816), .B (n_3104), .Y (n_3562));
XOR2X1 g59002(.A (WX9820), .B (n_3101), .Y (n_3561));
XOR2X1 g59004(.A (WX3301), .B (n_3099), .Y (n_3560));
XOR2X1 g59005(.A (WX11057), .B (n_3098), .Y (n_3559));
XOR2X1 g59012(.A (WX11059), .B (n_3095), .Y (n_3558));
XOR2X1 g59013(.A (WX3303), .B (n_3093), .Y (n_3557));
XOR2X1 g59014(.A (WX3305), .B (n_3092), .Y (n_3556));
XOR2X1 g59016(.A (WX11061), .B (n_3085), .Y (n_3555));
XOR2X1 g59017(.A (WX5883), .B (n_3087), .Y (n_3554));
XOR2X1 g59018(.A (WX5885), .B (n_2957), .Y (n_3553));
XOR2X1 g59019(.A (WX3307), .B (n_2969), .Y (n_3552));
XOR2X1 g59020(.A (WX11071), .B (n_3111), .Y (n_3551));
XOR2X1 g59023(.A (WX5887), .B (n_3083), .Y (n_3550));
XOR2X1 g59025(.A (WX5889), .B (n_3081), .Y (n_3549));
XOR2X1 g59026(.A (WX5891), .B (n_3022), .Y (n_3548));
XOR2X1 g59027(.A (WX11063), .B (n_2955), .Y (n_3547));
XOR2X1 g59029(.A (WX5893), .B (n_3080), .Y (n_3546));
XOR2X1 g59030(.A (WX3309), .B (n_3043), .Y (n_3545));
XOR2X1 g59033(.A (WX5895), .B (n_3076), .Y (n_3544));
XOR2X1 g59034(.A (WX5897), .B (n_3075), .Y (n_3543));
XOR2X1 g59038(.A (WX5899), .B (n_3029), .Y (n_3542));
XOR2X1 g59039(.A (WX11065), .B (n_2958), .Y (n_3541));
XOR2X1 g59040(.A (WX5901), .B (n_3015), .Y (n_3540));
XOR2X1 g59041(.A (WX3311), .B (n_3074), .Y (n_3539));
XOR2X1 g59046(.A (WX4650), .B (n_3110), .Y (n_3538));
XOR2X1 g59048(.A (WX5905), .B (n_3071), .Y (n_3537));
XOR2X1 g59049(.A (WX5907), .B (n_3069), .Y (n_3536));
XOR2X1 g59050(.A (WX11067), .B (n_3088), .Y (n_3535));
XOR2X1 g59052(.A (WX5911), .B (n_3114), .Y (n_3534));
XOR2X1 g59053(.A (WX5913), .B (n_3128), .Y (n_3533));
XOR2X1 g59058(.A (WX11069), .B (n_3064), .Y (n_3532));
XOR2X1 g59062(.A (WX3317), .B (n_3052), .Y (n_3531));
XOR2X1 g59065(.A (WX5925), .B (n_3062), .Y (n_3530));
XOR2X1 g59066(.A (WX5927), .B (n_3090), .Y (n_3529));
XOR2X1 g59072(.A (WX11073), .B (n_3054), .Y (n_3527));
XOR2X1 g59078(.A (WX3323), .B (n_3051), .Y (n_3526));
XOR2X1 g59079(.A (WX5939), .B (n_3115), .Y (n_3525));
XOR2X1 g59082(.A (WX5941), .B (n_3066), .Y (n_3524));
XOR2X1 g59083(.A (WX11075), .B (n_3049), .Y (n_3523));
XOR2X1 g59087(.A (WX5943), .B (n_3102), .Y (n_3522));
XOR2X1 g59089(.A (WX3325), .B (n_3039), .Y (n_3521));
XOR2X1 g59090(.A (WX11077), .B (n_3065), .Y (n_3520));
XOR2X1 g59092(.A (WX11079), .B (n_3047), .Y (n_3519));
XOR2X1 g59096(.A (WX3329), .B (n_3045), .Y (n_3518));
XOR2X1 g59099(.A (WX3331), .B (n_3037), .Y (n_3517));
XOR2X1 g59100(.A (WX7174), .B (n_3038), .Y (n_3516));
XOR2X1 g59105(.A (WX7178), .B (n_3032), .Y (n_3514));
XOR2X1 g59106(.A (WX7180), .B (n_3030), .Y (n_3513));
XOR2X1 g59108(.A (WX11083), .B (n_3028), .Y (n_3512));
XOR2X1 g59109(.A (WX7182), .B (n_3026), .Y (n_3511));
XOR2X1 g59110(.A (WX7184), .B (n_3024), .Y (n_3510));
XOR2X1 g59112(.A (WX7186), .B (n_3023), .Y (n_3509));
XOR2X1 g59114(.A (WX7188), .B (n_3020), .Y (n_3508));
XOR2X1 g59116(.A (WX7190), .B (n_3018), .Y (n_3507));
XOR2X1 g59118(.A (WX7192), .B (n_3014), .Y (n_3506));
XOR2X1 g59121(.A (WX7194), .B (n_3012), .Y (n_3505));
XOR2X1 g59122(.A (WX3337), .B (n_3011), .Y (n_3504));
XOR2X1 g59125(.A (WX7196), .B (n_3009), .Y (n_3503));
XOR2X1 g59126(.A (WX3339), .B (n_3007), .Y (n_3502));
XOR2X1 g59127(.A (WX5881), .B (n_3077), .Y (n_3501));
XOR2X1 g59128(.A (WX7198), .B (n_3003), .Y (n_3500));
XOR2X1 g59129(.A (WX7200), .B (n_3000), .Y (n_3499));
XOR2X1 g59131(.A (WX11087), .B (n_3005), .Y (n_3498));
XOR2X1 g59132(.A (WX7202), .B (n_2999), .Y (n_3497));
XOR2X1 g59134(.A (WX7204), .B (n_3040), .Y (n_3496));
XOR2X1 g59135(.A (WX7206), .B (n_2997), .Y (n_3495));
XOR2X1 g59138(.A (WX7208), .B (n_2995), .Y (n_3494));
XOR2X1 g59139(.A (WX7210), .B (n_2994), .Y (n_3493));
XOR2X1 g59140(.A (WX4648), .B (n_2998), .Y (n_3492));
XOR2X1 g59142(.A (WX7212), .B (n_2992), .Y (n_3491));
XOR2X1 g59144(.A (WX7214), .B (n_2991), .Y (n_3490));
XOR2X1 g59149(.A (WX7220), .B (n_2990), .Y (n_3489));
XOR2X1 g59150(.A (WX3345), .B (n_2987), .Y (n_3488));
XOR2X1 g59151(.A (WX7222), .B (n_2985), .Y (n_3487));
XOR2X1 g59152(.A (WX11093), .B (n_2984), .Y (n_3486));
XOR2X1 g59157(.A (WX7226), .B (n_2981), .Y (n_3485));
XOR2X1 g59162(.A (WX7230), .B (n_2979), .Y (n_3484));
XOR2X1 g59163(.A (WX11095), .B (n_2975), .Y (n_3483));
XOR2X1 g59164(.A (WX3349), .B (n_2978), .Y (n_3482));
XOR2X1 g59170(.A (WX7236), .B (n_2974), .Y (n_3481));
XOR2X1 g59172(.A (WX11097), .B (n_2971), .Y (n_3480));
XOR2X1 g59176(.A (WX11099), .B (n_3048), .Y (n_3479));
XOR2X1 g59182(.A (WX11101), .B (n_2968), .Y (n_3478));
XOR2X1 g59183(.A (WX3357), .B (n_2967), .Y (n_3477));
XOR2X1 g59185(.A (WX11103), .B (n_2966), .Y (n_3476));
XOR2X1 g59186(.A (WX5909), .B (n_3141), .Y (n_3475));
XOR2X1 g59188(.A (WX5929), .B (n_3059), .Y (n_3474));
XOR2X1 g59193(.A (WX8469), .B (n_2965), .Y (n_3472));
XOR2X1 g59194(.A (WX8471), .B (n_2963), .Y (n_3471));
XOR2X1 g59197(.A (WX8473), .B (n_2961), .Y (n_3470));
XOR2X1 g59198(.A (WX11109), .B (n_3108), .Y (n_3469));
XOR2X1 g59199(.A (WX8475), .B (n_2960), .Y (n_3468));
XOR2X1 g59201(.A (WX8477), .B (n_3136), .Y (n_3467));
XOR2X1 g59206(.A (WX8485), .B (n_2952), .Y (n_3466));
XOR2X1 g59209(.A (WX8487), .B (n_2950), .Y (n_3465));
XOR2X1 g59211(.A (WX8489), .B (n_2949), .Y (n_3464));
XOR2X1 g59215(.A (WX8491), .B (n_3061), .Y (n_3463));
XOR2X1 g59216(.A (WX4590), .B (n_2948), .Y (n_3462));
XOR2X1 g59217(.A (WX8493), .B (n_2947), .Y (n_3461));
XOR2X1 g59220(.A (WX8495), .B (n_2946), .Y (n_3460));
XOR2X1 g59221(.A (WX4592), .B (n_2944), .Y (n_3459));
XOR2X1 g59222(.A (WX8497), .B (n_3068), .Y (n_3458));
XOR2X1 g59224(.A (WX4594), .B (n_2941), .Y (n_3457));
XOR2X1 g59226(.A (WX8501), .B (n_2940), .Y (n_3456));
XOR2X1 g59227(.A (WX4596), .B (n_2939), .Y (n_3455));
XOR2X1 g59229(.A (WX8505), .B (n_2937), .Y (n_3454));
XOR2X1 g59231(.A (WX4598), .B (n_2934), .Y (n_3453));
XOR2X1 g59232(.A (WX8509), .B (n_2933), .Y (n_3452));
XOR2X1 g59234(.A (WX4600), .B (n_2932), .Y (n_3451));
XOR2X1 g59235(.A (WX8513), .B (n_2982), .Y (n_3450));
XOR2X1 g59237(.A (WX4602), .B (n_2931), .Y (n_3449));
DFFSRX1 _2241__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3200), .Q (_2241_), .QN ());
NOR2X1 g59499(.A (WX3099), .B (n_5500), .Y (n_3447));
NOR2X1 g59502(.A (WX8263), .B (n_5500), .Y (n_6663));
NOR2X1 g59508(.A (WX9554), .B (n_5811), .Y (n_6204));
NOR2X1 g59509(.A (WX5681), .B (n_5811), .Y (n_6206));
DFFSRX1 WX3133_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3167), .Q (), .QN (WX3133));
DFFSRX1 WX485_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3177), .Q (WX485), .QN ());
DFFSRX1 _2317__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3190), .Q (_2317_), .QN ());
DFFSRX1 _2120__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3213), .Q (_2120_), .QN ());
DFFSRX1 _2125__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3212), .Q (_2125_), .QN ());
DFFSRX1 _2145__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3211), .Q (_2145_), .QN ());
DFFSRX1 _2157__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3208), .Q (_2157_), .QN ());
DFFSRX1 _2177__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3207), .Q (_2177_), .QN ());
DFFSRX1 _2184__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3205), .Q (_2184_), .QN ());
DFFSRX1 _2209__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3203), .Q (_2209_), .QN ());
DFFSRX1 _2216__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3202), .Q (_2216_), .QN ());
DFFSRX1 _2221__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3201), .Q (_2221_), .QN ());
DFFSRX1 _2248__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3199), .Q (_2248_), .QN ());
DFFSRX1 _2273__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3197), .Q (_2273_), .QN ());
DFFSRX1 _2285__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3194), .Q (_2285_), .QN ());
DFFSRX1 _2305__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3192), .Q (_2305_), .QN ());
DFFSRX1 _2312__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3191), .Q (_2312_), .QN ());
DFFSRX1 _2337__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3189), .Q (_2337_), .QN ());
DFFSRX1 _2344__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3187), .Q (_2344_), .QN ());
DFFSRX1 _2349__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3186), .Q (_2349_), .QN ());
DFFSRX1 _2253__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3198), .Q (_2253_), .QN ());
DFFSRX1 _2280__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3195), .Q (_2280_), .QN ());
NOR2X1 g56885(.A (WX3073), .B (n_5427), .Y (n_3443));
DFFSRX1 WX5719_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3227), .Q (), .QN (WX5719));
AND2X1 g56933(.A (WX5657), .B (n_5828), .Y (n_6212));
DFFSRX1 WX1840_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2917), .Q (), .QN (WX1840));
DFFSRX1 WX10891_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2928), .Q (), .QN (WX10891));
DFFSRX1 WX547_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2927), .Q (WX547), .QN ());
AND2X1 g57000(.A (WX6950), .B (n_5828), .Y (n_6213));
DFFSRX1 _2087__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2843), .Q (_2087_), .QN ());
AND2X1 g57038(.A (WX8243), .B (n_5828), .Y (n_6183));
DFFSRX1 _2085__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2879), .Q (_2085_), .QN ());
AND2X1 g57103(.A (WX9536), .B (n_5828), .Y (n_3439));
DFFSRX1 _2083__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2881), .Q (_2083_), .QN ());
AND2X1 g61553(.A (WX5683), .B (n_5828), .Y (n_6208));
AND2X1 g55863(.A (WX1780), .B (n_5828), .Y (n_3437));
AND2X1 g55864(.A (WX10831), .B (n_5828), .Y (n_3436));
AND2X1 g61819(.A (WX1778), .B (n_5828), .Y (n_3435));
AND2X1 g61843(.A (WX4392), .B (n_5828), .Y (n_3434));
AND2X1 g62063(.A (WX3101), .B (n_5828), .Y (n_3433));
AND2X1 g62145(.A (WX6974), .B (n_5828), .Y (n_6664));
AND2X1 g62308(.A (WX10829), .B (n_5828), .Y (n_3431));
INVX4 g62383(.A (n_3428), .Y (n_5460));
INVX4 g62393(.A (n_3428), .Y (n_5619));
INVX4 g62398(.A (n_3428), .Y (n_5556));
INVX8 g62403(.A (n_3426), .Y (n_4860));
INVX4 g62439(.A (n_3421), .Y (n_5566));
INVX8 g62441(.A (n_3421), .Y (n_4947));
INVX8 g62445(.A (n_7088), .Y (n_5722));
INVX1 g62449(.A (n_7088), .Y (n_5706));
INVX1 g62452(.A (n_7088), .Y (n_5275));
XOR2X1 g58920(.A (WX2002), .B (n_2811), .Y (n_3414));
INVX1 g58925(.A (n_3410), .Y (n_3411));
XOR2X1 g58928(.A (WX8521), .B (n_2839), .Y (n_3409));
XOR2X1 g58929(.A (WX8523), .B (n_2836), .Y (n_3408));
DFFSRX1 _2077__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2887), .Q (_2077_), .QN ());
INVX1 g58942(.A (n_3404), .Y (n_3405));
XOR2X1 g58945(.A (WX4622), .B (n_2835), .Y (n_3403));
XOR2X1 g58947(.A (WX9760), .B (n_2831), .Y (n_3402));
XOR2X1 g58949(.A (WX4626), .B (n_2830), .Y (n_3401));
XOR2X1 g58952(.A (WX4628), .B (n_2824), .Y (n_3400));
XOR2X1 g58953(.A (WX9768), .B (n_2823), .Y (n_3399));
XOR2X1 g58955(.A (WX4630), .B (n_2820), .Y (n_3398));
XOR2X1 g58958(.A (WX4632), .B (n_2818), .Y (n_3397));
INVX1 g58960(.A (n_3395), .Y (n_3396));
XOR2X1 g58963(.A (WX4634), .B (n_2816), .Y (n_3394));
XOR2X1 g58966(.A (WX4636), .B (n_2814), .Y (n_3393));
XOR2X1 g58973(.A (WX9788), .B (n_2812), .Y (n_3390));
XOR2X1 g58975(.A (WX4640), .B (n_2810), .Y (n_3389));
XOR2X1 g58979(.A (WX2004), .B (n_2807), .Y (n_3388));
XOR2X1 g58981(.A (WX9798), .B (n_2699), .Y (n_3387));
XOR2X1 g58982(.A (WX4644), .B (n_2711), .Y (n_3386));
XOR2X1 g58984(.A (WX3297), .B (n_2709), .Y (n_3385));
XOR2X1 g58986(.A (WX9804), .B (n_2806), .Y (n_3384));
INVX1 g58987(.A (n_3382), .Y (n_3383));
XOR2X1 g58991(.A (WX9806), .B (n_2805), .Y (n_3379));
XOR2X1 g58992(.A (WX11055), .B (n_2801), .Y (n_3378));
XOR2X1 g58993(.A (WX2022), .B (n_2773), .Y (n_3377));
XOR2X1 g58994(.A (WX9808), .B (n_2749), .Y (n_3376));
XOR2X1 g58995(.A (WX3299), .B (n_2794), .Y (n_3375));
XOR2X1 g58996(.A (WX9810), .B (n_2797), .Y (n_3374));
XOR2X1 g58997(.A (WX9812), .B (n_2793), .Y (n_3373));
XOR2X1 g58999(.A (WX2006), .B (n_2803), .Y (n_3372));
XOR2X1 g59001(.A (WX9818), .B (n_2792), .Y (n_3371));
XOR2X1 g59003(.A (WX9822), .B (n_2694), .Y (n_3370));
XOR2X1 g59006(.A (WX2008), .B (n_2726), .Y (n_3369));
XOR2X1 g59009(.A (WX2010), .B (n_2786), .Y (n_3366));
INVX1 g59010(.A (n_3364), .Y (n_3365));
XOR2X1 g59015(.A (WX2012), .B (n_2791), .Y (n_3363));
INVX1 g59021(.A (n_3361), .Y (n_3362));
XOR2X1 g59024(.A (WX2014), .B (n_2789), .Y (n_3360));
XOR2X1 g59028(.A (WX2016), .B (n_2787), .Y (n_3359));
XOR2X1 g59035(.A (WX2018), .B (n_2714), .Y (n_3356));
XOR2X1 g59042(.A (WX5933), .B (n_2777), .Y (n_3353));
XOR2X1 g59043(.A (WX5903), .B (n_2784), .Y (n_3352));
XOR2X1 g59047(.A (WX2020), .B (n_2700), .Y (n_3349));
XOR2X1 g59051(.A (WX3313), .B (n_2783), .Y (n_3348));
INVX1 g59054(.A (n_3346), .Y (n_3347));
XOR2X1 g59056(.A (WX3315), .B (n_2763), .Y (n_3345));
XOR2X1 g59057(.A (WX5915), .B (n_2769), .Y (n_3344));
XOR2X1 g59059(.A (WX5917), .B (n_2799), .Y (n_3343));
XOR2X1 g59060(.A (WX2024), .B (n_2703), .Y (n_3342));
XOR2X1 g59061(.A (WX5919), .B (n_2822), .Y (n_3341));
XOR2X1 g59063(.A (WX5923), .B (n_2780), .Y (n_3340));
XOR2X1 g59064(.A (WX2026), .B (n_2778), .Y (n_3339));
INVX1 g59067(.A (n_3337), .Y (n_3338));
XOR2X1 g59070(.A (WX5931), .B (n_2771), .Y (n_3336));
XOR2X1 g59071(.A (WX3321), .B (n_2695), .Y (n_3335));
XOR2X1 g59073(.A (WX2028), .B (n_2768), .Y (n_3334));
XOR2X1 g59074(.A (WX5935), .B (n_2790), .Y (n_3333));
XOR2X1 g59077(.A (WX5937), .B (n_2765), .Y (n_3330));
XOR2X1 g59084(.A (WX2030), .B (n_2774), .Y (n_3327));
XOR2X1 g59088(.A (WX2032), .B (n_2827), .Y (n_3324));
XOR2X1 g59091(.A (WX3327), .B (n_2833), .Y (n_3323));
XOR2X1 g59093(.A (WX2036), .B (n_2788), .Y (n_3322));
INVX1 g59094(.A (n_3320), .Y (n_3321));
XOR2X1 g59097(.A (WX2038), .B (n_2767), .Y (n_3319));
XOR2X1 g59098(.A (WX11081), .B (n_2762), .Y (n_3318));
XOR2X1 g59104(.A (WX3333), .B (n_2761), .Y (n_3315));
XOR2X1 g59107(.A (WX2040), .B (n_2759), .Y (n_3314));
XOR2X1 g59111(.A (WX3335), .B (n_2756), .Y (n_3313));
XOR2X1 g59113(.A (WX2042), .B (n_2754), .Y (n_3312));
XOR2X1 g59115(.A (WX11085), .B (n_2752), .Y (n_3311));
XOR2X1 g59117(.A (WX2044), .B (n_2750), .Y (n_3310));
INVX1 g59119(.A (n_3308), .Y (n_3309));
INVX1 g59123(.A (n_3306), .Y (n_3307));
XOR2X1 g59130(.A (WX2046), .B (n_2745), .Y (n_3305));
XOR2X1 g59133(.A (WX2048), .B (n_2743), .Y (n_3304));
XOR2X1 g59136(.A (WX11089), .B (n_2742), .Y (n_3303));
XOR2X1 g59137(.A (WX3341), .B (n_2741), .Y (n_3302));
XOR2X1 g59141(.A (WX3343), .B (n_2738), .Y (n_3301));
XOR2X1 g59143(.A (WX2050), .B (n_2737), .Y (n_3300));
XOR2X1 g59145(.A (WX11091), .B (n_2736), .Y (n_3299));
XOR2X1 g59147(.A (WX2052), .B (n_2733), .Y (n_3297));
XOR2X1 g59148(.A (WX7218), .B (n_2732), .Y (n_3296));
XOR2X1 g59155(.A (WX2054), .B (n_2731), .Y (n_3293));
XOR2X1 g59156(.A (WX7224), .B (n_2730), .Y (n_3292));
XOR2X1 g59158(.A (WX3347), .B (n_2729), .Y (n_3291));
XOR2X1 g59159(.A (WX7228), .B (n_2728), .Y (n_3290));
XOR2X1 g59165(.A (WX7232), .B (n_2725), .Y (n_3287));
XOR2X1 g59166(.A (WX2056), .B (n_2724), .Y (n_3286));
XOR2X1 g59167(.A (WX7234), .B (n_2722), .Y (n_3285));
XOR2X1 g59171(.A (WX2058), .B (n_2721), .Y (n_3282));
XOR2X1 g59173(.A (WX3351), .B (n_2720), .Y (n_3281));
XOR2X1 g59174(.A (WX3353), .B (n_2719), .Y (n_3280));
INVX2 g63085(.A (n_5873), .Y (n_5822));
XOR2X1 g59175(.A (WX2060), .B (n_2718), .Y (n_3278));
INVX2 g63101(.A (n_4150), .Y (n_5052));
INVX4 g63107(.A (n_3221), .Y (n_5968));
XOR2X1 g59177(.A (WX2062), .B (n_2772), .Y (n_3276));
XOR2X1 g59180(.A (WX3355), .B (n_2717), .Y (n_3273));
XOR2X1 g59181(.A (WX2034), .B (n_2782), .Y (n_3272));
INVX8 g63165(.A (n_6440), .Y (n_4882));
INVX4 g63172(.A (n_3269), .Y (n_3828));
XOR2X1 g59184(.A (WX2064), .B (n_2715), .Y (n_3268));
INVX8 g63194(.A (n_3264), .Y (n_5662));
XOR2X1 g59187(.A (WX11105), .B (n_2713), .Y (n_3265));
INVX8 g63212(.A (n_3263), .Y (n_5479));
INVX1 g59189(.A (n_3261), .Y (n_3262));
XOR2X1 g59191(.A (WX11107), .B (n_2710), .Y (n_3260));
XOR2X1 g59200(.A (WX9802), .B (n_2708), .Y (n_3257));
XOR2X1 g59202(.A (WX8479), .B (n_2707), .Y (n_3256));
XOR2X1 g59203(.A (WX8481), .B (n_2706), .Y (n_3255));
XOR2X1 g59204(.A (WX11111), .B (n_2705), .Y (n_3254));
XOR2X1 g59205(.A (WX8483), .B (n_2704), .Y (n_3253));
XOR2X1 g59210(.A (WX4588), .B (n_2702), .Y (n_3250));
XOR2X1 g59212(.A (WX11113), .B (n_2701), .Y (n_3249));
XOR2X1 g59223(.A (WX11115), .B (n_2698), .Y (n_3244));
XOR2X1 g59225(.A (WX8499), .B (n_2697), .Y (n_3243));
XOR2X1 g59228(.A (WX8503), .B (n_2696), .Y (n_3242));
XOR2X1 g59230(.A (WX8507), .B (n_2712), .Y (n_3241));
XOR2X1 g59233(.A (WX8511), .B (n_2734), .Y (n_3240));
XOR2X1 g59236(.A (WX8515), .B (n_2739), .Y (n_3239));
XOR2X1 g59238(.A (WX8517), .B (n_2746), .Y (n_3238));
XOR2X1 g59239(.A (WX8519), .B (n_2760), .Y (n_3237));
NOR2X1 g59501(.A (WX8263), .B (n_5712), .Y (n_3236));
NOR2X1 g59504(.A (WX9554), .B (n_1648), .Y (n_3235));
NOR2X1 g59505(.A (WX4390), .B (n_3188), .Y (n_3234));
NOR2X1 g59507(.A (WX5681), .B (n_5712), .Y (n_3233));
NOR2X1 g59513(.A (WX6972), .B (n_5712), .Y (n_3231));
NOR2X1 g59516(.A (WX3099), .B (n_3188), .Y (n_3230));
DFFSRX1 _2094__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2872), .Q (_2094_), .QN ());
DFFSRX1 _2099__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2868), .Q (_2099_), .QN ());
DFFSRX1 _2103__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2846), .Q (_2103_), .QN ());
DFFSRX1 _2108__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2898), .Q (_2108_), .QN ());
DFFSRX1 _2118__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2861), .Q (_2118_), .QN ());
DFFSRX1 _2080__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2883), .Q (_2080_), .QN ());
DFFSRX1 _2078__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2885), .Q (_2078_), .QN ());
DFFSRX1 _2079__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2884), .Q (_2079_), .QN ());
DFFSRX1 _2082__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2882), .Q (_2082_), .QN ());
DFFSRX1 _2084__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2850), .Q (_2084_), .QN ());
DFFSRX1 _2086__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2878), .Q (_2086_), .QN ());
DFFSRX1 _2090__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2875), .Q (_2090_), .QN ());
DFFSRX1 _2091__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2852), .Q (_2091_), .QN ());
DFFSRX1 _2092__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2873), .Q (_2092_), .QN ());
DFFSRX1 _2095__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2870), .Q (_2095_), .QN ());
DFFSRX1 _2096__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2844), .Q (_2096_), .QN ());
DFFSRX1 _2098__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2893), .Q (_2098_), .QN ());
DFFSRX1 _2100__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2856), .Q (_2100_), .QN ());
DFFSRX1 _2101__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2867), .Q (_2101_), .QN ());
DFFSRX1 _2102__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2854), .Q (_2102_), .QN ());
DFFSRX1 _2104__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2866), .Q (_2104_), .QN ());
DFFSRX1 _2105__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2865), .Q (_2105_), .QN ());
DFFSRX1 _2106__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2864), .Q (_2106_), .QN ());
DFFSRX1 _2131__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2889), .Q (_2131_), .QN ());
AND2X1 g56826(.A (WX3071), .B (n_5828), .Y (n_6182));
DFFSRX1 _2183__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2860), .Q (_2183_), .QN ());
DFFSRX1 _2185__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2859), .Q (_2185_), .QN ());
DFFSRX1 _2198__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2892), .Q (_2198_), .QN ());
DFFSRX1 _2271__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2858), .Q (_2271_), .QN ());
DFFSRX1 _2272__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2857), .Q (_2272_), .QN ());
DFFSRX1 _2331__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2847), .Q (_2331_), .QN ());
DFFSRX1 _2362__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2848), .Q (_2362_), .QN ());
DFFSRX1 _2097__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2855), .Q (_2097_), .QN ());
DFFSRX1 _2089__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2876), .Q (_2089_), .QN ());
DFFSRX1 _2107__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2863), .Q (_2107_), .QN ());
DFFSRX1 WX721_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2907), .Q (WX721), .QN ());
DFFSRX1 WX725_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2914), .Q (WX725), .QN ());
DFFSRX1 WX727_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2916), .Q (WX727), .QN ());
DFFSRX1 WX745_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2903), .Q (WX745), .QN ());
DFFSRX1 WX831_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2911), .Q (WX831), .QN ());
DFFSRX1 WX835_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2909), .Q (WX835), .QN ());
DFFSRX1 WX899_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2912), .Q (WX899), .QN ());
DFFSRX1 WX845_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2908), .Q (WX845), .QN ());
DFFSRX1 WX873_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2902), .Q (WX873), .QN ());
DFFSRX1 WX895_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2906), .Q (WX895), .QN ());
DFFSRX1 WX2032_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2900), .Q (WX2032), .QN ());
DFFSRX1 WX715_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2905), .Q (WX715), .QN ());
DFFSRX1 WX4364_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_3163), .Q (WX4364), .QN ());
NOR2X1 g56932(.A (WX5657), .B (n_2605), .Y (n_3227));
DFFSRX1 _2334__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2583), .Q (_2334_), .QN ());
BUFX3 g63099(.A (n_3221), .Y (n_3840));
BUFX3 g63100(.A (n_3221), .Y (n_3835));
CLKBUFX3 g63103(.A (n_3221), .Y (n_4150));
BUFX3 g63094(.A (n_3221), .Y (n_4600));
BUFX3 g63092(.A (n_3221), .Y (n_4579));
BUFX3 g63093(.A (n_3221), .Y (n_4439));
BUFX3 g63090(.A (n_3221), .Y (n_4608));
NOR2X1 g56999(.A (WX6950), .B (n_2605), .Y (n_3219));
INVX4 g63058(.A (n_3831), .Y (n_3218));
NOR2X1 g57037(.A (WX8243), .B (n_2849), .Y (n_3217));
NOR2X1 g57102(.A (WX9536), .B (n_2605), .Y (n_3216));
DFFSRX1 _2308__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2567), .Q (_2308_), .QN ());
NOR2X1 g58575(.A (n_2658), .B (n_5712), .Y (n_3215));
NOR2X1 g58576(.A (n_2662), .B (n_5712), .Y (n_3213));
NOR2X1 g58577(.A (n_2656), .B (n_5712), .Y (n_3212));
NOR2X1 g58578(.A (n_2655), .B (n_5181), .Y (n_3211));
NOR2X1 g58579(.A (n_2654), .B (n_1425), .Y (n_3210));
NOR2X1 g58580(.A (n_2653), .B (n_3690), .Y (n_3208));
NOR2X1 g58581(.A (n_2652), .B (n_3690), .Y (n_3207));
NOR2X1 g58582(.A (n_2661), .B (n_2851), .Y (n_3205));
NOR2X1 g58583(.A (n_2651), .B (n_2849), .Y (n_3204));
NOR2X1 g58584(.A (n_2649), .B (n_1425), .Y (n_3203));
NOR2X1 g58585(.A (n_2647), .B (n_5181), .Y (n_3202));
NOR2X1 g58586(.A (n_2646), .B (n_5712), .Y (n_3201));
NOR2X1 g58587(.A (n_2644), .B (n_5712), .Y (n_3200));
NOR2X1 g58588(.A (n_2648), .B (n_1648), .Y (n_3199));
NOR2X1 g58589(.A (n_2643), .B (n_1425), .Y (n_3198));
NOR2X1 g58590(.A (n_2642), .B (n_1648), .Y (n_3197));
NOR2X1 g58591(.A (n_2641), .B (n_1425), .Y (n_3195));
NOR2X1 g58592(.A (n_2657), .B (n_5712), .Y (n_3194));
NOR2X1 g58593(.A (n_2635), .B (n_5712), .Y (n_3192));
NOR2X1 g58594(.A (n_2640), .B (n_3188), .Y (n_3191));
NOR2X1 g58595(.A (n_2634), .B (n_1425), .Y (n_3190));
NOR2X1 g58596(.A (n_2639), .B (n_3188), .Y (n_3189));
NOR2X1 g58597(.A (n_2637), .B (n_1425), .Y (n_3187));
NOR2X1 g58598(.A (n_2636), .B (n_3188), .Y (n_3186));
INVX4 g62395(.A (n_6614), .Y (n_3428));
INVX4 g62406(.A (n_6497), .Y (n_3426));
INVX8 g62432(.A (n_3183), .Y (n_3421));
XOR2X1 g58893(.A (_2080_), .B (n_2544), .Y (n_3181));
XOR2X1 g58898(.A (_2087_), .B (n_2540), .Y (n_3180));
XOR2X1 g58899(.A (_2092_), .B (n_2537), .Y (n_3179));
XOR2X1 g58921(.A (WX11053), .B (n_2496), .Y (n_3178));
MX2X1 g58926(.A (n_18), .B (WX753), .S0 (n_2514), .Y (n_3410));
MX2X1 g58943(.A (n_19), .B (WX755), .S0 (n_2406), .Y (n_3404));
AND2X1 g55873(.A (n_2378), .B (WX487), .Y (n_3177));
MX2X1 g58961(.A (n_67), .B (WX757), .S0 (n_2500), .Y (n_3395));
MX2X1 g58988(.A (n_12), .B (WX721), .S0 (n_2487), .Y (n_3382));
MX2X1 g59011(.A (n_71), .B (WX715), .S0 (n_2471), .Y (n_3364));
MX2X1 g59022(.A (n_112), .B (WX763), .S0 (n_2477), .Y (n_3361));
MX2X1 g59055(.A (n_85), .B (WX767), .S0 (n_2470), .Y (n_3346));
MX2X1 g59068(.A (n_87), .B (WX769), .S0 (n_2480), .Y (n_3337));
MX2X1 g59095(.A (n_20), .B (WX741), .S0 (n_2462), .Y (n_3320));
MX2X1 g59120(.A (n_2), .B (WX717), .S0 (n_2445), .Y (n_3308));
MX2X1 g59124(.A (n_16), .B (WX743), .S0 (n_2448), .Y (n_3306));
INVX8 g63064(.A (n_3173), .Y (n_5889));
INVX2 g63083(.A (n_6626), .Y (n_5873));
BUFX3 g63091(.A (n_3221), .Y (n_4468));
BUFX3 g63095(.A (n_3221), .Y (n_4603));
BUFX3 g63096(.A (n_3221), .Y (n_4586));
BUFX3 g63097(.A (n_3221), .Y (n_4615));
INVX8 g63116(.A (n_3222), .Y (n_5427));
INVX8 g63127(.A (n_3223), .Y (n_5811));
INVX8 g63135(.A (n_3224), .Y (n_5500));
INVX8 g63145(.A (n_3225), .Y (n_5838));
INVX4 g63189(.A (n_3169), .Y (n_4015));
INVX4 g63213(.A (n_3168), .Y (n_3263));
MX2X1 g59190(.A (n_106), .B (WX749), .S0 (n_2424), .Y (n_3261));
DFFSRX1 _2332__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2585), .Q (_2332_), .QN ());
DFFSRX1 _2363__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2572), .Q (_2363_), .QN ());
DFFSRX1 _2328__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2587), .Q (_2328_), .QN ());
DFFSRX1 _2140__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2631), .Q (_2140_), .QN ());
DFFSRX1 WX11181_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2678), .Q (), .QN (WX11181));
DFFSRX1 _2150__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2571), .Q (_2150_), .QN ());
DFFSRX1 _2293__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2596), .Q (_2293_), .QN ());
DFFSRX1 _2119__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2621), .Q (_2119_), .QN ());
DFFSRX1 _2121__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2619), .Q (_2121_), .QN ());
DFFSRX1 _2139__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2629), .Q (_2139_), .QN ());
DFFSRX1 _2162__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2618), .Q (_2162_), .QN ());
DFFSRX1 _2163__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2617), .Q (_2163_), .QN ());
DFFSRX1 _2171__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2622), .Q (_2171_), .QN ());
DFFSRX1 _2174__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2616), .Q (_2174_), .QN ());
DFFSRX1 _2175__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2615), .Q (_2175_), .QN ());
DFFSRX1 _2181__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2563), .Q (_2181_), .QN ());
DFFSRX1 _2194__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2613), .Q (_2194_), .QN ());
DFFSRX1 _2201__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2612), .Q (_2201_), .QN ());
DFFSRX1 _2202__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2611), .Q (_2202_), .QN ());
DFFSRX1 _2205__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2610), .Q (_2205_), .QN ());
DFFSRX1 _2207__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2609), .Q (_2207_), .QN ());
DFFSRX1 _2218__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2608), .Q (_2218_), .QN ());
DFFSRX1 _2220__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2565), .Q (_2220_), .QN ());
DFFSRX1 _2224__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2607), .Q (_2224_), .QN ());
DFFSRX1 _2232__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2600), .Q (_2232_), .QN ());
DFFSRX1 _2237__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2606), .Q (_2237_), .QN ());
DFFSRX1 _2240__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2604), .Q (_2240_), .QN ());
DFFSRX1 _2244__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2564), .Q (_2244_), .QN ());
DFFSRX1 _2246__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2566), .Q (_2246_), .QN ());
DFFSRX1 _2250__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2625), .Q (_2250_), .QN ());
DFFSRX1 _2258__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2602), .Q (_2258_), .QN ());
DFFSRX1 _2262__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2601), .Q (_2262_), .QN ());
DFFSRX1 _2263__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2626), .Q (_2263_), .QN ());
DFFSRX1 _2268__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2599), .Q (_2268_), .QN ());
DFFSRX1 _2281__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2570), .Q (_2281_), .QN ());
DFFSRX1 _2289__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2598), .Q (_2289_), .QN ());
DFFSRX1 _2292__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2597), .Q (_2292_), .QN ());
DFFSRX1 _2295__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2624), .Q (_2295_), .QN ());
DFFSRX1 _2298__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2628), .Q (_2298_), .QN ());
DFFSRX1 _2301__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2595), .Q (_2301_), .QN ());
DFFSRX1 _2302__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2594), .Q (_2302_), .QN ());
DFFSRX1 _2303__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2593), .Q (_2303_), .QN ());
DFFSRX1 _2306__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2591), .Q (_2306_), .QN ());
DFFSRX1 _2307__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2590), .Q (_2307_), .QN ());
DFFSRX1 _2309__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2627), .Q (_2309_), .QN ());
DFFSRX1 _2319__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2589), .Q (_2319_), .QN ());
DFFSRX1 _2327__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2588), .Q (_2327_), .QN ());
DFFSRX1 _2333__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2584), .Q (_2333_), .QN ());
DFFSRX1 _2335__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2582), .Q (_2335_), .QN ());
DFFSRX1 _2348__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2581), .Q (_2348_), .QN ());
DFFSRX1 _2350__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2579), .Q (_2350_), .QN ());
DFFSRX1 _2352__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2576), .Q (_2352_), .QN ());
DFFSRX1 _2353__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2575), .Q (_2353_), .QN ());
DFFSRX1 _2354__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2574), .Q (_2354_), .QN ());
DFFSRX1 _2264__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2568), .Q (_2264_), .QN ());
DFFSRX1 WX11115_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2663), .Q (WX11115), .QN ());
DFFSRX1 WX11153_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2689), .Q (WX11153), .QN ());
DFFSRX1 WX7216_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2677), .Q (WX7216), .QN ());
DFFSRX1 WX7272_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2630), .Q (WX7272), .QN ());
DFFSRX1 WX4606_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2682), .Q (WX4606), .QN ());
DFFSRX1 WX11199_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2686), .Q (WX11199), .QN ());
DFFSRX1 WX11235_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2650), .Q (WX11235), .QN ());
DFFSRX1 WX11239_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2690), .Q (WX11239), .QN ());
DFFSRX1 WX4674_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2665), .Q (WX4674), .QN ());
DFFSRX1 WX3369_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2666), .Q (WX3369), .QN ());
DFFSRX1 WX3401_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2645), .Q (WX3401), .QN ());
DFFSRX1 WX3433_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2667), .Q (WX3433), .QN ());
DFFSRX1 WX3439_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2668), .Q (WX3439), .QN ());
DFFSRX1 WX11169_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2680), .Q (WX11169), .QN ());
DFFSRX1 WX8649_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2660), .Q (WX8649), .QN ());
DFFSRX1 WX8651_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2659), .Q (WX8651), .QN ());
DFFSRX1 WX9804_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2562), .Q (WX9804), .QN ());
DFFSRX1 WX9828_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2671), .Q (WX9828), .QN ());
DFFSRX1 WX9834_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2687), .Q (WX9834), .QN ());
DFFSRX1 WX9872_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2681), .Q (WX9872), .QN ());
DFFSRX1 WX9926_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2673), .Q (WX9926), .QN ());
DFFSRX1 WX4620_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2685), .Q (WX4620), .QN ());
DFFSRX1 WX4638_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2614), .Q (WX4638), .QN ());
DFFSRX1 WX4746_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2670), .Q (WX4746), .QN ());
DFFSRX1 WX4754_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2669), .Q (WX4754), .QN ());
DFFSRX1 WX5927_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2638), .Q (WX5927), .QN ());
DFFSRX1 WX6051_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2664), .Q (WX6051), .QN ());
DFFSRX1 WX2050_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2692), .Q (WX2050), .QN ());
DFFSRX1 WX2064_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2676), .Q (WX2064), .QN ());
DFFSRX1 WX2098_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2633), .Q (WX2098), .QN ());
DFFSRX1 WX2146_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2632), .Q (WX2146), .QN ());
DFFSRX1 WX11207_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2684), .Q (WX11207), .QN ());
INVX4 g63208(.A (n_3168), .Y (n_3264));
DFFSRX1 _2242__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2603), .Q (_2242_), .QN ());
NOR2X1 g56825(.A (WX3071), .B (n_2849), .Y (n_3167));
DFFSRX1 _2355__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2573), .Q (_2355_), .QN ());
DFFSRX1 _2351__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2577), .Q (_2351_), .QN ());
INVX2 g63177(.A (n_4184), .Y (n_5990));
INVX2 g63174(.A (n_4670), .Y (n_3269));
INVX2 g63162(.A (n_6438), .Y (n_6440));
DFFSRX1 WX9816_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1678), .Q (WX9816), .QN ());
NOR2X1 g56925(.A (WX4366), .B (n_2849), .Y (n_3163));
DFFSRX1 WX9924_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2307), .Q (WX9924), .QN ());
DFFSRX1 WX8263_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1487), .Q (), .QN (WX8263));
DFFSRX1 WX7206_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1956), .Q (WX7206), .QN ());
DFFSRX1 WX11237_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1830), .Q (WX11237), .QN ());
DFFSRX1 WX6972_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1720), .Q (), .QN (WX6972));
BUFX3 g63138(.A (n_3162), .Y (n_3224));
DFFSRX1 WX7202_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2196), .Q (WX7202), .QN ());
DFFSRX1 WX1778_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2405), .Q (WX1778), .QN ());
DFFSRX1 _2346__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1524), .Q (_2346_), .QN ());
DFFSRX1 WX4758_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1928), .Q (WX4758), .QN ());
DFFSRX1 _2270__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1565), .Q (_2270_), .QN ());
DFFSRX1 _2296__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1688), .Q (_2296_), .QN ());
DFFSRX1 _2347__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1694), .Q (_2347_), .QN ());
BUFX3 g63129(.A (n_3162), .Y (n_3223));
DFFSRX1 _2196__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1605), .Q (_2196_), .QN ());
DFFSRX1 WX6025_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1905), .Q (WX6025), .QN ());
DFFSRX1 WX3099_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1900), .Q (), .QN (WX3099));
DFFSRX1 _2235__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1582), .Q (_2235_), .QN ());
DFFSRX1 WX8631_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2094), .Q (WX8631), .QN ());
BUFX3 g63120(.A (n_3162), .Y (n_3222));
INVX4 g63109(.A (n_6626), .Y (n_3221));
DFFSRX1 WX2166_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2055), .Q (WX2166), .QN ());
DFFSRX1 _2161__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1633), .Q (_2161_), .QN ());
DFFSRX1 _2127__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1658), .Q (_2127_), .QN ());
DFFSRX1 WX11079_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2085), .Q (WX11079), .QN ());
DFFSRX1 WX5893_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2525), .Q (WX5893), .QN ());
DFFSRX1 WX8543_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1891), .Q (WX8543), .QN ());
DFFSRX1 _2182__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1615), .Q (_2182_), .QN ());
DFFSRX1 _2158__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1636), .Q (_2158_), .QN ());
DFFSRX1 WX2174_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1922), .Q (WX2174), .QN ());
DFFSRX1 WX2156_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2002), .Q (WX2156), .QN ());
DFFSRX1 _2124__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1660), .Q (_2124_), .QN ());
DFFSRX1 _2160__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1503), .Q (_2160_), .QN ());
BUFX3 g63074(.A (n_4562), .Y (n_4628));
BUFX3 g63088(.A (n_6626), .Y (n_4105));
DFFSRX1 WX11063_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2013), .Q (WX11063), .QN ());
DFFSRX1 _2197__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1604), .Q (_2197_), .QN ());
DFFSRX1 WX2192_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2247), .Q (WX2192), .QN ());
DFFSRX1 WX2182_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2194), .Q (WX2182), .QN ());
BUFX3 g63076(.A (n_4562), .Y (n_4471));
DFFSRX1 _2236__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1581), .Q (_2236_), .QN ());
DFFSRX1 WX11129_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1951), .Q (WX11129), .QN ());
INVX2 g63065(.A (n_3158), .Y (n_3173));
DFFSRX1 WX4734_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2067), .Q (WX4734), .QN ());
DFFSRX1 WX11071_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1737), .Q (WX11071), .QN ());
DFFSRX1 WX2124_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2172), .Q (WX2124), .QN ());
DFFSRX1 _2212__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1597), .Q (_2212_), .QN ());
DFFSRX1 WX4690_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2193), .Q (WX4690), .QN ());
DFFSRX1 WX4596_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1723), .Q (WX4596), .QN ());
DFFSRX1 WX4716_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2143), .Q (WX4716), .QN ());
CLKBUFX3 g63060(.A (n_3158), .Y (n_3831));
MX2X1 g60707(.A (n_3027), .B (n_6422), .S0 (WX4540), .Y (n_3157));
MX2X1 g60711(.A (n_3140), .B (n_2938), .S0 (WX4554), .Y (n_3156));
DFFSRX1 WX4612_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2035), .Q (WX4612), .QN ());
MX2X1 g60716(.A (n_3058), .B (n_2775), .S0 (WX8461), .Y (n_3155));
MX2X1 g60718(.A (n_3106), .B (n_2837), .S0 (WX8463), .Y (n_3154));
MX2X1 g60719(.A (n_3137), .B (n_3086), .S0 (WX4544), .Y (n_3153));
MX2X1 g60722(.A (n_2776), .B (n_2996), .S0 (WX8465), .Y (n_3152));
MX2X1 g60726(.A (n_3137), .B (n_2938), .S0 (WX4546), .Y (n_3151));
DFFSRX1 _2278__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1500), .Q (_2278_), .QN ());
MX2X1 g60729(.A (n_3137), .B (n_3072), .S0 (WX4548), .Y (n_3149));
MX2X1 g60733(.A (n_3021), .B (n_3086), .S0 (WX4550), .Y (n_3147));
MX2X1 g60735(.A (n_3021), .B (n_3041), .S0 (WX4552), .Y (n_3145));
MX2X1 g60739(.A (n_2798), .B (n_3004), .S0 (WX4556), .Y (n_3142));
DFFSRX1 WX4652_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2159), .Q (WX4652), .QN ());
MX2X1 g60745(.A (n_3140), .B (n_3086), .S0 (WX5845), .Y (n_3141));
MX2X1 g60746(.A (n_2986), .B (n_3056), .S0 (WX4560), .Y (n_3139));
MX2X1 g60751(.A (n_3137), .B (n_3086), .S0 (WX9698), .Y (n_3138));
DFFSRX1 WX4654_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1870), .Q (WX4654), .QN ());
MX2X1 g60755(.A (n_3137), .B (n_7488), .S0 (WX8413), .Y (n_3136));
MX2X1 g60758(.A (n_3031), .B (n_2938), .S0 (WX9700), .Y (n_3135));
MX2X1 g60761(.A (n_3031), .B (n_3041), .S0 (WX9702), .Y (n_3134));
MX2X1 g60769(.A (n_3027), .B (n_6422), .S0 (WX9706), .Y (n_3131));
MX2X1 g60774(.A (n_2815), .B (n_2976), .S0 (WX5849), .Y (n_3128));
MX2X1 g60776(.A (n_3137), .B (n_2945), .S0 (WX9708), .Y (n_3127));
MX2X1 g60780(.A (n_2838), .B (n_3044), .S0 (WX9730), .Y (n_3126));
DFFSRX1 WX7244_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1672), .Q (WX7244), .QN ());
DFFSRX1 WX9786_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2138), .Q (WX9786), .QN ());
MX2X1 g60782(.A (n_3137), .B (n_6422), .S0 (WX9712), .Y (n_3125));
MX2X1 g60788(.A (n_3120), .B (n_7488), .S0 (WX3231), .Y (n_3123));
MX2X1 g60793(.A (n_3120), .B (n_3086), .S0 (WX9722), .Y (n_3121));
MX2X1 g60801(.A (n_3140), .B (n_3072), .S0 (WX9726), .Y (n_3118));
DFFSRX1 _2287__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1557), .Q (_2287_), .QN ());
MX2X1 g60805(.A (n_3058), .B (n_3105), .S0 (WX9728), .Y (n_3117));
MX2X1 g60810(.A (n_3106), .B (n_3103), .S0 (WX4578), .Y (n_3116));
DFFSRX1 WX7290_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2305), .Q (WX7290), .QN ());
MX2X1 g60811(.A (n_3106), .B (n_2775), .S0 (WX5875), .Y (n_3115));
MX2X1 g60816(.A (n_3031), .B (n_2945), .S0 (WX5847), .Y (n_3114));
MX2X1 g60821(.A (n_3058), .B (n_2837), .S0 (WX4582), .Y (n_3113));
DFFSRX1 WX7294_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2320), .Q (WX7294), .QN ());
MX2X1 g60828(.A (n_3031), .B (n_3041), .S0 (WX11007), .Y (n_3111));
DFFSRX1 WX7330_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1709), .Q (WX7330), .QN ());
DFFSRX1 WX4702_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2233), .Q (WX4702), .QN ());
MX2X1 g60838(.A (n_3106), .B (n_2837), .S0 (WX4586), .Y (n_3110));
MX2X1 g60843(.A (n_3106), .B (n_3089), .S0 (WX11045), .Y (n_3108));
MX2X1 g60846(.A (n_3106), .B (n_3105), .S0 (WX9750), .Y (n_3107));
MX2X1 g60848(.A (n_2935), .B (n_3103), .S0 (WX9752), .Y (n_3104));
MX2X1 g60856(.A (n_2798), .B (n_3105), .S0 (WX5879), .Y (n_3102));
MX2X1 g60857(.A (n_3106), .B (n_3089), .S0 (WX9756), .Y (n_3101));
DFFSRX1 WX7196_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2181), .Q (WX7196), .QN ());
MX2X1 g60860(.A (n_3027), .B (n_3041), .S0 (WX3237), .Y (n_3099));
MX2X1 g60861(.A (n_3027), .B (n_2945), .S0 (WX10993), .Y (n_3098));
MX2X1 g60866(.A (n_3027), .B (n_3072), .S0 (WX9710), .Y (n_3096));
MX2X1 g60867(.A (n_3027), .B (n_2945), .S0 (WX10995), .Y (n_3095));
MX2X1 g60868(.A (n_3027), .B (n_3072), .S0 (WX3239), .Y (n_3093));
MX2X1 g60874(.A (n_3027), .B (n_2945), .S0 (WX3241), .Y (n_3092));
MX2X1 g60875(.A (n_3058), .B (n_3089), .S0 (WX5863), .Y (n_3090));
MX2X1 g60877(.A (n_3021), .B (n_2945), .S0 (WX11003), .Y (n_3088));
MX2X1 g60884(.A (n_3021), .B (n_3086), .S0 (WX5819), .Y (n_3087));
MX2X1 g60885(.A (n_3120), .B (n_3072), .S0 (WX10997), .Y (n_3085));
DFFSRX1 WX7286_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2300), .Q (WX7286), .QN ());
DFFSRX1 WX4636_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1931), .Q (WX4636), .QN ());
MX2X1 g60897(.A (n_3120), .B (n_3072), .S0 (WX5823), .Y (n_3083));
DFFSRX1 WX11163_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2240), .Q (WX11163), .QN ());
MX2X1 g60900(.A (n_3027), .B (n_3041), .S0 (WX5825), .Y (n_3081));
MX2X1 g60910(.A (n_3027), .B (n_3072), .S0 (WX5829), .Y (n_3080));
MX2X1 g60911(.A (n_3137), .B (n_3041), .S0 (WX5817), .Y (n_3077));
MX2X1 g60912(.A (n_3137), .B (n_3086), .S0 (WX5831), .Y (n_3076));
MX2X1 g60916(.A (n_3137), .B (n_3072), .S0 (WX5833), .Y (n_3075));
DFFSRX1 _2267__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1515), .Q (_2267_), .QN ());
MX2X1 g60918(.A (n_3137), .B (n_3072), .S0 (WX3247), .Y (n_3074));
MX2X1 g60922(.A (n_3027), .B (n_2945), .S0 (WX5841), .Y (n_3071));
DFFSRX1 WX8601_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2015), .Q (WX8601), .QN ());
MX2X1 g60924(.A (n_3137), .B (n_2945), .S0 (WX5843), .Y (n_3069));
MX2X1 g60925(.A (n_3137), .B (n_3072), .S0 (WX8433), .Y (n_3068));
DFFSRX1 WX3365_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2201), .Q (WX3365), .QN ());
MX2X1 g60929(.A (n_3106), .B (n_2988), .S0 (WX5877), .Y (n_3066));
MX2X1 g60932(.A (n_3021), .B (n_3072), .S0 (WX11013), .Y (n_3065));
MX2X1 g60936(.A (n_3021), .B (n_3072), .S0 (WX11005), .Y (n_3064));
DFFSRX1 WX2092_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1801), .Q (WX2092), .QN ());
MX2X1 g60946(.A (n_3106), .B (n_3089), .S0 (WX5861), .Y (n_3062));
MX2X1 g60948(.A (n_3021), .B (n_3072), .S0 (WX8427), .Y (n_3061));
MX2X1 g60952(.A (n_3058), .B (n_2953), .S0 (WX5865), .Y (n_3059));
MX2X1 g60953(.A (n_2829), .B (n_3056), .S0 (WX4574), .Y (n_3057));
MX2X1 g60954(.A (n_3021), .B (n_2945), .S0 (WX4542), .Y (n_3055));
MX2X1 g60958(.A (n_3021), .B (n_3041), .S0 (WX11009), .Y (n_3054));
MX2X1 g60960(.A (n_3137), .B (n_3041), .S0 (WX3253), .Y (n_3052));
DFFSRX1 WX2086_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1885), .Q (WX2086), .QN ());
MX2X1 g60962(.A (n_3137), .B (n_2938), .S0 (WX3259), .Y (n_3051));
MX2X1 g60967(.A (n_3120), .B (n_2945), .S0 (WX11011), .Y (n_3049));
DFFSRX1 WX2150_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2080), .Q (WX2150), .QN ());
DFFSRX1 WX11125_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1988), .Q (WX11125), .QN ());
MX2X1 g60980(.A (n_2986), .B (n_3056), .S0 (WX11035), .Y (n_3048));
MX2X1 g60983(.A (n_3120), .B (n_3072), .S0 (WX11015), .Y (n_3047));
MX2X1 g60989(.A (n_2829), .B (n_3044), .S0 (WX3265), .Y (n_3045));
DFFSRX1 WX3385_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2205), .Q (WX3385), .QN ());
DFFSRX1 WX7336_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2197), .Q (WX7336), .QN ());
DFFSRX1 WX2138_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1948), .Q (WX2138), .QN ());
MX2X1 g60992(.A (n_6423), .B (n_3041), .S0 (WX3245), .Y (n_3043));
MX2X1 g60993(.A (n_3137), .B (n_3072), .S0 (WX7140), .Y (n_3040));
MX2X1 g60994(.A (n_3137), .B (n_3041), .S0 (WX3261), .Y (n_3039));
DFFSRX1 WX7332_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1999), .Q (WX7332), .QN ());
MX2X1 g61003(.A (n_7483), .B (n_3072), .S0 (WX7110), .Y (n_3038));
MX2X1 g61004(.A (n_3058), .B (n_2828), .S0 (WX3267), .Y (n_3037));
MX2X1 g61009(.A (n_3031), .B (n_3072), .S0 (WX7112), .Y (n_3034));
MX2X1 g61014(.A (n_3031), .B (n_3086), .S0 (WX7114), .Y (n_3032));
MX2X1 g61018(.A (n_3031), .B (n_2945), .S0 (WX7116), .Y (n_3030));
MX2X1 g61023(.A (n_3027), .B (n_3072), .S0 (WX5835), .Y (n_3029));
MX2X1 g61024(.A (n_3027), .B (n_3086), .S0 (WX11019), .Y (n_3028));
MX2X1 g61026(.A (n_7483), .B (n_3072), .S0 (WX7118), .Y (n_3026));
MX2X1 g61031(.A (n_7483), .B (n_3041), .S0 (WX7120), .Y (n_3024));
MX2X1 g61037(.A (n_3021), .B (n_3072), .S0 (WX7122), .Y (n_3023));
MX2X1 g61039(.A (n_3021), .B (n_3072), .S0 (WX5827), .Y (n_3022));
MX2X1 g61041(.A (n_3021), .B (n_3041), .S0 (WX7124), .Y (n_3020));
MX2X1 g61045(.A (n_3021), .B (n_3041), .S0 (WX7126), .Y (n_3018));
MX2X1 g61046(.A (n_3021), .B (n_7488), .S0 (WX9720), .Y (n_3017));
MX2X1 g61049(.A (n_3021), .B (n_3086), .S0 (WX5837), .Y (n_3015));
MX2X1 g61053(.A (n_3021), .B (n_3072), .S0 (WX7128), .Y (n_3014));
DFFSRX1 WX9920_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2299), .Q (WX9920), .QN ());
DFFSRX1 _2304__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1509), .Q (_2304_), .QN ());
DFFSRX1 WX8605_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1913), .Q (WX8605), .QN ());
MX2X1 g61059(.A (n_3027), .B (n_3086), .S0 (WX7130), .Y (n_3012));
MX2X1 g61060(.A (n_2986), .B (n_3044), .S0 (WX3273), .Y (n_3011));
MX2X1 g61067(.A (n_3027), .B (n_3072), .S0 (WX7132), .Y (n_3009));
DFFSRX1 _2117__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1510), .Q (_2117_), .QN ());
MX2X1 g61070(.A (n_3058), .B (n_2993), .S0 (WX3275), .Y (n_3007));
MX2X1 g61071(.A (n_2776), .B (n_3004), .S0 (WX11023), .Y (n_3005));
MX2X1 g61072(.A (n_3021), .B (n_3072), .S0 (WX7134), .Y (n_3003));
MX2X1 g61076(.A (n_3021), .B (n_3041), .S0 (WX9718), .Y (n_3001));
MX2X1 g61077(.A (n_3021), .B (n_3086), .S0 (WX7136), .Y (n_3000));
MX2X1 g61082(.A (n_3021), .B (n_3072), .S0 (WX7138), .Y (n_2999));
MX2X1 g61087(.A (n_3106), .B (n_2817), .S0 (WX4584), .Y (n_2998));
MX2X1 g61094(.A (n_3058), .B (n_2996), .S0 (WX7142), .Y (n_2997));
MX2X1 g61099(.A (n_3106), .B (n_3105), .S0 (WX7144), .Y (n_2995));
MX2X1 g61104(.A (n_2813), .B (n_2993), .S0 (WX7146), .Y (n_2994));
MX2X1 g61108(.A (n_3106), .B (n_2770), .S0 (WX7148), .Y (n_2992));
DFFSRX1 WX7242_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1807), .Q (WX7242), .QN ());
DFFSRX1 _2341__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1529), .Q (_2341_), .QN ());
MX2X1 g61112(.A (n_2986), .B (n_2996), .S0 (WX7150), .Y (n_2991));
MX2X1 g61126(.A (n_3058), .B (n_2988), .S0 (WX7156), .Y (n_2990));
DFFSRX1 _2153__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1691), .Q (_2153_), .QN ());
MX2X1 g61127(.A (n_2986), .B (n_3103), .S0 (WX3281), .Y (n_2987));
MX2X1 g61129(.A (n_6513), .B (n_3004), .S0 (WX7158), .Y (n_2985));
MX2X1 g61131(.A (n_2798), .B (n_3103), .S0 (WX11029), .Y (n_2984));
MX2X1 g61132(.A (n_2986), .B (n_2993), .S0 (WX8449), .Y (n_2982));
DFFSRX1 _2190__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1611), .Q (_2190_), .QN ());
DFFSRX1 WX8633_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1986), .Q (WX8633), .QN ());
MX2X1 g61139(.A (n_3106), .B (n_2755), .S0 (WX7162), .Y (n_2981));
MX2X1 g61147(.A (n_3106), .B (n_3056), .S0 (WX7166), .Y (n_2979));
MX2X1 g61149(.A (n_2829), .B (n_2976), .S0 (WX3285), .Y (n_2978));
MX2X1 g61150(.A (n_3058), .B (n_2755), .S0 (WX11031), .Y (n_2975));
DFFSRX1 WX9916_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2392), .Q (WX9916), .QN ());
DFFSRX1 WX8493_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1964), .Q (WX8493), .QN ());
MX2X1 g61166(.A (n_3058), .B (n_2795), .S0 (WX7172), .Y (n_2974));
MX2X1 g61169(.A (n_3021), .B (n_3072), .S0 (WX9716), .Y (n_2972));
MX2X1 g61171(.A (n_3058), .B (n_2755), .S0 (WX11033), .Y (n_2971));
DFFSRX1 WX3345_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2179), .Q (WX3345), .QN ());
MX2X1 g61187(.A (n_3137), .B (n_3072), .S0 (WX3243), .Y (n_2969));
MX2X1 g61188(.A (n_3058), .B (n_3044), .S0 (WX11037), .Y (n_2968));
MX2X1 g61189(.A (n_3058), .B (n_2988), .S0 (WX3293), .Y (n_2967));
MX2X1 g61197(.A (n_3058), .B (n_2795), .S0 (WX11039), .Y (n_2966));
DFFSRX1 WX9790_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2253), .Q (WX9790), .QN ());
DFFSRX1 WX9794_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2231), .Q (WX9794), .QN ());
MX2X1 g61212(.A (n_3137), .B (n_3072), .S0 (WX8405), .Y (n_2965));
MX2X1 g61215(.A (n_3137), .B (n_2938), .S0 (WX8407), .Y (n_2963));
DFFSRX1 WX9868_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1965), .Q (WX9868), .QN ());
MX2X1 g61218(.A (n_3021), .B (n_2938), .S0 (WX8409), .Y (n_2961));
DFFSRX1 _2231__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1584), .Q (_2231_), .QN ());
MX2X1 g61221(.A (n_3021), .B (n_2938), .S0 (WX8411), .Y (n_2960));
DFFSRX1 _2310__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1551), .Q (_2310_), .QN ());
MX2X1 g61225(.A (n_3137), .B (n_2945), .S0 (WX11001), .Y (n_2958));
MX2X1 g61226(.A (n_3137), .B (n_3041), .S0 (WX5821), .Y (n_2957));
DFFSRX1 WX9824_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2129), .Q (WX9824), .QN ());
MX2X1 g61228(.A (n_3021), .B (n_3072), .S0 (WX10999), .Y (n_2955));
MX2X1 g61238(.A (n_3058), .B (n_2953), .S0 (WX9732), .Y (n_2954));
MX2X1 g61244(.A (n_3137), .B (n_3072), .S0 (WX8421), .Y (n_2952));
DFFSRX1 WX9832_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2124), .Q (WX9832), .QN ());
MX2X1 g61248(.A (n_3137), .B (n_3072), .S0 (WX8423), .Y (n_2950));
DFFSRX1 WX11175_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2379), .Q (WX11175), .QN ());
DFFSRX1 WX3311_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2178), .Q (WX3311), .QN ());
MX2X1 g61252(.A (n_3140), .B (n_2938), .S0 (WX8425), .Y (n_2949));
MX2X1 g61259(.A (n_3137), .B (n_3072), .S0 (WX4526), .Y (n_2948));
DFFSRX1 WX2134_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1895), .Q (WX2134), .QN ());
MX2X1 g61266(.A (n_3137), .B (n_2938), .S0 (WX8429), .Y (n_2947));
MX2X1 g61269(.A (n_3021), .B (n_2945), .S0 (WX8431), .Y (n_2946));
MX2X1 g61272(.A (n_3021), .B (n_3041), .S0 (WX4528), .Y (n_2944));
MX2X1 g61277(.A (n_3021), .B (n_2945), .S0 (WX9714), .Y (n_2943));
MX2X1 g61278(.A (n_3021), .B (n_2945), .S0 (WX4530), .Y (n_2941));
DFFSRX1 _2229__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1587), .Q (_2229_), .QN ());
MX2X1 g61283(.A (n_2809), .B (n_3004), .S0 (WX8437), .Y (n_2940));
DFFSRX1 WX11121_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1974), .Q (WX11121), .QN ());
MX2X1 g61287(.A (n_3021), .B (n_2938), .S0 (WX4532), .Y (n_2939));
MX2X1 g61291(.A (n_3106), .B (n_2993), .S0 (WX8441), .Y (n_2937));
DFFSRX1 _2192__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1608), .Q (_2192_), .QN ());
MX2X1 g61293(.A (n_2935), .B (n_2976), .S0 (WX9736), .Y (n_2936));
MX2X1 g61294(.A (n_3021), .B (n_2938), .S0 (WX4534), .Y (n_2934));
MX2X1 g61296(.A (n_3106), .B (n_2976), .S0 (WX8445), .Y (n_2933));
MX2X1 g61299(.A (n_3137), .B (n_2938), .S0 (WX4536), .Y (n_2932));
MX2X1 g61305(.A (n_3031), .B (n_2945), .S0 (WX4538), .Y (n_2931));
MX2X1 g61308(.A (n_6513), .B (n_2996), .S0 (WX5857), .Y (n_2930));
NOR2X1 g61336(.A (WX10829), .B (n_2849), .Y (n_2928));
NOR2X1 g61341(.A (n_2849), .B (WX485), .Y (n_2927));
DFFSRX1 WX9826_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2312), .Q (WX9826), .QN ());
DFFSRX1 WX8575_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1904), .Q (WX8575), .QN ());
DFFSRX1 WX2108_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1750), .Q (WX2108), .QN ());
INVX2 g61376(.A (n_2926), .Y (n_5493));
INVX2 g61377(.A (n_2926), .Y (n_5183));
INVX1 g61378(.A (n_2926), .Y (n_5085));
INVX2 g61379(.A (n_2926), .Y (n_4803));
INVX1 g61380(.A (n_2926), .Y (n_5254));
INVX1 g61385(.A (n_2925), .Y (n_5474));
INVX1 g61386(.A (n_2925), .Y (n_5600));
INVX1 g61387(.A (n_2925), .Y (n_5918));
INVX1 g61388(.A (n_2925), .Y (n_5320));
INVX1 g61389(.A (n_2925), .Y (n_5598));
INVX1 g61390(.A (n_2925), .Y (n_5239));
INVX1 g61391(.A (n_2925), .Y (n_4866));
INVX1 g61392(.A (n_2925), .Y (n_5549));
INVX2 g61395(.A (n_2924), .Y (n_5415));
INVX2 g61396(.A (n_2924), .Y (n_5928));
INVX1 g61397(.A (n_2924), .Y (n_5196));
DFFSRX1 WX3415_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2275), .Q (WX3415), .QN ());
INVX1 g61398(.A (n_2924), .Y (n_5317));
INVX1 g61399(.A (n_2924), .Y (n_4868));
INVX1 g61400(.A (n_2924), .Y (n_5630));
INVX1 g61404(.A (n_6482), .Y (n_5750));
INVX1 g61405(.A (n_6482), .Y (n_5334));
INVX4 g61406(.A (n_6482), .Y (n_5439));
INVX1 g61408(.A (n_6482), .Y (n_5649));
INVX1 g61410(.A (n_6482), .Y (n_5158));
INVX8 g61418(.A (n_2922), .Y (n_4697));
INVX2 g61421(.A (n_2921), .Y (n_5235));
INVX1 g61422(.A (n_2921), .Y (n_5576));
INVX1 g61424(.A (n_2921), .Y (n_5886));
INVX1 g61425(.A (n_2921), .Y (n_5845));
INVX1 g61426(.A (n_2921), .Y (n_5729));
INVX1 g61427(.A (n_2921), .Y (n_5418));
INVX1 g61428(.A (n_2921), .Y (n_5482));
INVX1 g61430(.A (n_7090), .Y (n_5393));
INVX1 g61432(.A (n_7090), .Y (n_5882));
INVX1 g61433(.A (n_7090), .Y (n_5185));
INVX4 g61435(.A (n_7090), .Y (n_5841));
INVX1 g61437(.A (n_7090), .Y (n_6106));
INVX4 g61440(.A (n_6503), .Y (n_5535));
INVX2 g61441(.A (n_6503), .Y (n_5468));
INVX1 g61444(.A (n_6503), .Y (n_5830));
INVX1 g61445(.A (n_6503), .Y (n_6050));
INVX1 g61446(.A (n_6503), .Y (n_5490));
INVX2 g61448(.A (n_2920), .Y (n_5879));
INVX1 g61451(.A (n_2920), .Y (n_5825));
INVX2 g61452(.A (n_2920), .Y (n_5105));
INVX2 g61454(.A (n_2920), .Y (n_5892));
INVX1 g61455(.A (n_2920), .Y (n_5834));
DFFSRX1 _2144__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1645), .Q (_2144_), .QN ());
NOR2X1 g61468(.A (WX1778), .B (n_2849), .Y (n_2917));
DFFSRX1 WX6065_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1962), .Q (WX6065), .QN ());
DFFSRX1 WX5997_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2323), .Q (WX5997), .QN ());
DFFSRX1 _2187__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1613), .Q (_2187_), .QN ());
DFFSRX1 WX9944_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1977), .Q (WX9944), .QN ());
DFFSRX1 WX6017_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2353), .Q (WX6017), .QN ());
DFFSRX1 WX3451_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2010), .Q (WX3451), .QN ());
DFFSRX1 WX7190_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2176), .Q (WX7190), .QN ());
DFFSRX1 WX8655_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2110), .Q (WX8655), .QN ());
DFFSRX1 WX7278_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2290), .Q (WX7278), .QN ());
DFFSRX1 WX7232_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1840), .Q (WX7232), .QN ());
DFFSRX1 WX9774_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1671), .Q (WX9774), .QN ());
DFFSRX1 WX8597_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1485), .Q (WX8597), .QN ());
DFFSRX1 WX9860_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2133), .Q (WX9860), .QN ());
DFFSRX1 WX11229_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1791), .Q (WX11229), .QN ());
NOR2X1 g61699(.A (n_2849), .B (n_920), .Y (n_2916));
NOR2X1 g61737(.A (n_2849), .B (n_935), .Y (n_2914));
NOR2X1 g61760(.A (n_2849), .B (n_126), .Y (n_2912));
DFFSRX1 WX8653_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2116), .Q (WX8653), .QN ());
DFFSRX1 WX6053_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1959), .Q (WX6053), .QN ());
NOR2X1 g61771(.A (n_2849), .B (n_85), .Y (n_2911));
DFFSRX1 WX3485_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2363), .Q (WX3485), .QN ());
NOR2X1 g61774(.A (n_2849), .B (n_120), .Y (n_2909));
NOR2X1 g61775(.A (n_2849), .B (n_40), .Y (n_2908));
DFFSRX1 WX9782_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2120), .Q (WX9782), .QN ());
NOR2X1 g61806(.A (n_2849), .B (n_977), .Y (n_2907));
NOR2X1 g61808(.A (n_2849), .B (n_5), .Y (n_2906));
DFFSRX1 WX8619_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2054), .Q (WX8619), .QN ());
DFFSRX1 WX3471_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2057), .Q (WX3471), .QN ());
DFFSRX1 WX6021_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2142), .Q (WX6021), .QN ());
DFFSRX1 WX2100_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2408), .Q (WX2100), .QN ());
DFFSRX1 WX6049_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2258), .Q (WX6049), .QN ());
DFFSRX1 WX2078_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1754), .Q (WX2078), .QN ());
DFFSRX1 WX4666_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2027), .Q (WX4666), .QN ());
DFFSRX1 _2261__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1620), .Q (_2261_), .QN ());
DFFSRX1 _2300__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1552), .Q (_2300_), .QN ());
DFFSRX1 WX7236_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1765), .Q (WX7236), .QN ());
DFFSRX1 _2225__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1590), .Q (_2225_), .QN ());
DFFSRX1 WX5885_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1471), .Q (WX5885), .QN ());
DFFSRX1 WX8623_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2101), .Q (WX8623), .QN ());
NOR2X1 g62112(.A (n_2849), .B (n_927), .Y (n_2905));
NOR2X1 g62114(.A (n_2849), .B (n_924), .Y (n_2903));
DFFSRX1 WX5903_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1738), .Q (WX5903), .QN ());
DFFSRX1 WX4630_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2061), .Q (WX4630), .QN ());
DFFSRX1 WX3399_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2073), .Q (WX3399), .QN ());
DFFSRX1 WX11113_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2394), .Q (WX11113), .QN ());
NOR2X1 g62151(.A (n_2849), .B (n_33), .Y (n_2902));
DFFSRX1 WX6001_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2175), .Q (WX6001), .QN ());
DFFSRX1 WX4592_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1788), .Q (WX4592), .QN ());
DFFSRX1 WX5907_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1787), .Q (WX5907), .QN ());
DFFSRX1 WX5955_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1825), .Q (WX5955), .QN ());
DFFSRX1 WX2082_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1814), .Q (WX2082), .QN ());
DFFSRX1 WX2074_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2117), .Q (WX2074), .QN ());
DFFSRX1 WX8591_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1710), .Q (WX8591), .QN ());
DFFSRX1 WX8567_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1813), .Q (WX8567), .QN ());
DFFSRX1 WX3419_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2160), .Q (WX3419), .QN ());
DFFSRX1 WX7302_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2559), .Q (WX7302), .QN ());
DFFSRX1 WX8565_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1873), .Q (WX8565), .QN ());
DFFSRX1 WX9902_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2068), .Q (WX9902), .QN ());
BUFX3 g62443(.A (n_7086), .Y (n_3183));
DFFSRX1 WX4588_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1883), .Q (WX4588), .QN ());
DFFSRX1 WX9820_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1955), .Q (WX9820), .QN ());
DFFSRX1 WX8539_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2442), .Q (WX8539), .QN ());
DFFSRX1 WX11109_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1483), .Q (WX11109), .QN ());
DFFSRX1 WX8537_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2369), .Q (WX8537), .QN ());
DFFSRX1 WX5979_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1878), .Q (WX5979), .QN ());
DFFSRX1 WX3347_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2167), .Q (WX3347), .QN ());
DFFSRX1 WX4750_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2074), .Q (WX4750), .QN ());
DFFSRX1 WX8467_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1833), .Q (WX8467), .QN ());
DFFSRX1 WX5931_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2136), .Q (WX5931), .QN ());
DFFSRX1 WX8501_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1875), .Q (WX8501), .QN ());
NOR2X1 g62618(.A (n_2825), .B (n_2849), .Y (n_2900));
DFFSRX1 WX3295_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1993), .Q (WX3295), .QN ());
DFFSRX1 _2111__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1668), .Q (_2111_), .QN ());
DFFSRX1 WX3319_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2228), .Q (WX3319), .QN ());
DFFSRX1 _2336__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1534), .Q (_2336_), .QN ());
DFFSRX1 _2147__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1644), .Q (_2147_), .QN ());
DFFSRX1 _2114__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1665), .Q (_2114_), .QN ());
DFFSRX1 WX4726_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2123), .Q (WX4726), .QN ());
DFFSRX1 WX3359_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2053), .Q (WX3359), .QN ());
DFFSRX1 WX4634_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2147), .Q (WX4634), .QN ());
DFFSRX1 WX4682_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1996), .Q (WX4682), .QN ());
DFFSRX1 WX11105_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1481), .Q (WX11105), .QN ());
DFFSRX1 WX3307_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2113), .Q (WX3307), .QN ());
DFFSRX1 WX3313_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1837), .Q (WX3313), .QN ());
DFFSRX1 WX3351_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2141), .Q (WX3351), .QN ());
DFFSRX1 _2339__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1531), .Q (_2339_), .QN ());
DFFSRX1 WX3431_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1989), .Q (WX3431), .QN ());
DFFSRX1 WX3379_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1896), .Q (WX3379), .QN ());
DFFSRX1 WX3299_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2095), .Q (WX3299), .QN ());
DFFSRX1 WX3303_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2109), .Q (WX3303), .QN ());
DFFSRX1 WX3355_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1717), .Q (WX3355), .QN ());
DFFSRX1 _2138__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1650), .Q (_2138_), .QN ());
DFFSRX1 WX8559_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1877), .Q (WX8559), .QN ());
DFFSRX1 WX3459_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2127), .Q (WX3459), .QN ());
DFFSRX1 WX6057_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1958), .Q (WX6057), .QN ());
DFFSRX1 WX8531_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1969), .Q (WX8531), .QN ());
DFFSRX1 WX8579_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1762), .Q (WX8579), .QN ());
DFFSRX1 WX4762_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2111), .Q (WX4762), .QN ());
DFFSRX1 _2219__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1693), .Q (_2219_), .QN ());
DFFSRX1 WX7248_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1792), .Q (WX7248), .QN ());
DFFSRX1 WX8589_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1991), .Q (WX8589), .QN ());
DFFSRX1 WX4626_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2274), .Q (WX4626), .QN ());
DFFSRX1 _2142__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1647), .Q (_2142_), .QN ());
DFFSRX1 WX7262_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1491), .Q (WX7262), .QN ());
DFFSRX1 _2252__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1498), .Q (_2252_), .QN ());
DFFSRX1 WX9852_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2070), .Q (WX9852), .QN ());
DFFSRX1 _2361__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1517), .Q (_2361_), .QN ());
DFFSRX1 _2109__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1670), .Q (_2109_), .QN ());
DFFSRX1 WX9806_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2170), .Q (WX9806), .QN ());
DFFSRX1 WX7268_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2356), .Q (WX7268), .QN ());
NOR2X1 g57537(.A (n_1473), .B (n_5181), .Y (n_2898));
DFFSRX1 _2215__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1593), .Q (_2215_), .QN ());
DFFSRX1 WX7180_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2134), .Q (WX7180), .QN ());
DFFSRX1 WX7364_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1980), .Q (WX7364), .QN ());
BUFX3 g63072(.A (n_4562), .Y (n_4593));
DFFSRX1 WX9940_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2390), .Q (WX9940), .QN ());
BUFX3 g63075(.A (n_4562), .Y (n_4644));
BUFX3 g63080(.A (n_6626), .Y (n_4096));
DFFSRX1 _2313__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1550), .Q (_2313_), .QN ());
DFFSRX1 WX9894_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2071), .Q (WX9894), .QN ());
BUFX3 g63147(.A (n_3162), .Y (n_3225));
INVX4 g63153(.A (n_2897), .Y (n_5965));
INVX4 g63155(.A (n_2897), .Y (n_6091));
BUFX3 g63159(.A (n_6437), .Y (n_4184));
BUFX3 g63181(.A (n_6437), .Y (n_5828));
BUFX3 g63187(.A (n_6452), .Y (n_4099));
BUFX3 g63215(.A (n_2894), .Y (n_4078));
BUFX3 g63217(.A (n_2894), .Y (n_4016));
DFFSRX1 WX6061_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2243), .Q (WX6061), .QN ());
DFFSRX1 WX9836_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2277), .Q (WX9836), .QN ());
DFFSRX1 WX6033_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1912), .Q (WX6033), .QN ());
DFFSRX1 WX6041_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1920), .Q (WX6041), .QN ());
DFFSRX1 WX6037_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1797), .Q (WX6037), .QN ());
DFFSRX1 WX11223_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1990), .Q (WX11223), .QN ());
DFFSRX1 WX8545_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1724), .Q (WX8545), .QN ());
DFFSRX1 WX7184_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2182), .Q (WX7184), .QN ());
DFFSRX1 WX7326_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1489), .Q (WX7326), .QN ());
DFFSRX1 _2180__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1617), .Q (_2180_), .QN ());
DFFSRX1 WX9798_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1848), .Q (WX9798), .QN ());
NOR2X1 g59247(.A (n_2535), .B (n_1648), .Y (n_2893));
NOR2X1 g59258(.A (n_1235), .B (n_2605), .Y (n_2892));
DFFSRX1 WX11187_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2276), .Q (WX11187), .QN ());
DFFSRX1 WX8523_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1772), .Q (WX8523), .QN ());
NOR2X1 g59262(.A (n_1026), .B (n_2849), .Y (n_2889));
INVX1 g55889(.A (WX487), .Y (n_2888));
DFFSRX1 WX7224_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2364), .Q (WX7224), .QN ());
DFFSRX1 _2129__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1504), .Q (_2129_), .QN ());
DFFSRX1 WX7228_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2350), .Q (WX7228), .QN ());
DFFSRX1 WX7270_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1719), .Q (WX7270), .QN ());
NOR2X1 g59268(.A (n_2546), .B (n_1648), .Y (n_2887));
NOR2X1 g59269(.A (n_2523), .B (n_1425), .Y (n_2885));
NOR2X1 g59270(.A (n_2545), .B (n_1425), .Y (n_2884));
NOR2X1 g59271(.A (n_2524), .B (n_5181), .Y (n_2883));
DFFSRX1 WX4700_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2154), .Q (WX4700), .QN ());
NOR2X1 g59272(.A (n_2517), .B (n_1425), .Y (n_2882));
DFFSRX1 WX5899_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1784), .Q (WX5899), .QN ());
NOR2X1 g59273(.A (n_2519), .B (n_1425), .Y (n_2881));
NOR2X1 g59274(.A (n_2542), .B (n_1425), .Y (n_2879));
NOR2X1 g59275(.A (n_2541), .B (n_5181), .Y (n_2878));
NOR2X1 g59276(.A (n_2539), .B (n_2849), .Y (n_2876));
NOR2X1 g59277(.A (n_2516), .B (n_1425), .Y (n_2875));
NOR2X1 g59278(.A (n_2551), .B (n_2849), .Y (n_2873));
NOR2X1 g59279(.A (n_2536), .B (n_1425), .Y (n_2872));
NOR2X1 g59280(.A (n_2518), .B (n_5181), .Y (n_2870));
NOR2X1 g59281(.A (n_2547), .B (n_1425), .Y (n_2868));
NOR2X1 g59282(.A (n_2557), .B (n_1425), .Y (n_2867));
NOR2X1 g59283(.A (n_2532), .B (n_1425), .Y (n_2866));
NOR2X1 g59284(.A (n_2548), .B (n_2849), .Y (n_2865));
DFFSRX1 WX7274_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1721), .Q (WX7274), .QN ());
NOR2X1 g59285(.A (n_2531), .B (n_5712), .Y (n_2864));
NOR2X1 g59286(.A (n_2552), .B (n_5712), .Y (n_2863));
NOR2X1 g59293(.A (n_1029), .B (n_2605), .Y (n_2861));
DFFSRX1 _2277__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1563), .Q (_2277_), .QN ());
DFFSRX1 WX9936_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2151), .Q (WX9936), .QN ());
DFFSRX1 WX5987_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2248), .Q (WX5987), .QN ());
DFFSRX1 WX2130_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2226), .Q (), .QN (WX2130));
NOR2X1 g59338(.A (n_1167), .B (n_2605), .Y (n_2860));
NOR2X1 g59339(.A (n_1234), .B (n_2605), .Y (n_2859));
DFFSRX1 WX11159_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2553), .Q (WX11159), .QN ());
DFFSRX1 WX3375_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1741), .Q (WX3375), .QN ());
DFFSRX1 WX3443_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2322), .Q (WX3443), .QN ());
DFFSRX1 WX7318_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1785), .Q (WX7318), .QN ());
DFFSRX1 WX8585_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1961), .Q (WX8585), .QN ());
DFFSRX1 WX8647_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2107), .Q (WX8647), .QN ());
DFFSRX1 WX9760_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2062), .Q (WX9760), .QN ());
DFFSRX1 WX5963_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2020), .Q (WX5963), .QN ());
DFFSRX1 WX8617_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2046), .Q (WX8617), .QN ());
DFFSRX1 WX3411_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2173), .Q (WX3411), .QN ());
NOR2X1 g59396(.A (n_1121), .B (n_2849), .Y (n_2858));
NOR2X1 g59397(.A (n_1222), .B (n_2849), .Y (n_2857));
DFFSRX1 WX5993_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2344), .Q (WX5993), .QN ());
DFFSRX1 WX8611_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2148), .Q (WX8611), .QN ());
DFFSRX1 WX11157_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2366), .Q (WX11157), .QN ());
DFFSRX1 WX11145_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2528), .Q (WX11145), .QN ());
DFFSRX1 WX9848_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1820), .Q (WX9848), .QN ());
DFFSRX1 WX11171_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2285), .Q (WX11171), .QN ());
DFFSRX1 WX7176_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1898), .Q (WX7176), .QN ());
DFFSRX1 _2257__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1507), .Q (_2257_), .QN ());
DFFSRX1 _2324__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1540), .Q (_2324_), .QN ());
DFFSRX1 _2330__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1535), .Q (_2330_), .QN ());
NOR2X1 g59466(.A (n_2521), .B (n_5712), .Y (n_2856));
NOR2X1 g59467(.A (n_2555), .B (n_5712), .Y (n_2855));
DFFSRX1 WX9766_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2391), .Q (WX9766), .QN ());
NOR2X1 g59470(.A (n_2533), .B (n_5181), .Y (n_2854));
DFFSRX1 _2297__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1690), .Q (_2297_), .QN ());
DFFSRX1 WX9802_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1889), .Q (WX9802), .QN ());
NOR2X1 g59479(.A (n_2538), .B (n_2851), .Y (n_2852));
NOR2X1 g59480(.A (n_2543), .B (n_2849), .Y (n_2850));
NOR2X1 g59481(.A (n_1043), .B (n_2849), .Y (n_2848));
DFFSRX1 WX7360_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2064), .Q (WX7360), .QN ());
NOR2X1 g59482(.A (n_1042), .B (n_2849), .Y (n_2847));
DFFSRX1 WX5971_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1838), .Q (WX5971), .QN ());
DFFSRX1 _2326__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1537), .Q (_2326_), .QN ());
NOR2X1 g59488(.A (n_2522), .B (n_5712), .Y (n_2846));
NOR2X1 g59491(.A (n_2520), .B (n_1648), .Y (n_2844));
NOR2X1 g59494(.A (n_2554), .B (n_5712), .Y (n_2843));
DFFSRX1 _2290__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1555), .Q (_2290_), .QN ());
DFFSRX1 WX3425_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2281), .Q (WX3425), .QN ());
DFFSRX1 _2291__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1554), .Q (_2291_), .QN ());
DFFSRX1 WX8645_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1729), .Q (WX8645), .QN ());
DFFSRX1 WX8527_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2041), .Q (WX8527), .QN ());
DFFSRX1 _2255__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1681), .Q (_2255_), .QN ());
DFFSRX1 WX6009_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2308), .Q (WX6009), .QN ());
DFFSRX1 WX3323_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2241), .Q (WX3323), .QN ());
DFFSRX1 _2133__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1654), .Q (_2133_), .QN ());
DFFSRX1 _2247__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1508), .Q (_2247_), .QN ());
DFFSRX1 _2283__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1559), .Q (_2283_), .QN ());
DFFSRX1 _2251__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1575), .Q (_2251_), .QN ());
DFFSRX1 _2137__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1514), .Q (_2137_), .QN ());
DFFSRX1 _2199__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1496), .Q (_2199_), .QN ());
DFFSRX1 WX3341_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2331), .Q (WX3341), .QN ());
DFFSRX1 _2320__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1545), .Q (_2320_), .QN ());
DFFSRX1 WX8487_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2303), .Q (WX8487), .QN ());
DFFSRX1 WX8477_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1984), .Q (WX8477), .QN ());
DFFSRX1 WX8511_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2166), .Q (WX8511), .QN ());
DFFSRX1 WX2066_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1493), .Q (WX2066), .QN ());
DFFSRX1 WX7254_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2264), .Q (WX7254), .QN ());
DFFSRX1 WX5939_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2270), .Q (WX5939), .QN ());
DFFSRX1 WX8639_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1725), .Q (WX8639), .QN ());
DFFSRX1 WX5947_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1847), .Q (WX5947), .QN ());
DFFSRX1 WX9906_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2207), .Q (WX9906), .QN ());
DFFSRX1 WX8513_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2221), .Q (WX8513), .QN ());
DFFSRX1 WX3337_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2309), .Q (WX3337), .QN ());
DFFSRX1 WX8475_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1972), .Q (WX8475), .QN ());
DFFSRX1 _2239__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1580), .Q (_2239_), .QN ());
DFFSRX1 WX9840_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2132), .Q (WX9840), .QN ());
DFFSRX1 WX4600_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1924), .Q (WX4600), .QN ());
DFFSRX1 WX4670_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1925), .Q (WX4670), .QN ());
DFFSRX1 WX7316_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2399), .Q (WX7316), .QN ());
DFFSRX1 WX8553_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1992), .Q (WX8553), .QN ());
DFFSRX1 WX11101_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2393), .Q (WX11101), .QN ());
DFFSRX1 WX3333_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1732), .Q (WX3333), .QN ());
DFFSRX1 WX10829_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2452), .Q (WX10829), .QN ());
DFFSRX1 WX5923_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2036), .Q (WX5923), .QN ());
DFFSRX1 WX8519_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2096), .Q (WX8519), .QN ());
DFFSRX1 WX8551_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1856), .Q (WX8551), .QN ());
DFFSRX1 _2359__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1519), .Q (_2359_), .QN ());
DFFSRX1 WX7344_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2237), .Q (WX7344), .QN ());
DFFSRX1 WX7352_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1901), .Q (WX7352), .QN ());
DFFSRX1 _2170__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1696), .Q (_2170_), .QN ());
DFFSRX1 WX7296_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2337), .Q (WX7296), .QN ());
DFFSRX1 _2172__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1624), .Q (_2172_), .QN ());
DFFSRX1 WX7212_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2206), .Q (WX7212), .QN ());
DFFSRX1 _2210__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1676), .Q (_2210_), .QN ());
DFFSRX1 _2214__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1594), .Q (_2214_), .QN ());
DFFSRX1 WX2116_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1818), .Q (WX2116), .QN ());
DFFSRX1 WX2070_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2011), .Q (WX2070), .QN ());
DFFSRX1 WX2184_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1935), .Q (WX2184), .QN ());
DFFSRX1 _2357__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1522), .Q (_2357_), .QN ());
DFFSRX1 _2173__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1623), .Q (_2173_), .QN ());
DFFSRX1 _2294__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1673), .Q (_2294_), .QN ());
DFFSRX1 _2364__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1706), .Q (_2364_), .QN ());
DFFSRX1 _2176__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1622), .Q (_2176_), .QN ());
DFFSRX1 _2243__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1579), .Q (_2243_), .QN ());
DFFSRX1 WX11117_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1495), .Q (WX11117), .QN ());
DFFSRX1 _2110__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1669), .Q (_2110_), .QN ());
DFFSRX1 _2112__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1666), .Q (_2112_), .QN ());
DFFSRX1 _2116__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1512), .Q (_2116_), .QN ());
DFFSRX1 _2115__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1664), .Q (_2115_), .QN ());
DFFSRX1 _2122__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1662), .Q (_2122_), .QN ());
DFFSRX1 _2123__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1661), .Q (_2123_), .QN ());
DFFSRX1 _2126__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1659), .Q (_2126_), .QN ());
DFFSRX1 _2128__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1656), .Q (_2128_), .QN ());
DFFSRX1 _2130__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1516), .Q (_2130_), .QN ());
DFFSRX1 _2132__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1655), .Q (_2132_), .QN ());
DFFSRX1 _2134__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1652), .Q (_2134_), .QN ());
DFFSRX1 _2136__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1651), .Q (_2136_), .QN ());
DFFSRX1 _2141__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1682), .Q (_2141_), .QN ());
DFFSRX1 _2143__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1646), .Q (_2143_), .QN ());
DFFSRX1 _2146__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1697), .Q (_2146_), .QN ());
DFFSRX1 _2148__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1642), .Q (_2148_), .QN ());
DFFSRX1 _2149__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1641), .Q (_2149_), .QN ());
DFFSRX1 _2151__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1640), .Q (_2151_), .QN ());
DFFSRX1 _2154__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1639), .Q (_2154_), .QN ());
DFFSRX1 _2155__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1638), .Q (_2155_), .QN ());
DFFSRX1 _2156__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1637), .Q (_2156_), .QN ());
DFFSRX1 _2159__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1635), .Q (_2159_), .QN ());
DFFSRX1 _2164__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1631), .Q (_2164_), .QN ());
DFFSRX1 _2165__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1629), .Q (_2165_), .QN ());
DFFSRX1 _2167__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1627), .Q (_2167_), .QN ());
DFFSRX1 _2169__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1625), .Q (_2169_), .QN ());
DFFSRX1 _2178__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1619), .Q (_2178_), .QN ());
DFFSRX1 _2179__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1618), .Q (_2179_), .QN ());
DFFSRX1 _2186__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1614), .Q (_2186_), .QN ());
DFFSRX1 _2188__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1612), .Q (_2188_), .QN ());
DFFSRX1 _2191__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1609), .Q (_2191_), .QN ());
DFFSRX1 _2193__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1607), .Q (_2193_), .QN ());
DFFSRX1 _2195__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1606), .Q (_2195_), .QN ());
DFFSRX1 _2200__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1603), .Q (_2200_), .QN ());
DFFSRX1 _2203__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1601), .Q (_2203_), .QN ());
DFFSRX1 _2284__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1558), .Q (_2284_), .QN ());
DFFSRX1 _2208__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1599), .Q (_2208_), .QN ());
DFFSRX1 _2211__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1598), .Q (_2211_), .QN ());
DFFSRX1 _2213__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1595), .Q (_2213_), .QN ());
DFFSRX1 _2217__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1592), .Q (_2217_), .QN ());
DFFSRX1 _2223__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1591), .Q (_2223_), .QN ());
DFFSRX1 _2222__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1687), .Q (_2222_), .QN ());
DFFSRX1 _2226__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1588), .Q (_2226_), .QN ());
DFFSRX1 _2227__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1568), .Q (_2227_), .QN ());
DFFSRX1 _2228__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1577), .Q (_2228_), .QN ());
DFFSRX1 _2230__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1585), .Q (_2230_), .QN ());
DFFSRX1 _2233__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1583), .Q (_2233_), .QN ());
DFFSRX1 _2234__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1506), .Q (_2234_), .QN ());
DFFSRX1 WX3371_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1946), .Q (WX3371), .QN ());
DFFSRX1 _2238__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1684), .Q (_2238_), .QN ());
DFFSRX1 _2245__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1649), .Q (_2245_), .QN ());
DFFSRX1 _2249__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1677), .Q (_2249_), .QN ());
DFFSRX1 _2254__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1574), .Q (_2254_), .QN ());
DFFSRX1 _2256__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1573), .Q (_2256_), .QN ());
DFFSRX1 _2259__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1572), .Q (_2259_), .QN ());
DFFSRX1 _2260__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1571), .Q (_2260_), .QN ());
DFFSRX1 _2266__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1567), .Q (_2266_), .QN ());
DFFSRX1 _2269__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1675), .Q (_2269_), .QN ());
DFFSRX1 _2274__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1576), .Q (_2274_), .QN ());
DFFSRX1 _2275__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1564), .Q (_2275_), .QN ());
DFFSRX1 _2279__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1561), .Q (_2279_), .QN ());
DFFSRX1 _2282__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1560), .Q (_2282_), .QN ());
DFFSRX1 _2288__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1685), .Q (_2288_), .QN ());
DFFSRX1 _2286__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1511), .Q (_2286_), .QN ());
DFFSRX1 _2299__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1553), .Q (_2299_), .QN ());
DFFSRX1 _2311__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1679), .Q (_2311_), .QN ());
DFFSRX1 _2314__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1502), .Q (_2314_), .QN ());
DFFSRX1 _2316__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1547), .Q (_2316_), .QN ());
DFFSRX1 _2321__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1544), .Q (_2321_), .QN ());
DFFSRX1 _2322__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1542), .Q (_2322_), .QN ());
DFFSRX1 _2323__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1541), .Q (_2323_), .QN ());
DFFSRX1 _2325__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1539), .Q (_2325_), .QN ());
DFFSRX1 _2329__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1536), .Q (_2329_), .QN ());
DFFSRX1 _2338__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1533), .Q (_2338_), .QN ());
DFFSRX1 _2340__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1530), .Q (_2340_), .QN ());
DFFSRX1 _2342__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1528), .Q (_2342_), .QN ());
DFFSRX1 _2343__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1527), .Q (_2343_), .QN ());
DFFSRX1 _2345__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1525), .Q (_2345_), .QN ());
DFFSRX1 _2356__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1523), .Q (_2356_), .QN ());
DFFSRX1 _2358__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1521), .Q (_2358_), .QN ());
DFFSRX1 _2360__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1518), .Q (_2360_), .QN ());
DFFSRX1 _2265__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1499), .Q (_2265_), .QN ());
DFFSRX1 WX11107_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2168), .Q (WX11107), .QN ());
DFFSRX1 WX11111_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1906), .Q (WX11111), .QN ());
DFFSRX1 WX11119_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1970), .Q (WX11119), .QN ());
DFFSRX1 WX11123_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2404), .Q (WX11123), .QN ());
DFFSRX1 WX11127_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2043), .Q (WX11127), .QN ());
DFFSRX1 WX11131_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2164), .Q (WX11131), .QN ());
DFFSRX1 WX11133_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1482), .Q (WX11133), .QN ());
DFFSRX1 WX11135_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2130), .Q (WX11135), .QN ());
DFFSRX1 WX11139_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1742), .Q (WX11139), .QN ());
DFFSRX1 WX11143_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2376), .Q (WX11143), .QN ());
DFFSRX1 WX7174_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2375), .Q (WX7174), .QN ());
DFFSRX1 WX7178_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2387), .Q (WX7178), .QN ());
DFFSRX1 WX11147_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2372), .Q (WX11147), .QN ());
DFFSRX1 WX7182_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2297), .Q (WX7182), .QN ());
DFFSRX1 WX11151_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2203), .Q (WX11151), .QN ());
DFFSRX1 WX7186_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2155), .Q (WX7186), .QN ());
DFFSRX1 WX7188_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2202), .Q (WX7188), .QN ());
DFFSRX1 WX7192_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2174), .Q (WX7192), .QN ());
DFFSRX1 WX11149_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2169), .Q (WX11149), .QN ());
DFFSRX1 WX7194_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2171), .Q (WX7194), .QN ());
DFFSRX1 WX7198_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2212), .Q (WX7198), .QN ());
DFFSRX1 WX7200_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2000), .Q (WX7200), .QN ());
DFFSRX1 WX7204_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1699), .Q (WX7204), .QN ());
DFFSRX1 WX11155_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1894), .Q (WX11155), .QN ());
DFFSRX1 WX7214_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2208), .Q (WX7214), .QN ());
DFFSRX1 WX7218_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2214), .Q (WX7218), .QN ());
DFFSRX1 WX7220_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2215), .Q (WX7220), .QN ());
DFFSRX1 WX7222_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2220), .Q (WX7222), .QN ());
DFFSRX1 WX7226_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1865), .Q (WX7226), .QN ());
DFFSRX1 WX7230_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2266), .Q (WX7230), .QN ());
DFFSRX1 WX7234_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1828), .Q (WX7234), .QN ());
DFFSRX1 WX11161_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1824), .Q (WX11161), .QN ());
DFFSRX1 WX7238_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1730), .Q (WX7238), .QN ());
DFFSRX1 WX7240_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1815), .Q (WX7240), .QN ());
DFFSRX1 WX11165_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1773), .Q (WX11165), .QN ());
DFFSRX1 WX7246_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2360), .Q (WX7246), .QN ());
DFFSRX1 WX7250_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2250), .Q (WX7250), .QN ());
DFFSRX1 WX7252_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1713), .Q (WX7252), .QN ());
DFFSRX1 WX11167_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2359), .Q (WX11167), .QN ());
DFFSRX1 WX7256_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2257), .Q (WX7256), .QN ());
DFFSRX1 WX7260_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2357), .Q (WX7260), .QN ());
DFFSRX1 WX7264_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1731), .Q (WX7264), .QN ());
DFFSRX1 WX7266_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1632), .Q (WX7266), .QN ());
DFFSRX1 WX11173_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2304), .Q (WX11173), .QN ());
DFFSRX1 WX7276_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2008), .Q (WX7276), .QN ());
DFFSRX1 WX7280_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1886), .Q (WX7280), .QN ());
DFFSRX1 WX7282_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2296), .Q (WX7282), .QN ());
DFFSRX1 WX7284_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2384), .Q (WX7284), .QN ());
DFFSRX1 WX7288_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2295), .Q (WX7288), .QN ());
DFFSRX1 WX7292_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2306), .Q (WX7292), .QN ());
DFFSRX1 WX11179_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2395), .Q (WX11179), .QN ());
DFFSRX1 WX7298_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2347), .Q (WX7298), .QN ());
DFFSRX1 WX11177_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2348), .Q (WX11177), .QN ());
DFFSRX1 WX7304_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2373), .Q (WX7304), .QN ());
DFFSRX1 WX7308_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2343), .Q (WX7308), .QN ());
DFFSRX1 WX7310_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2211), .Q (WX7310), .QN ());
DFFSRX1 WX7312_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2341), .Q (WX7312), .QN ());
DFFSRX1 WX7314_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2012), .Q (WX7314), .QN ());
DFFSRX1 WX11185_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2389), .Q (WX11185), .QN ());
DFFSRX1 WX7320_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2260), .Q (WX7320), .QN ());
DFFSRX1 WX7322_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1976), .Q (WX7322), .QN ());
DFFSRX1 WX7324_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1954), .Q (WX7324), .QN ());
DFFSRX1 WX7328_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1967), .Q (WX7328), .QN ());
DFFSRX1 WX11189_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1985), .Q (WX11189), .QN ());
DFFSRX1 WX7334_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1960), .Q (WX7334), .QN ());
DFFSRX1 WX7338_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1921), .Q (WX7338), .QN ());
DFFSRX1 WX7340_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2332), .Q (WX7340), .QN ());
DFFSRX1 WX11191_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1804), .Q (WX11191), .QN ());
DFFSRX1 WX7342_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2244), .Q (WX7342), .QN ());
DFFSRX1 WX7346_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2022), .Q (WX7346), .QN ());
DFFSRX1 WX11193_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1494), .Q (WX11193), .QN ());
DFFSRX1 WX7348_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1472), .Q (WX7348), .QN ());
DFFSRX1 WX7354_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1774), .Q (WX7354), .QN ());
DFFSRX1 WX7358_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2349), .Q (WX7358), .QN ());
DFFSRX1 WX4662_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2288), .Q (WX4662), .QN ());
DFFSRX1 WX11197_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2328), .Q (WX11197), .QN ());
DFFSRX1 WX11201_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2326), .Q (WX11201), .QN ());
DFFSRX1 WX11203_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2145), .Q (WX11203), .QN ());
DFFSRX1 WX11205_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2190), .Q (WX11205), .QN ());
DFFSRX1 WX11209_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1745), .Q (WX11209), .QN ());
DFFSRX1 WX11211_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2156), .Q (WX11211), .QN ());
DFFSRX1 WX7300_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1761), .Q (WX7300), .QN ());
DFFSRX1 WX11213_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2140), .Q (WX11213), .QN ());
DFFSRX1 WX11215_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1822), .Q (WX11215), .QN ());
DFFSRX1 WX11217_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2361), .Q (WX11217), .QN ());
DFFSRX1 WX11219_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1490), .Q (WX11219), .QN ());
DFFSRX1 WX4710_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1978), .Q (WX4710), .QN ());
DFFSRX1 WX11221_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1861), .Q (WX11221), .QN ());
DFFSRX1 WX11225_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2324), .Q (WX11225), .QN ());
DFFSRX1 WX11227_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2280), .Q (WX11227), .QN ());
DFFSRX1 WX11231_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1470), .Q (WX11231), .QN ());
DFFSRX1 WX11233_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2513), .Q (WX11233), .QN ());
DFFSRX1 WX4646_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1944), .Q (WX4646), .QN ());
DFFSRX1 WX11241_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2329), .Q (WX11241), .QN ());
DFFSRX1 WX11243_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1746), .Q (WX11243), .QN ());
DFFSRX1 WX4658_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2351), .Q (WX4658), .QN ());
DFFSRX1 WX3327_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2267), .Q (WX3327), .QN ());
DFFSRX1 WX3321_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2398), .Q (WX3321), .QN ());
DFFSRX1 WX4640_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2128), .Q (WX4640), .QN ());
DFFSRX1 WX4708_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1936), .Q (WX4708), .QN ());
DFFSRX1 WX7210_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1914), .Q (WX7210), .QN ());
DFFSRX1 WX3297_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2098), .Q (WX3297), .QN ());
DFFSRX1 WX3301_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2318), .Q (WX3301), .QN ());
DFFSRX1 WX3305_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2112), .Q (WX3305), .QN ());
DFFSRX1 WX3309_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2118), .Q (WX3309), .QN ());
DFFSRX1 WX3315_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1714), .Q (WX3315), .QN ());
DFFSRX1 WX3317_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2066), .Q (WX3317), .QN ());
DFFSRX1 WX3325_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1793), .Q (WX3325), .QN ());
DFFSRX1 WX3329_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2191), .Q (WX3329), .QN ());
DFFSRX1 WX3331_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2183), .Q (WX3331), .QN ());
DFFSRX1 WX3335_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2403), .Q (WX3335), .QN ());
DFFSRX1 WX3339_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2433), .Q (WX3339), .QN ());
DFFSRX1 WX3343_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2355), .Q (WX3343), .QN ());
DFFSRX1 WX3349_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2352), .Q (WX3349), .QN ());
DFFSRX1 WX3353_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2234), .Q (WX3353), .QN ());
DFFSRX1 WX7306_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2086), .Q (WX7306), .QN ());
DFFSRX1 WX3357_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1783), .Q (WX3357), .QN ());
DFFSRX1 WX3361_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2048), .Q (WX3361), .QN ());
DFFSRX1 WX3363_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2038), .Q (WX3363), .QN ());
DFFSRX1 WX8469_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2026), .Q (WX8469), .QN ());
DFFSRX1 WX8471_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2149), .Q (WX8471), .QN ());
DFFSRX1 WX8473_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1997), .Q (WX8473), .QN ());
DFFSRX1 WX3367_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1957), .Q (WX3367), .QN ());
DFFSRX1 WX8479_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1734), .Q (WX8479), .QN ());
DFFSRX1 WX11195_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2282), .Q (WX11195), .QN ());
DFFSRX1 WX8483_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1790), .Q (WX8483), .QN ());
DFFSRX1 WX3373_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1735), .Q (WX3373), .QN ());
DFFSRX1 WX8489_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1829), .Q (WX8489), .QN ());
DFFSRX1 WX8491_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1930), .Q (WX8491), .QN ());
DFFSRX1 WX3377_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1876), .Q (WX3377), .QN ());
DFFSRX1 WX8495_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1903), .Q (WX8495), .QN ());
DFFSRX1 WX8497_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1907), .Q (WX8497), .QN ());
DFFSRX1 WX8499_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2016), .Q (WX8499), .QN ());
DFFSRX1 WX3381_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1755), .Q (WX3381), .QN ());
DFFSRX1 WX8503_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1890), .Q (WX8503), .QN ());
DFFSRX1 WX8505_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2249), .Q (WX8505), .QN ());
DFFSRX1 WX3383_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2289), .Q (WX3383), .QN ());
DFFSRX1 WX8509_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2255), .Q (WX8509), .QN ());
DFFSRX1 WX3387_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1816), .Q (WX3387), .QN ());
DFFSRX1 WX8515_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1764), .Q (WX8515), .QN ());
DFFSRX1 WX3389_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1767), .Q (WX3389), .QN ());
DFFSRX1 WX8517_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2163), .Q (WX8517), .QN ());
DFFSRX1 WX3391_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2302), .Q (WX3391), .QN ());
DFFSRX1 WX3393_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1849), .Q (WX3393), .QN ());
DFFSRX1 _2135__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1513), .Q (_2135_), .QN ());
DFFSRX1 WX8525_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1850), .Q (WX8525), .QN ());
DFFSRX1 WX3395_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2039), .Q (WX3395), .QN ());
DFFSRX1 WX3397_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2004), .Q (WX3397), .QN ());
DFFSRX1 WX8535_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1775), .Q (WX8535), .QN ());
DFFSRX1 WX3403_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2530), .Q (WX3403), .QN ());
DFFSRX1 WX8541_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1880), .Q (WX8541), .QN ());
DFFSRX1 WX3405_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1817), .Q (WX3405), .QN ());
DFFSRX1 WX8547_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1947), .Q (WX8547), .QN ());
DFFSRX1 WX3407_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1899), .Q (WX3407), .QN ());
DFFSRX1 WX8549_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1726), .Q (WX8549), .QN ());
DFFSRX1 WX3409_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1853), .Q (WX3409), .QN ());
DFFSRX1 WX8555_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2370), .Q (WX8555), .QN ());
DFFSRX1 WX8557_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1860), .Q (WX8557), .QN ());
DFFSRX1 WX3413_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2362), .Q (WX3413), .QN ());
DFFSRX1 WX8561_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1863), .Q (WX8561), .QN ());
DFFSRX1 WX8563_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1867), .Q (WX8563), .QN ());
DFFSRX1 WX3417_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1933), .Q (WX3417), .QN ());
DFFSRX1 WX8569_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2558), .Q (WX8569), .QN ());
DFFSRX1 WX8571_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1918), .Q (WX8571), .QN ());
DFFSRX1 WX8573_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1908), .Q (WX8573), .QN ());
DFFSRX1 WX3421_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2180), .Q (WX3421), .QN ());
DFFSRX1 WX8577_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1909), .Q (WX8577), .QN ());
DFFSRX1 WX3423_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1492), .Q (WX3423), .QN ());
DFFSRX1 WX8581_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2279), .Q (WX8581), .QN ());
DFFSRX1 WX4706_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1998), .Q (WX4706), .QN ());
DFFSRX1 WX3427_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2242), .Q (WX3427), .QN ());
DFFSRX1 WX3429_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2283), .Q (WX3429), .QN ());
DFFSRX1 WX8593_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2224), .Q (WX8593), .QN ());
DFFSRX1 WX3435_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1973), .Q (WX3435), .QN ());
DFFSRX1 WX3437_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1911), .Q (WX3437), .QN ());
DFFSRX1 WX8603_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2031), .Q (WX8603), .QN ());
DFFSRX1 WX11183_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2177), .Q (WX11183), .QN ());
DFFSRX1 WX3441_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1893), .Q (WX3441), .QN ());
DFFSRX1 WX8613_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2037), .Q (WX8613), .QN ());
DFFSRX1 WX7258_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2256), .Q (WX7258), .QN ());
DFFSRX1 WX8615_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2152), .Q (WX8615), .QN ());
DFFSRX1 WX3445_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2262), .Q (WX3445), .QN ());
DFFSRX1 WX3447_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2102), .Q (WX3447), .QN ());
DFFSRX1 WX8621_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2139), .Q (WX8621), .QN ());
DFFSRX1 WX3449_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2083), .Q (WX3449), .QN ());
DFFSRX1 WX8625_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2077), .Q (WX8625), .QN ());
DFFSRX1 WX8627_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1736), .Q (WX8627), .QN ());
DFFSRX1 WX8629_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2104), .Q (WX8629), .QN ());
DFFSRX1 WX3453_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1698), .Q (WX3453), .QN ());
DFFSRX1 WX8635_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2090), .Q (WX8635), .QN ());
DFFSRX1 WX8637_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2093), .Q (WX8637), .QN ());
DFFSRX1 WX3457_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2097), .Q (WX3457), .QN ());
DFFSRX1 WX8641_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1708), .Q (WX8641), .QN ());
DFFSRX1 WX8643_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2103), .Q (WX8643), .QN ());
DFFSRX1 WX3461_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1981), .Q (WX3461), .QN ());
DFFSRX1 WX3463_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1776), .Q (WX3463), .QN ());
DFFSRX1 WX3465_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2045), .Q (WX3465), .QN ());
DFFSRX1 WX8657_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1975), .Q (WX8657), .QN ());
DFFSRX1 WX3467_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2397), .Q (WX3467), .QN ());
DFFSRX1 WX3469_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2119), .Q (WX3469), .QN ());
DFFSRX1 WX3473_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2200), .Q (WX3473), .QN ());
DFFSRX1 WX3475_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1864), .Q (WX3475), .QN ());
DFFSRX1 WX3477_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1718), .Q (WX3477), .QN ());
DFFSRX1 WX3479_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2229), .Q (WX3479), .QN ());
DFFSRX1 WX3481_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1919), .Q (WX3481), .QN ());
DFFSRX1 WX3483_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2034), .Q (WX3483), .QN ());
DFFSRX1 WX9876_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2059), .Q (WX9876), .QN ());
DFFSRX1 WX9904_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2137), .Q (WX9904), .QN ());
DFFSRX1 WX9764_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2042), .Q (WX9764), .QN ());
DFFSRX1 WX9928_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2084), .Q (WX9928), .QN ());
DFFSRX1 WX9762_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2284), .Q (WX9762), .QN ());
DFFSRX1 WX9768_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2252), .Q (WX9768), .QN ());
DFFSRX1 WX9770_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2114), .Q (WX9770), .QN ());
DFFSRX1 WX9772_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2556), .Q (WX9772), .QN ());
DFFSRX1 WX9776_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2345), .Q (WX9776), .QN ());
DFFSRX1 WX9778_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2475), .Q (WX9778), .QN ());
DFFSRX1 WX9780_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2316), .Q (WX9780), .QN ());
DFFSRX1 WX9784_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1917), .Q (WX9784), .QN ());
DFFSRX1 WX9788_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2158), .Q (WX9788), .QN ());
DFFSRX1 WX9792_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2121), .Q (WX9792), .QN ());
DFFSRX1 WX9796_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1805), .Q (WX9796), .QN ());
DFFSRX1 WX9800_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2209), .Q (WX9800), .QN ());
DFFSRX1 WX9808_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2313), .Q (WX9808), .QN ());
DFFSRX1 WX9810_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1766), .Q (WX9810), .QN ());
DFFSRX1 WX9814_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2321), .Q (WX9814), .QN ());
DFFSRX1 WX9822_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1982), .Q (WX9822), .QN ());
DFFSRX1 WX9830_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1897), .Q (WX9830), .QN ());
DFFSRX1 WX9838_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2261), .Q (WX9838), .QN ());
DFFSRX1 WX9842_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2199), .Q (WX9842), .QN ());
DFFSRX1 WX9846_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1727), .Q (WX9846), .QN ());
DFFSRX1 WX9850_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1480), .Q (WX9850), .QN ());
DFFSRX1 WX9854_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2125), .Q (WX9854), .QN ());
DFFSRX1 WX9856_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1868), .Q (WX9856), .QN ());
DFFSRX1 WX9858_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1488), .Q (WX9858), .QN ());
DFFSRX1 WX9862_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1712), .Q (WX9862), .QN ());
DFFSRX1 WX9864_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2238), .Q (WX9864), .QN ());
DFFSRX1 WX9866_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2386), .Q (WX9866), .QN ());
DFFSRX1 WX9870_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2504), .Q (WX9870), .QN ());
DFFSRX1 WX9874_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1733), .Q (WX9874), .QN ());
DFFSRX1 WX9880_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2213), .Q (WX9880), .QN ());
DFFSRX1 WX9882_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1740), .Q (WX9882), .QN ());
DFFSRX1 WX9884_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2287), .Q (WX9884), .QN ());
DFFSRX1 WX9888_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2385), .Q (WX9888), .QN ());
DFFSRX1 WX9890_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2003), .Q (WX9890), .QN ());
DFFSRX1 WX9892_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1859), .Q (WX9892), .QN ());
DFFSRX1 WX9896_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2222), .Q (WX9896), .QN ());
DFFSRX1 WX9898_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1887), .Q (WX9898), .QN ());
DFFSRX1 WX9900_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1971), .Q (WX9900), .QN ());
DFFSRX1 WX9908_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1768), .Q (WX9908), .QN ());
DFFSRX1 WX9910_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1782), .Q (WX9910), .QN ());
DFFSRX1 WX9914_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2377), .Q (WX9914), .QN ());
DFFSRX1 WX9918_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2014), .Q (WX9918), .QN ());
DFFSRX1 WX2140_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2135), .Q (WX2140), .QN ());
DFFSRX1 WX9930_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1945), .Q (WX9930), .QN ());
DFFSRX1 WX9932_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1846), .Q (WX9932), .QN ());
DFFSRX1 WX9934_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1968), .Q (WX9934), .QN ());
DFFSRX1 WX9938_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1484), .Q (WX9938), .QN ());
DFFSRX1 WX9942_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2380), .Q (WX9942), .QN ());
DFFSRX1 WX9946_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2340), .Q (WX9946), .QN ());
DFFSRX1 WX9948_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2021), .Q (WX9948), .QN ());
DFFSRX1 WX8587_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1810), .Q (WX8587), .QN ());
DFFSRX1 WX8609_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2033), .Q (WX8609), .QN ());
DFFSRX1 WX4680_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2019), .Q (WX4680), .QN ());
DFFSRX1 WX4610_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1949), .Q (WX4610), .QN ());
DFFSRX1 WX8599_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2009), .Q (WX8599), .QN ());
DFFSRX1 WX8595_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2056), .Q (WX8595), .QN ());
DFFSRX1 WX8583_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2236), .Q (WX8583), .QN ());
DFFSRX1 WX4590_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2126), .Q (WX4590), .QN ());
DFFSRX1 WX4594_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1826), .Q (WX4594), .QN ());
DFFSRX1 WX4602_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2162), .Q (WX4602), .QN ());
DFFSRX1 WX4604_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2273), .Q (WX4604), .QN ());
DFFSRX1 WX4608_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2293), .Q (WX4608), .QN ());
DFFSRX1 WX4618_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1841), .Q (WX4618), .QN ());
DFFSRX1 WX4614_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2338), .Q (WX4614), .QN ());
DFFSRX1 WX4622_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2310), .Q (WX4622), .QN ());
DFFSRX1 WX4624_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2292), .Q (WX4624), .QN ());
DFFSRX1 WX4628_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2165), .Q (WX4628), .QN ());
DFFSRX1 WX4632_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1716), .Q (WX4632), .QN ());
DFFSRX1 WX4642_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1806), .Q (WX4642), .QN ());
DFFSRX1 WX4644_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2122), .Q (WX4644), .QN ());
DFFSRX1 WX4648_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2185), .Q (WX4648), .QN ());
DFFSRX1 WX4656_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1566), .Q (WX4656), .QN ());
DFFSRX1 WX4660_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1942), .Q (WX4660), .QN ());
DFFSRX1 WX4668_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1966), .Q (WX4668), .QN ());
DFFSRX1 WX4672_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1879), .Q (WX4672), .QN ());
DFFSRX1 WX4676_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1995), .Q (WX4676), .QN ());
DFFSRX1 WX4678_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1770), .Q (WX4678), .QN ());
DFFSRX1 WX4684_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2058), .Q (WX4684), .QN ());
DFFSRX1 WX4686_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2032), .Q (WX4686), .QN ());
DFFSRX1 WX4688_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2001), .Q (WX4688), .QN ());
DFFSRX1 WX4692_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2153), .Q (WX4692), .QN ());
DFFSRX1 WX4694_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1836), .Q (WX4694), .QN ());
DFFSRX1 WX4696_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1799), .Q (WX4696), .QN ());
DFFSRX1 WX8607_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2024), .Q (WX8607), .QN ());
DFFSRX1 WX4704_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1943), .Q (WX4704), .QN ());
DFFSRX1 WX4714_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2025), .Q (WX4714), .QN ());
DFFSRX1 WX4720_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2005), .Q (WX4720), .QN ());
DFFSRX1 WX4722_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1778), .Q (WX4722), .QN ());
DFFSRX1 WX4724_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2063), .Q (WX4724), .QN ());
DFFSRX1 WX4728_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2065), .Q (WX4728), .QN ());
DFFSRX1 WX4730_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2072), .Q (WX4730), .QN ());
DFFSRX1 WX4732_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1771), .Q (WX4732), .QN ());
DFFSRX1 WX4736_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1769), .Q (WX4736), .QN ());
DFFSRX1 WX4738_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2069), .Q (WX4738), .QN ());
DFFSRX1 WX4740_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2217), .Q (WX4740), .QN ());
DFFSRX1 WX4744_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2079), .Q (WX4744), .QN ());
DFFSRX1 WX4748_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1929), .Q (WX4748), .QN ());
DFFSRX1 WX4752_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2115), .Q (WX4752), .QN ());
DFFSRX1 WX4756_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1759), .Q (WX4756), .QN ());
DFFSRX1 WX2188_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1869), .Q (WX2188), .QN ());
DFFSRX1 WX4760_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2078), .Q (WX4760), .QN ());
DFFSRX1 WX4764_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1760), .Q (WX4764), .QN ());
DFFSRX1 WX4768_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2108), .Q (WX4768), .QN ());
DFFSRX1 WX4770_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1821), .Q (WX4770), .QN ());
DFFSRX1 WX4772_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1751), .Q (WX4772), .QN ());
DFFSRX1 WX4776_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2105), .Q (WX4776), .QN ());
DFFSRX1 WX4778_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1844), .Q (WX4778), .QN ());
DFFSRX1 WX7362_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1941), .Q (WX7362), .QN ());
DFFSRX1 WX4698_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2204), .Q (WX4698), .QN ());
DFFSRX1 WX9950_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1927), .Q (WX9950), .QN ());
DFFSRX1 WX4650_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2006), .Q (WX4650), .QN ());
DFFSRX1 WX4664_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2028), .Q (WX4664), .QN ());
DFFSRX1 WX9818_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2230), .Q (WX9818), .QN ());
DFFSRX1 WX11137_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2382), .Q (WX11137), .QN ());
DFFSRX1 WX8533_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1802), .Q (WX8533), .QN ());
DFFSRX1 WX5881_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1477), .Q (WX5881), .QN ());
DFFSRX1 WX5883_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2291), .Q (WX5883), .QN ());
DFFSRX1 WX5887_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2515), .Q (WX5887), .QN ());
DFFSRX1 WX5889_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1777), .Q (WX5889), .QN ());
DFFSRX1 WX5891_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1786), .Q (WX5891), .QN ());
DFFSRX1 WX5895_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2235), .Q (WX5895), .QN ());
DFFSRX1 WX5897_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1795), .Q (WX5897), .QN ());
DFFSRX1 WX8529_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1827), .Q (WX8529), .QN ());
DFFSRX1 WX5901_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1476), .Q (WX5901), .QN ());
DFFSRX1 WX5905_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1798), .Q (WX5905), .QN ());
DFFSRX1 WX5909_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1728), .Q (WX5909), .QN ());
DFFSRX1 WX5911_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1803), .Q (WX5911), .QN ());
DFFSRX1 WX5913_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2047), .Q (WX5913), .QN ());
DFFSRX1 WX5917_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1882), .Q (WX5917), .QN ());
DFFSRX1 WX5919_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2017), .Q (WX5919), .QN ());
DFFSRX1 WX5921_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1789), .Q (WX5921), .QN ());
DFFSRX1 WX5925_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2150), .Q (WX5925), .QN ());
DFFSRX1 WX5929_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1809), .Q (WX5929), .QN ());
DFFSRX1 WX5933_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1747), .Q (WX5933), .QN ());
DFFSRX1 WX5935_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2315), .Q (WX5935), .QN ());
DFFSRX1 WX5937_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1702), .Q (WX5937), .QN ());
DFFSRX1 WX5915_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2330), .Q (WX5915), .QN ());
DFFSRX1 WX5941_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1963), .Q (WX5941), .QN ());
DFFSRX1 WX5943_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2271), .Q (WX5943), .QN ());
DFFSRX1 WX5945_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1937), .Q (WX5945), .QN ());
DFFSRX1 WX5949_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1808), .Q (WX5949), .QN ());
DFFSRX1 WX5951_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1834), .Q (WX5951), .QN ());
DFFSRX1 WX5953_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1881), .Q (WX5953), .QN ());
DFFSRX1 WX5957_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1781), .Q (WX5957), .QN ());
DFFSRX1 WX5959_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1835), .Q (WX5959), .QN ());
DFFSRX1 WX5961_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1831), .Q (WX5961), .QN ());
DFFSRX1 WX5965_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2420), .Q (WX5965), .QN ());
DFFSRX1 WX5967_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1953), .Q (WX5967), .QN ());
DFFSRX1 WX5969_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1854), .Q (WX5969), .QN ());
DFFSRX1 WX5973_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1763), .Q (WX5973), .QN ());
DFFSRX1 WX5975_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1858), .Q (WX5975), .QN ());
DFFSRX1 WX5977_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1855), .Q (WX5977), .QN ());
DFFSRX1 WX5981_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1862), .Q (WX5981), .QN ());
DFFSRX1 WX5983_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2365), .Q (WX5983), .QN ());
DFFSRX1 WX5985_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1701), .Q (WX5985), .QN ());
DFFSRX1 WX5989_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2358), .Q (WX5989), .QN ());
DFFSRX1 WX8521_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2018), .Q (WX8521), .QN ());
DFFSRX1 WX5991_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2335), .Q (WX5991), .QN ());
DFFSRX1 WX5995_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1871), .Q (WX5995), .QN ());
DFFSRX1 WX5999_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1874), .Q (WX5999), .QN ());
DFFSRX1 WX6003_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2317), .Q (WX6003), .QN ());
DFFSRX1 WX6005_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2534), .Q (WX6005), .QN ());
DFFSRX1 WX6007_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1892), .Q (WX6007), .QN ());
DFFSRX1 WX6011_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2189), .Q (WX6011), .QN ());
DFFSRX1 WX6013_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2192), .Q (WX6013), .QN ());
DFFSRX1 WX6015_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2050), .Q (WX6015), .QN ());
DFFSRX1 WX6019_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1811), .Q (WX6019), .QN ());
DFFSRX1 WX6023_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2161), .Q (WX6023), .QN ());
DFFSRX1 WX6027_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1910), .Q (WX6027), .QN ());
DFFSRX1 WX6029_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2157), .Q (WX6029), .QN ());
DFFSRX1 WX6031_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1915), .Q (WX6031), .QN ());
DFFSRX1 WX6035_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1916), .Q (WX6035), .QN ());
DFFSRX1 WX6039_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1923), .Q (WX6039), .QN ());
DFFSRX1 WX6043_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2286), .Q (WX6043), .QN ());
DFFSRX1 WX6045_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2007), .Q (WX6045), .QN ());
DFFSRX1 WX6047_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1932), .Q (WX6047), .QN ());
DFFSRX1 WX6055_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2269), .Q (WX6055), .QN ());
DFFSRX1 WX6059_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1794), .Q (WX6059), .QN ());
DFFSRX1 WX6063_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2254), .Q (WX6063), .QN ());
DFFSRX1 WX6067_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1979), .Q (WX6067), .QN ());
DFFSRX1 WX6069_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1812), .Q (WX6069), .QN ());
DFFSRX1 WX6071_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1752), .Q (WX6071), .QN ());
DFFSRX1 WX4718_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1934), .Q (WX4718), .QN ());
DFFSRX1 WX8507_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1758), .Q (WX8507), .QN ());
DFFSRX1 WX9812_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1852), .Q (WX9812), .QN ());
DFFSRX1 WX2068_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2476), .Q (WX2068), .QN ());
DFFSRX1 WX2072_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2087), .Q (WX2072), .QN ());
DFFSRX1 WX2076_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2081), .Q (WX2076), .QN ());
DFFSRX1 WX2080_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2044), .Q (WX2080), .QN ());
DFFSRX1 WX2084_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1753), .Q (WX2084), .QN ());
DFFSRX1 WX2088_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1832), .Q (WX2088), .QN ());
DFFSRX1 WX4616_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1926), .Q (WX4616), .QN ());
DFFSRX1 WX2090_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1739), .Q (WX2090), .QN ());
DFFSRX1 WX2096_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1757), .Q (WX2096), .QN ());
DFFSRX1 WX2094_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1743), .Q (WX2094), .QN ());
DFFSRX1 WX2102_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1939), .Q (WX2102), .QN ());
DFFSRX1 WX2104_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1857), .Q (WX2104), .QN ());
DFFSRX1 WX2106_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2301), .Q (WX2106), .QN ());
DFFSRX1 WX2110_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1749), .Q (WX2110), .QN ());
DFFSRX1 WX2112_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2029), .Q (WX2112), .QN ());
DFFSRX1 WX2114_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1779), .Q (WX2114), .QN ());
DFFSRX1 _2276__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1497), .Q (_2276_), .QN ());
DFFSRX1 WX2118_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1748), .Q (WX2118), .QN ());
DFFSRX1 WX2120_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2268), .Q (WX2120), .QN ());
DFFSRX1 WX2122_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1851), .Q (WX2122), .QN ());
DFFSRX1 WX2126_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1983), .Q (WX2126), .QN ());
DFFSRX1 WX2128_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2336), .Q (WX2128), .QN ());
DFFSRX1 WX2132_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2368), .Q (WX2132), .QN ());
DFFSRX1 WX2136_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1479), .Q (WX2136), .QN ());
DFFSRX1 WX2142_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1940), .Q (WX2142), .QN ());
DFFSRX1 WX2144_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1744), .Q (WX2144), .QN ());
DFFSRX1 WX2148_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2259), .Q (WX2148), .QN ());
DFFSRX1 WX2152_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2239), .Q (WX2152), .QN ());
DFFSRX1 WX2154_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1843), .Q (WX2154), .QN ());
DFFSRX1 WX2158_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2030), .Q (WX2158), .QN ());
DFFSRX1 WX2160_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2040), .Q (WX2160), .QN ());
DFFSRX1 WX2162_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2049), .Q (WX2162), .QN ());
DFFSRX1 WX2164_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2052), .Q (WX2164), .QN ());
DFFSRX1 WX2168_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2100), .Q (WX2168), .QN ());
DFFSRX1 WX2170_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2075), .Q (WX2170), .QN ());
DFFSRX1 WX2172_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2089), .Q (WX2172), .QN ());
DFFSRX1 WX2176_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2232), .Q (WX2176), .QN ());
DFFSRX1 WX2178_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2186), .Q (WX2178), .QN ());
DFFSRX1 WX2180_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1823), .Q (WX2180), .QN ());
DFFSRX1 WX9912_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1486), .Q (WX9912), .QN ());
DFFSRX1 WX2186_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2225), .Q (WX2186), .QN ());
DFFSRX1 WX2190_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2245), .Q (WX2190), .QN ());
DFFSRX1 WX11095_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1722), .Q (WX11095), .QN ());
DFFSRX1 WX8481_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1845), .Q (WX8481), .QN ());
DFFSRX1 WX11055_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1866), .Q (WX11055), .QN ());
DFFSRX1 WX11057_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1707), .Q (WX11057), .QN ());
DFFSRX1 WX11061_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2023), .Q (WX11061), .QN ());
DFFSRX1 WX11059_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2091), .Q (WX11059), .QN ());
DFFSRX1 WX11065_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2060), .Q (WX11065), .QN ());
DFFSRX1 WX11067_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1938), .Q (WX11067), .QN ());
DFFSRX1 WX11069_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2441), .Q (WX11069), .QN ());
DFFSRX1 WX11073_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1872), .Q (WX11073), .QN ());
DFFSRX1 WX11075_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2219), .Q (WX11075), .QN ());
DFFSRX1 WX11077_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1819), .Q (WX11077), .QN ());
DFFSRX1 WX11081_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2051), .Q (WX11081), .QN ());
DFFSRX1 WX11085_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1800), .Q (WX11085), .QN ());
DFFSRX1 WX11089_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2187), .Q (WX11089), .QN ());
DFFSRX1 WX11093_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2106), .Q (WX11093), .QN ());
DFFSRX1 WX11097_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2401), .Q (WX11097), .QN ());
DFFSRX1 WX11099_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1715), .Q (WX11099), .QN ());
DFFSRX1 WX11103_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1711), .Q (WX11103), .QN ());
DFFSRX1 WX9554_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1526), .Q (), .QN (WX9554));
DFFSRX1 WX4390_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1987), .Q (), .QN (WX4390));
DFFSRX1 WX3455_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2092), .Q (WX3455), .QN ());
DFFSRX1 WX4598_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1950), .Q (WX4598), .QN ());
DFFSRX1 WX11083_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1796), .Q (WX11083), .QN ());
DFFSRX1 WX11087_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1756), .Q (WX11087), .QN ());
DFFSRX1 WX7350_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1902), .Q (WX7350), .QN ());
DFFSRX1 WX11091_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2146), .Q (WX11091), .QN ());
DFFSRX1 _2166__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1628), .Q (_2166_), .QN ());
DFFSRX1 WX4712_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1478), .Q (WX4712), .QN ());
DFFSRX1 _2168__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1626), .Q (_2168_), .QN ());
DFFSRX1 _2204__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1600), .Q (_2204_), .QN ());
DFFSRX1 WX8485_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1842), .Q (WX8485), .QN ());
BUFX3 g63216(.A (n_2894), .Y (n_4058));
CLKBUFX3 g63214(.A (n_2894), .Y (n_3168));
DFFSRX1 WX9886_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2334), .Q (WX9886), .QN ());
DFFSRX1 _2315__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1548), .Q (_2315_), .QN ());
DFFSRX1 WX4742_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2099), .Q (WX4742), .QN ());
INVX4 g63152(.A (n_2897), .Y (n_5242));
DFFSRX1 WX5681_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2144), .Q (), .QN (WX5681));
INVX2 g63175(.A (n_6437), .Y (n_4670));
BUFX3 g63192(.A (n_6452), .Y (n_4017));
INVX2 g63190(.A (n_6452), .Y (n_3169));
BUFX3 g63191(.A (n_6452), .Y (n_4095));
DFFSRX1 WX11141_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2076), .Q (WX11141), .QN ());
BUFX3 g63186(.A (n_6452), .Y (n_4103));
DFFSRX1 WX9844_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1700), .Q (WX9844), .QN ());
DFFSRX1 _2318__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1546), .Q (_2318_), .QN ());
BUFX3 g63185(.A (n_6452), .Y (n_4104));
DFFSRX1 _2206__reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1570), .Q (_2206_), .QN ());
DFFSRX1 WX7356_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1994), .Q (WX7356), .QN ());
DFFSRX1 WX9922_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1888), .Q (WX9922), .QN ());
INVX2 g63154(.A (n_2897), .Y (n_5709));
DFFSRX1 WX9878_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1780), .Q (WX9878), .QN ());
DFFSRX1 WX4774_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2082), .Q (WX4774), .QN ());
DFFSRX1 WX7208_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_2210), .Q (WX7208), .QN ());
DFFSRX1 WX4766_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1884), .Q (WX4766), .QN ());
INVX1 g63156(.A (n_2897), .Y (n_5843));
DFFSRX1 WX2040_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1287), .Q (WX2040), .QN ());
DFFSRX1 WX5657_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1464), .Q (WX5657), .QN ());
DFFSRX1 WX877_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1280), .Q (WX877), .QN ());
DFFSRX1 WX887_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1448), .Q (WX887), .QN ());
DFFSRX1 WX711_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1326), .Q (WX711), .QN ());
DFFSRX1 WX857_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1366), .Q (WX857), .QN ());
INVX8 g63078(.A (n_2840), .Y (n_4562));
DFFSRX1 WX799_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1407), .Q (WX799), .QN ());
DFFSRX1 WX743_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1330), .Q (WX743), .QN ());
INVX1 g63071(.A (n_2840), .Y (n_3158));
DFFSRX1 WX6950_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1459), .Q (WX6950), .QN ());
MX2X1 g60709(.A (n_2838), .B (n_2837), .S0 (WX8457), .Y (n_2839));
MX2X1 g60712(.A (n_2813), .B (n_2953), .S0 (WX8459), .Y (n_2836));
DFFSRX1 WX875_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1353), .Q (WX875), .QN ());
MX2X1 g60741(.A (n_2813), .B (n_2817), .S0 (WX4558), .Y (n_2835));
MX2X1 g60744(.A (n_2935), .B (n_2770), .S0 (WX3263), .Y (n_2833));
MX2X1 g60747(.A (n_3140), .B (n_2826), .S0 (WX9696), .Y (n_2831));
DFFSRX1 WX713_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1382), .Q (WX713), .QN ());
BUFX3 g63052(.A (n_2840), .Y (n_4100));
MX2X1 g60754(.A (n_2829), .B (n_2828), .S0 (WX4562), .Y (n_2830));
MX2X1 g60757(.A (n_2826), .B (n_860), .S0 (n_2825), .Y (n_2827));
BUFX3 g63050(.A (n_2840), .Y (n_4094));
MX2X1 g60765(.A (n_2838), .B (n_3089), .S0 (WX4564), .Y (n_2824));
MX2X1 g60766(.A (n_3137), .B (n_2800), .S0 (WX9704), .Y (n_2823));
MX2X1 g60770(.A (n_2776), .B (n_2770), .S0 (WX5855), .Y (n_2822));
MX2X1 g60773(.A (n_2809), .B (n_3089), .S0 (WX4566), .Y (n_2820));
MX2X1 g60781(.A (n_2776), .B (n_2817), .S0 (WX4568), .Y (n_2818));
MX2X1 g60784(.A (n_2815), .B (n_2828), .S0 (WX4570), .Y (n_2816));
MX2X1 g60787(.A (n_2813), .B (n_2770), .S0 (WX4572), .Y (n_2814));
MX2X1 g60797(.A (n_3140), .B (n_2826), .S0 (WX9724), .Y (n_2812));
MX2X1 g60800(.A (n_6422), .B (n_3140), .S0 (n_1337), .Y (n_2811));
MX2X1 g60803(.A (n_2809), .B (n_2775), .S0 (WX4576), .Y (n_2810));
MX2X1 g60813(.A (n_2826), .B (n_860), .S0 (n_1335), .Y (n_2807));
MX2X1 g60822(.A (n_2935), .B (n_3089), .S0 (WX9740), .Y (n_2806));
MX2X1 g60827(.A (n_2716), .B (n_2795), .S0 (WX9742), .Y (n_2805));
MX2X1 g60832(.A (n_6422), .B (n_860), .S0 (n_1359), .Y (n_2803));
MX2X1 g60833(.A (n_3120), .B (n_2800), .S0 (WX10991), .Y (n_2801));
MX2X1 g60834(.A (n_2798), .B (n_2795), .S0 (WX5853), .Y (n_2799));
MX2X1 g60835(.A (n_2935), .B (n_2795), .S0 (WX9746), .Y (n_2797));
MX2X1 g60837(.A (n_3120), .B (n_2800), .S0 (WX3235), .Y (n_2794));
MX2X1 g60840(.A (n_2798), .B (n_2770), .S0 (WX9748), .Y (n_2793));
DFFSRX1 WX8243_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1454), .Q (WX8243), .QN ());
MX2X1 g60853(.A (n_2813), .B (n_2837), .S0 (WX9754), .Y (n_2792));
MX2X1 g60880(.A (n_6422), .B (n_860), .S0 (n_1357), .Y (n_2791));
MX2X1 g60888(.A (n_2815), .B (n_6512), .S0 (WX5871), .Y (n_2790));
MX2X1 g60899(.A (n_2826), .B (n_6432), .S0 (n_1284), .Y (n_2789));
MX2X1 g60905(.A (n_2744), .B (n_2757), .S0 (n_1431), .Y (n_2788));
MX2X1 g60907(.A (n_2826), .B (n_858), .S0 (n_1341), .Y (n_2787));
MX2X1 g60909(.A (n_2826), .B (n_3140), .S0 (n_1412), .Y (n_2786));
DFFSRX1 WX753_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1389), .Q (WX753), .QN ());
MX2X1 g60920(.A (n_3027), .B (n_2826), .S0 (WX5839), .Y (n_2784));
MX2X1 g60926(.A (n_3021), .B (n_2826), .S0 (WX3249), .Y (n_2783));
DFFSRX1 WX733_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1404), .Q (WX733), .QN ());
MX2X1 g60938(.A (n_2744), .B (n_2757), .S0 (n_1350), .Y (n_2782));
MX2X1 g60944(.A (n_2829), .B (n_2953), .S0 (WX5859), .Y (n_2780));
MX2X1 g60945(.A (n_2826), .B (n_858), .S0 (n_1345), .Y (n_2778));
MX2X1 g60957(.A (n_2776), .B (n_2775), .S0 (WX5869), .Y (n_2777));
DFFSRX1 WX751_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1418), .Q (WX751), .QN ());
MX2X1 g60966(.A (n_2826), .B (n_858), .S0 (n_1427), .Y (n_2774));
MX2X1 g60970(.A (n_2826), .B (n_6432), .S0 (n_1419), .Y (n_2773));
MX2X1 g60971(.A (n_2744), .B (n_2757), .S0 (n_1451), .Y (n_2772));
MX2X1 g60975(.A (n_2776), .B (n_2770), .S0 (WX5867), .Y (n_2771));
MX2X1 g60978(.A (n_2776), .B (n_2795), .S0 (WX5851), .Y (n_2769));
MX2X1 g60981(.A (n_2826), .B (n_858), .S0 (n_1323), .Y (n_2768));
MX2X1 g60995(.A (n_2744), .B (n_2757), .S0 (n_1348), .Y (n_2767));
MX2X1 g60996(.A (n_2838), .B (n_2817), .S0 (WX5873), .Y (n_2765));
DFFSRX1 WX2060_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1319), .Q (WX2060), .QN ());
MX2X1 g61001(.A (n_6423), .B (n_2800), .S0 (WX3251), .Y (n_2763));
MX2X1 g61002(.A (n_6423), .B (n_2800), .S0 (WX11017), .Y (n_2762));
MX2X1 g61013(.A (n_2813), .B (n_2837), .S0 (WX3269), .Y (n_2761));
MX2X1 g61021(.A (n_2716), .B (n_2988), .S0 (WX8455), .Y (n_2760));
MX2X1 g61022(.A (n_2744), .B (n_2757), .S0 (n_1286), .Y (n_2759));
MX2X1 g61032(.A (n_2829), .B (n_2755), .S0 (WX3271), .Y (n_2756));
MX2X1 g61040(.A (n_2744), .B (n_2757), .S0 (n_1374), .Y (n_2754));
MX2X1 g61044(.A (n_2815), .B (n_3089), .S0 (WX11021), .Y (n_2752));
MX2X1 g61048(.A (n_2744), .B (n_2757), .S0 (n_1288), .Y (n_2750));
DFFSRX1 WX2008_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1340), .Q (WX2008), .QN ());
MX2X1 g61051(.A (n_2809), .B (n_2988), .S0 (WX9744), .Y (n_2749));
MX2X1 g61056(.A (n_2809), .B (n_2817), .S0 (WX8453), .Y (n_2746));
DFFSRX1 WX9536_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1453), .Q (WX9536), .QN ());
MX2X1 g61080(.A (n_2744), .B (n_2757), .S0 (n_1309), .Y (n_2745));
MX2X1 g61088(.A (n_2744), .B (n_2757), .S0 (n_1282), .Y (n_2743));
MX2X1 g61095(.A (n_2986), .B (n_2953), .S0 (WX11025), .Y (n_2742));
MX2X1 g61097(.A (n_2986), .B (n_6512), .S0 (WX3277), .Y (n_2741));
MX2X1 g61103(.A (n_2776), .B (n_6512), .S0 (WX8451), .Y (n_2739));
MX2X1 g61106(.A (n_6513), .B (n_2770), .S0 (WX3279), .Y (n_2738));
MX2X1 g61113(.A (n_2744), .B (n_2757), .S0 (n_2691), .Y (n_2737));
MX2X1 g61115(.A (n_2813), .B (n_2953), .S0 (WX11027), .Y (n_2736));
MX2X1 g61121(.A (n_2829), .B (n_2953), .S0 (WX8447), .Y (n_2734));
MX2X1 g61122(.A (n_2744), .B (n_2757), .S0 (n_1442), .Y (n_2733));
MX2X1 g61123(.A (n_2798), .B (n_2837), .S0 (WX7154), .Y (n_2732));
MX2X1 g61133(.A (n_2744), .B (n_2757), .S0 (n_1328), .Y (n_2731));
MX2X1 g61134(.A (n_2815), .B (n_2988), .S0 (WX7160), .Y (n_2730));
MX2X1 g61142(.A (n_2935), .B (n_2775), .S0 (WX3283), .Y (n_2729));
MX2X1 g61144(.A (n_2716), .B (n_2817), .S0 (WX7164), .Y (n_2728));
MX2X1 g61146(.A (n_6422), .B (n_860), .S0 (n_1339), .Y (n_2726));
MX2X1 g61154(.A (n_2809), .B (n_2755), .S0 (WX7168), .Y (n_2725));
MX2X1 g61160(.A (n_2744), .B (n_2757), .S0 (n_1437), .Y (n_2724));
MX2X1 g61161(.A (n_2798), .B (n_2775), .S0 (WX7170), .Y (n_2722));
MX2X1 g61170(.A (n_2744), .B (n_2757), .S0 (n_1429), .Y (n_2721));
MX2X1 g61173(.A (n_2815), .B (n_2988), .S0 (WX3287), .Y (n_2720));
DFFSRX1 WX833_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1447), .Q (WX833), .QN ());
MX2X1 g61177(.A (n_2716), .B (n_2770), .S0 (WX3289), .Y (n_2719));
MX2X1 g61178(.A (n_2744), .B (n_2757), .S0 (n_1318), .Y (n_2718));
DFFSRX1 WX2024_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1321), .Q (WX2024), .QN ());
MX2X1 g61184(.A (n_2716), .B (n_2775), .S0 (WX3291), .Y (n_2717));
MX2X1 g61192(.A (n_2744), .B (n_2757), .S0 (n_2675), .Y (n_2715));
DFFSRX1 WX2044_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1289), .Q (WX2044), .QN ());
MX2X1 g61200(.A (n_2826), .B (n_3140), .S0 (n_1449), .Y (n_2714));
MX2X1 g61201(.A (n_2815), .B (n_2795), .S0 (WX11041), .Y (n_2713));
MX2X1 g61202(.A (n_2798), .B (n_2837), .S0 (WX8443), .Y (n_2712));
MX2X1 g61206(.A (n_2815), .B (n_2817), .S0 (WX4580), .Y (n_2711));
MX2X1 g61208(.A (n_2813), .B (n_2988), .S0 (WX11043), .Y (n_2710));
MX2X1 g61213(.A (n_3137), .B (n_2826), .S0 (WX3233), .Y (n_2709));
MX2X1 g61227(.A (n_2809), .B (n_2828), .S0 (WX9738), .Y (n_2708));
MX2X1 g61230(.A (n_3021), .B (n_2826), .S0 (WX8415), .Y (n_2707));
MX2X1 g61234(.A (n_3137), .B (n_2826), .S0 (WX8417), .Y (n_2706));
MX2X1 g61237(.A (n_2716), .B (n_2795), .S0 (WX11047), .Y (n_2705));
MX2X1 g61239(.A (n_3137), .B (n_2826), .S0 (WX8419), .Y (n_2704));
DFFSRX1 WX803_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1388), .Q (WX803), .QN ());
MX2X1 g61246(.A (n_2826), .B (n_3140), .S0 (n_1320), .Y (n_2703));
MX2X1 g61249(.A (n_3140), .B (n_2800), .S0 (WX4524), .Y (n_2702));
MX2X1 g61258(.A (n_2716), .B (n_2775), .S0 (WX11049), .Y (n_2701));
MX2X1 g61265(.A (n_2826), .B (n_6432), .S0 (n_1421), .Y (n_2700));
DFFSRX1 WX2062_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1452), .Q (WX2062), .QN ());
DFFSRX1 WX719_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1365), .Q (WX719), .QN ());
MX2X1 g61274(.A (n_2809), .B (n_2755), .S0 (WX9734), .Y (n_2699));
MX2X1 g61276(.A (n_2829), .B (n_2755), .S0 (WX11051), .Y (n_2698));
MX2X1 g61279(.A (n_2935), .B (n_2817), .S0 (WX8435), .Y (n_2697));
MX2X1 g61288(.A (n_2716), .B (n_2755), .S0 (WX8439), .Y (n_2696));
MX2X1 g61300(.A (n_3137), .B (n_2800), .S0 (WX3257), .Y (n_2695));
MX2X1 g61304(.A (n_2935), .B (n_2953), .S0 (WX9758), .Y (n_2694));
DFFSRX1 WX723_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1423), .Q (WX723), .QN ());
DFFSRX1 WX889_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1380), .Q (WX889), .QN ());
BUFX3 g61384(.A (n_7089), .Y (n_2926));
BUFX3 g61393(.A (n_7089), .Y (n_2925));
BUFX3 g61402(.A (n_7089), .Y (n_2924));
BUFX3 g61420(.A (n_7089), .Y (n_2922));
BUFX3 g61429(.A (n_7089), .Y (n_2921));
BUFX3 g61456(.A (n_7089), .Y (n_2920));
DFFSRX1 WX2028_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1324), .Q (WX2028), .QN ());
NOR2X1 g61542(.A (n_2691), .B (n_3188), .Y (n_2692));
DFFSRX1 WX871_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1435), .Q (WX871), .QN ());
AND2X1 g61572(.A (WX11175), .B (n_2298), .Y (n_2690));
AND2X1 g61573(.A (WX11089), .B (n_2298), .Y (n_2689));
AND2X1 g61577(.A (WX9770), .B (n_2298), .Y (n_2687));
DFFSRX1 WX865_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1399), .Q (WX865), .QN ());
AND2X1 g61638(.A (WX11135), .B (n_2298), .Y (n_2686));
DFFSRX1 WX897_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1362), .Q (WX897), .QN ());
AND2X1 g61647(.A (WX4556), .B (n_2298), .Y (n_2685));
AND2X1 g61648(.A (WX11143), .B (n_2298), .Y (n_2684));
DFFSRX1 WX793_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1400), .Q (WX793), .QN ());
AND2X1 g61675(.A (WX4542), .B (n_2298), .Y (n_2682));
AND2X1 g61676(.A (WX9808), .B (n_2298), .Y (n_2681));
AND2X1 g61716(.A (WX11105), .B (n_2298), .Y (n_2680));
AND2X1 g58600(.A (WX11117), .B (n_2298), .Y (n_2678));
DFFSRX1 WX869_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1398), .Q (WX869), .QN ());
AND2X1 g61801(.A (WX7152), .B (n_2298), .Y (n_2677));
NOR2X1 g61817(.A (n_2675), .B (n_3188), .Y (n_2676));
DFFSRX1 WX2002_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1338), .Q (WX2002), .QN ());
DFFSRX1 WX2020_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1422), .Q (WX2020), .QN ());
DFFSRX1 WX3071_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1279), .Q (WX3071), .QN ());
AND2X1 g61914(.A (WX9862), .B (n_2378), .Y (n_2673));
AND2X1 g61934(.A (WX9764), .B (n_2378), .Y (n_2671));
AND2X1 g61960(.A (WX4682), .B (n_2298), .Y (n_2670));
AND2X1 g61964(.A (WX4690), .B (n_2378), .Y (n_2669));
AND2X1 g62074(.A (WX3375), .B (n_2298), .Y (n_2668));
AND2X1 g62097(.A (WX3369), .B (n_2298), .Y (n_2667));
AND2X1 g62137(.A (WX3305), .B (n_2298), .Y (n_2666));
DFFSRX1 WX2054_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1329), .Q (WX2054), .QN ());
DFFSRX1 WX2056_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1438), .Q (WX2056), .QN ());
AND2X1 g62215(.A (WX4610), .B (n_2378), .Y (n_2665));
AND2X1 g62219(.A (WX5987), .B (n_2378), .Y (n_2664));
AND2X1 g62221(.A (WX11051), .B (n_2378), .Y (n_2663));
DFFSRX1 WX853_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1327), .Q (WX853), .QN ());
DFFSRX1 WX2036_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1432), .Q (WX2036), .QN ());
DFFSRX1 WX849_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1333), .Q (WX849), .QN ());
XOR2X1 g58894(.A (_2119_), .B (n_1221), .Y (n_2662));
XOR2X1 g58895(.A (_2183_), .B (n_1044), .Y (n_2661));
AND2X1 g62490(.A (WX8585), .B (n_2298), .Y (n_2660));
AND2X1 g62491(.A (WX8587), .B (n_2298), .Y (n_2659));
XOR2X1 g58896(.A (_2112_), .B (n_1254), .Y (n_2658));
XOR2X1 g58897(.A (_2284_), .B (n_1111), .Y (n_2657));
XOR2X1 g58900(.A (_2124_), .B (n_1231), .Y (n_2656));
XOR2X1 g58901(.A (_2144_), .B (n_1047), .Y (n_2655));
XOR2X1 g58902(.A (_2151_), .B (n_1186), .Y (n_2654));
XOR2X1 g58903(.A (_2156_), .B (n_1181), .Y (n_2653));
XOR2X1 g58904(.A (_2176_), .B (n_1210), .Y (n_2652));
XOR2X1 g58905(.A (_2188_), .B (n_1257), .Y (n_2651));
AND2X1 g62520(.A (WX11171), .B (n_2298), .Y (n_2650));
XOR2X1 g58906(.A (_2208_), .B (n_1154), .Y (n_2649));
XOR2X1 g58907(.A (_2247_), .B (n_1237), .Y (n_2648));
XOR2X1 g58908(.A (_2215_), .B (n_1150), .Y (n_2647));
XOR2X1 g58909(.A (_2220_), .B (n_1148), .Y (n_2646));
AND2X1 g62532(.A (WX3337), .B (n_2298), .Y (n_2645));
XOR2X1 g58910(.A (_2240_), .B (n_1135), .Y (n_2644));
XOR2X1 g58911(.A (_2252_), .B (n_1116), .Y (n_2643));
XOR2X1 g58912(.A (_2272_), .B (n_1120), .Y (n_2642));
XOR2X1 g58913(.A (_2279_), .B (n_1114), .Y (n_2641));
XOR2X1 g58914(.A (_2311_), .B (n_1094), .Y (n_2640));
XOR2X1 g58915(.A (_2336_), .B (n_1082), .Y (n_2639));
AND2X1 g62550(.A (WX5863), .B (n_2298), .Y (n_2638));
XOR2X1 g58916(.A (_2343_), .B (n_1079), .Y (n_2637));
XOR2X1 g58917(.A (_2348_), .B (n_1076), .Y (n_2636));
XOR2X1 g58918(.A (_2304_), .B (n_1051), .Y (n_2635));
XOR2X1 g58919(.A (_2316_), .B (n_1091), .Y (n_2634));
DFFSRX1 WX829_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1314), .Q (WX829), .QN ());
AND2X1 g62615(.A (WX2034), .B (n_2298), .Y (n_2633));
AND2X1 g62680(.A (WX2082), .B (n_2298), .Y (n_2632));
DFFSRX1 WX827_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1458), .Q (WX827), .QN ());
DFFSRX1 WX2030_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1428), .Q (WX2030), .QN ());
DFFSRX1 WX747_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1373), .Q (WX747), .QN ());
DFFSRX1 WX2016_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1342), .Q (WX2016), .QN ());
DFFSRX1 WX861_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1347), .Q (WX861), .QN ());
DFFSRX1 WX795_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1415), .Q (WX795), .QN ());
DFFSRX1 WX735_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1332), .Q (WX735), .QN ());
DFFSRX1 WX883_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1410), .Q (WX883), .QN ());
DFFSRX1 WX787_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1378), .Q (WX787), .QN ());
DFFSRX1 WX825_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1411), .Q (WX825), .QN ());
CLKBUFX1 g63148(.A (n_6437), .Y (n_3162));
DFFSRX1 WX839_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1354), .Q (WX839), .QN ());
DFFSRX1 WX821_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1436), .Q (WX821), .QN ());
DFFSRX1 WX757_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1409), .Q (WX757), .QN ());
NOR2X1 g57541(.A (n_848), .B (n_3188), .Y (n_2631));
BUFX3 g63051(.A (n_2840), .Y (n_4101));
BUFX3 g63053(.A (n_2840), .Y (n_4106));
DFFSRX1 WX731_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1433), .Q (WX731), .QN ());
DFFSRX1 WX783_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1444), .Q (WX783), .QN ());
AND2X1 g62721(.A (WX7208), .B (n_2298), .Y (n_2630));
NOR2X1 g59242(.A (n_1195), .B (n_3188), .Y (n_2629));
NOR2X1 g59244(.A (n_1104), .B (n_2620), .Y (n_2628));
DFFSRX1 WX737_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1364), .Q (WX737), .QN ());
NOR2X1 g59248(.A (n_1097), .B (n_3188), .Y (n_2627));
NOR2X1 g59249(.A (n_1065), .B (n_3690), .Y (n_2626));
NOR2X1 g59250(.A (n_1131), .B (n_3690), .Y (n_2625));
NOR2X1 g59251(.A (n_1245), .B (n_2851), .Y (n_2624));
NOR2X1 g59257(.A (n_1233), .B (n_3690), .Y (n_2622));
NOR2X1 g59266(.A (n_1205), .B (n_2620), .Y (n_2621));
DFFSRX1 WX487_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1456), .Q (WX487), .QN ());
DFFSRX1 WX855_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1465), .Q (WX855), .QN ());
DFFSRX1 WX717_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1393), .Q (WX717), .QN ());
DFFSRX1 WX837_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1424), .Q (WX837), .QN ());
NOR2X1 g59294(.A (n_1023), .B (n_3188), .Y (n_2619));
DFFSRX1 WX823_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1377), .Q (WX823), .QN ());
NOR2X1 g59320(.A (n_1176), .B (n_2620), .Y (n_2618));
NOR2X1 g59321(.A (n_1227), .B (n_2620), .Y (n_2617));
NOR2X1 g59330(.A (n_1170), .B (n_2620), .Y (n_2616));
NOR2X1 g59331(.A (n_1066), .B (n_2620), .Y (n_2615));
AND2X1 g62701(.A (WX4574), .B (n_2298), .Y (n_2614));
NOR2X1 g59347(.A (n_1032), .B (n_2620), .Y (n_2613));
NOR2X1 g59352(.A (n_1158), .B (n_2851), .Y (n_2612));
NOR2X1 g59353(.A (n_1119), .B (n_2851), .Y (n_2611));
NOR2X1 g59356(.A (n_1033), .B (n_2605), .Y (n_2610));
NOR2X1 g59357(.A (n_1155), .B (n_2851), .Y (n_2609));
NOR2X1 g59365(.A (n_1019), .B (n_3188), .Y (n_2608));
NOR2X1 g59367(.A (n_1145), .B (n_3188), .Y (n_2607));
NOR2X1 g59376(.A (n_1054), .B (n_2605), .Y (n_2606));
NOR2X1 g59378(.A (n_1136), .B (n_2851), .Y (n_2604));
NOR2X1 g59379(.A (n_1226), .B (n_2851), .Y (n_2603));
NOR2X1 g59386(.A (n_1128), .B (n_2620), .Y (n_2602));
NOR2X1 g59390(.A (n_1055), .B (n_3188), .Y (n_2601));
NOR2X1 g59391(.A (n_1142), .B (n_3188), .Y (n_2600));
NOR2X1 g59394(.A (n_1265), .B (n_2620), .Y (n_2599));
NOR2X1 g59405(.A (n_1108), .B (n_3188), .Y (n_2598));
NOR2X1 g59408(.A (n_1106), .B (n_2851), .Y (n_2597));
NOR2X1 g59409(.A (n_1228), .B (n_2620), .Y (n_2596));
NOR2X1 g59412(.A (n_1102), .B (n_2605), .Y (n_2595));
NOR2X1 g59413(.A (n_1101), .B (n_2851), .Y (n_2594));
NOR2X1 g59414(.A (n_1244), .B (n_3188), .Y (n_2593));
NOR2X1 g59415(.A (n_1182), .B (n_3188), .Y (n_2591));
NOR2X1 g59416(.A (n_1099), .B (n_3188), .Y (n_2590));
NOR2X1 g59422(.A (n_1048), .B (n_3188), .Y (n_2589));
NOR2X1 g59430(.A (n_1086), .B (n_3690), .Y (n_2588));
NOR2X1 g59431(.A (n_1020), .B (n_3690), .Y (n_2587));
NOR2X1 g59434(.A (n_1064), .B (n_3690), .Y (n_2585));
NOR2X1 g59435(.A (n_1084), .B (n_2605), .Y (n_2584));
NOR2X1 g59436(.A (n_1230), .B (n_3690), .Y (n_2583));
NOR2X1 g59437(.A (n_1083), .B (n_3690), .Y (n_2582));
NOR2X1 g59447(.A (n_1264), .B (n_2851), .Y (n_2581));
NOR2X1 g59448(.A (n_1075), .B (n_3690), .Y (n_2579));
NOR2X1 g59449(.A (n_1015), .B (n_3690), .Y (n_2577));
NOR2X1 g59450(.A (n_1074), .B (n_2620), .Y (n_2576));
NOR2X1 g59451(.A (n_1247), .B (n_2851), .Y (n_2575));
NOR2X1 g59452(.A (n_1073), .B (n_2851), .Y (n_2574));
NOR2X1 g59453(.A (n_1072), .B (n_3690), .Y (n_2573));
NOR2X1 g59460(.A (n_1132), .B (n_3690), .Y (n_2572));
NOR2X1 g59464(.A (n_1068), .B (n_2851), .Y (n_2571));
NOR2X1 g59465(.A (n_1113), .B (n_2851), .Y (n_2570));
NOR2X1 g59468(.A (n_1242), .B (n_2851), .Y (n_2568));
NOR2X1 g59469(.A (n_1268), .B (n_2851), .Y (n_2567));
NOR2X1 g59475(.A (n_1035), .B (n_3690), .Y (n_2566));
NOR2X1 g59476(.A (n_1263), .B (n_2851), .Y (n_2565));
NOR2X1 g59477(.A (n_1027), .B (n_2851), .Y (n_2564));
NOR2X1 g59478(.A (n_1168), .B (n_3690), .Y (n_2563));
DFFSRX1 WX779_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1355), .Q (WX779), .QN ());
DFFSRX1 WX819_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1405), .Q (WX819), .QN ());
DFFSRX1 WX771_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1275), .Q (WX771), .QN ());
AND2X1 g62661(.A (WX9740), .B (n_2378), .Y (n_2562));
DFFSRX1 WX891_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1344), .Q (WX891), .QN ());
DFFSRX1 WX879_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1369), .Q (WX879), .QN ());
DFFSRX1 WX863_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1313), .Q (WX863), .QN ());
DFFSRX1 WX773_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1290), .Q (WX773), .QN ());
DFFSRX1 WX805_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1312), .Q (WX805), .QN ());
DFFSRX1 WX2048_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1283), .Q (WX2048), .QN ());
DFFSRX1 WX815_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1307), .Q (WX815), .QN ());
DFFSRX1 WX813_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1311), .Q (WX813), .QN ());
DFFSRX1 WX741_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1367), .Q (WX741), .QN ());
DFFSRX1 WX739_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1372), .Q (WX739), .QN ());
DFFSRX1 WX749_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1403), .Q (WX749), .QN ());
DFFSRX1 WX755_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1396), .Q (WX755), .QN ());
DFFSRX1 WX759_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1402), .Q (WX759), .QN ());
DFFSRX1 WX765_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1291), .Q (WX765), .QN ());
DFFSRX1 WX769_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1441), .Q (WX769), .QN ());
DFFSRX1 WX777_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1322), .Q (WX777), .QN ());
DFFSRX1 WX775_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1306), .Q (WX775), .QN ());
DFFSRX1 WX781_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1462), .Q (WX781), .QN ());
DFFSRX1 WX785_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1426), .Q (WX785), .QN ());
DFFSRX1 WX789_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1334), .Q (WX789), .QN ());
DFFSRX1 WX791_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1414), .Q (WX791), .QN ());
DFFSRX1 WX797_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1385), .Q (WX797), .QN ());
DFFSRX1 WX801_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1325), .Q (WX801), .QN ());
DFFSRX1 WX807_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1391), .Q (WX807), .QN ());
DFFSRX1 WX809_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1308), .Q (WX809), .QN ());
DFFSRX1 WX811_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1356), .Q (WX811), .QN ());
DFFSRX1 WX817_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1386), .Q (WX817), .QN ());
DFFSRX1 WX843_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1387), .Q (WX843), .QN ());
DFFSRX1 WX11053_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1316), .Q (WX11053), .QN ());
DFFSRX1 WX851_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1417), .Q (WX851), .QN ());
DFFSRX1 WX859_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1379), .Q (WX859), .QN ());
DFFSRX1 WX841_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1446), .Q (WX841), .QN ());
DFFSRX1 WX847_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1371), .Q (WX847), .QN ());
DFFSRX1 WX881_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1370), .Q (WX881), .QN ());
DFFSRX1 WX885_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1384), .Q (WX885), .QN ());
DFFSRX1 WX893_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1381), .Q (WX893), .QN ());
DFFSRX1 WX867_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1395), .Q (WX867), .QN ());
DFFSRX1 WX761_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1461), .Q (WX761), .QN ());
DFFSRX1 WX709_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1440), .Q (WX709), .QN ());
DFFSRX1 WX2004_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1336), .Q (WX2004), .QN ());
DFFSRX1 WX2006_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1360), .Q (WX2006), .QN ());
DFFSRX1 WX2010_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1413), .Q (WX2010), .QN ());
DFFSRX1 WX2012_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1358), .Q (WX2012), .QN ());
DFFSRX1 WX2014_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1285), .Q (WX2014), .QN ());
DFFSRX1 WX2018_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1450), .Q (WX2018), .QN ());
DFFSRX1 WX2022_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1420), .Q (WX2022), .QN ());
DFFSRX1 WX2026_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1346), .Q (WX2026), .QN ());
DFFSRX1 WX2034_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1351), .Q (WX2034), .QN ());
DFFSRX1 WX2038_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1349), .Q (WX2038), .QN ());
DFFSRX1 WX2042_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1375), .Q (WX2042), .QN ());
DFFSRX1 WX2046_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1310), .Q (WX2046), .QN ());
DFFSRX1 WX2052_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1443), .Q (WX2052), .QN ());
DFFSRX1 WX2058_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1430), .Q (WX2058), .QN ());
DFFSRX1 WX763_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1317), .Q (WX763), .QN ());
DFFSRX1 WX767_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1352), .Q (WX767), .QN ());
INVX2 g63218(.A (n_6446), .Y (n_2894));
DFFSRX1 WX729_reg(.RN (n_6171), .SN (1'b1), .CK (blif_clk_net), .D(n_1277), .Q (WX729), .QN ());
BUFX3 g63157(.A (n_6437), .Y (n_2897));
AND2X1 g61592(.A (WX7238), .B (n_2527), .Y (n_2559));
AND2X1 g62609(.A (WX8505), .B (n_2346), .Y (n_2558));
AOI21X1 g60399(.A0 (_2100_), .A1 (WX851), .B0 (n_897), .Y (n_2557));
AND2X1 g61587(.A (WX9708), .B (n_2400), .Y (n_2556));
AOI21X1 g60402(.A0 (_2096_), .A1 (WX859), .B0 (n_895), .Y (n_2555));
AOI21X1 g60405(.A0 (_2086_), .A1 (WX879), .B0 (n_900), .Y (n_2554));
AND2X1 g61585(.A (WX11095), .B (n_2346), .Y (n_2553));
AOI21X1 g60428(.A0 (_2106_), .A1 (WX839), .B0 (n_883), .Y (n_2552));
AOI21X1 g60431(.A0 (_2091_), .A1 (WX869), .B0 (n_877), .Y (n_2551));
AOI21X1 g60440(.A0 (_2104_), .A1 (WX843), .B0 (n_885), .Y (n_2548));
AOI21X1 g60449(.A0 (_2098_), .A1 (WX855), .B0 (n_875), .Y (n_2547));
AOI21X1 g60451(.A0 (_2108_), .A1 (WX899), .B0 (n_882), .Y (n_2546));
AOI21X1 g60452(.A0 (_2078_), .A1 (WX895), .B0 (n_1272), .Y (n_2545));
AOI21X1 g60453(.A0 (_2108_), .A1 (WX891), .B0 (n_887), .Y (n_2544));
AOI21X1 g60455(.A0 (_2083_), .A1 (WX885), .B0 (n_901), .Y (n_2543));
AOI21X1 g60456(.A0 (_2084_), .A1 (WX883), .B0 (n_852), .Y (n_2542));
AOI21X1 g60457(.A0 (_2085_), .A1 (WX881), .B0 (n_846), .Y (n_2541));
AOI21X1 g60458(.A0 (_2108_), .A1 (WX877), .B0 (n_898), .Y (n_2540));
AOI21X1 g60459(.A0 (_2088_), .A1 (WX875), .B0 (n_892), .Y (n_2539));
AOI21X1 g60460(.A0 (_2090_), .A1 (WX871), .B0 (n_894), .Y (n_2538));
AOI21X1 g60461(.A0 (_2108_), .A1 (WX867), .B0 (n_878), .Y (n_2537));
AOI21X1 g60462(.A0 (_2093_), .A1 (WX865), .B0 (n_890), .Y (n_2536));
AOI21X1 g60463(.A0 (_2097_), .A1 (WX857), .B0 (n_893), .Y (n_2535));
AND2X1 g61580(.A (WX5941), .B (n_2378), .Y (n_2534));
AOI21X1 g60464(.A0 (_2101_), .A1 (WX849), .B0 (n_873), .Y (n_2533));
AOI21X1 g60465(.A0 (_2103_), .A1 (WX845), .B0 (n_886), .Y (n_2532));
AOI21X1 g60466(.A0 (_2105_), .A1 (WX841), .B0 (n_889), .Y (n_2531));
AND2X1 g61570(.A (WX3339), .B (n_2529), .Y (n_2530));
AND2X1 g61566(.A (WX11081), .B (n_2527), .Y (n_2528));
CLKBUFX3 g63079(.A (n_6624), .Y (n_2840));
AND2X1 g62582(.A (WX5829), .B (n_2378), .Y (n_2525));
AOI21X1 g60623(.A0 (_2079_), .A1 (WX893), .B0 (n_881), .Y (n_2524));
AOI21X1 g60635(.A0 (_2077_), .A1 (WX897), .B0 (n_896), .Y (n_2523));
AOI21X1 g60649(.A0 (_2102_), .A1 (WX847), .B0 (n_888), .Y (n_2522));
AOI21X1 g60650(.A0 (_2099_), .A1 (WX853), .B0 (n_879), .Y (n_2521));
AOI21X1 g60657(.A0 (_2095_), .A1 (WX861), .B0 (n_874), .Y (n_2520));
AOI21X1 g60658(.A0 (_2082_), .A1 (WX887), .B0 (n_884), .Y (n_2519));
AOI21X1 g60662(.A0 (_2094_), .A1 (WX863), .B0 (n_876), .Y (n_2518));
AOI21X1 g60672(.A0 (_2081_), .A1 (WX889), .B0 (n_891), .Y (n_2517));
AOI21X1 g60673(.A0 (_2089_), .A1 (WX873), .B0 (n_899), .Y (n_2516));
AND2X1 g62596(.A (WX5823), .B (n_2527), .Y (n_2515));
NAND2X1 g60710(.A (n_1005), .B (n_1003), .Y (n_2514));
AND2X1 g61558(.A (WX11169), .B (n_2227), .Y (n_2513));
INVX1 g60724(.A (n_2511), .Y (n_2512));
NAND2X1 g60731(.A (n_1002), .B (n_999), .Y (n_2508));
NAND2X1 g60743(.A (n_998), .B (n_908), .Y (n_2505));
AND2X1 g61552(.A (WX9806), .B (n_2383), .Y (n_2504));
NAND2X1 g60764(.A (n_988), .B (n_910), .Y (n_2503));
NAND2X1 g60785(.A (n_986), .B (n_984), .Y (n_2500));
INVX1 g60795(.A (n_2498), .Y (n_2499));
NAND2X1 g60802(.A (n_982), .B (n_980), .Y (n_2497));
XOR2X1 g60804(.A (n_1315), .B (n_2800), .Y (n_2496));
INVX1 g60807(.A (n_2494), .Y (n_2495));
NAND2X1 g60818(.A (n_923), .B (n_941), .Y (n_2493));
NAND2X1 g60830(.A (n_976), .B (n_955), .Y (n_2488));
NAND2X1 g60842(.A (n_6696), .B (n_6697), .Y (n_2487));
NAND2X1 g60863(.A (n_969), .B (n_971), .Y (n_2484));
NAND2X1 g60872(.A (n_949), .B (n_904), .Y (n_2481));
NAND2X1 g60889(.A (n_952), .B (n_950), .Y (n_2480));
NAND2X1 g60896(.A (n_974), .B (n_967), .Y (n_2477));
AND2X1 g61532(.A (WX2004), .B (n_2216), .Y (n_2476));
AND2X1 g61531(.A (WX9714), .B (n_2383), .Y (n_2475));
INVX1 g60902(.A (n_2472), .Y (n_2473));
NAND2X1 g60906(.A (n_903), .B (n_928), .Y (n_2471));
NAND2X1 g60933(.A (n_957), .B (n_915), .Y (n_2470));
INVX1 g60950(.A (n_2468), .Y (n_2469));
INVX1 g60964(.A (n_2466), .Y (n_2467));
NAND2X1 g60968(.A (n_945), .B (n_942), .Y (n_2465));
NAND2X1 g60991(.A (n_939), .B (n_937), .Y (n_2462));
INVX1 g61010(.A (n_2458), .Y (n_2459));
NAND2X1 g61020(.A (n_6698), .B (n_6699), .Y (n_2457));
INVX1 g61057(.A (n_2453), .Y (n_2454));
AND2X1 g55856(.A (WX10831), .B (n_2346), .Y (n_2452));
NAND2X1 g61069(.A (n_933), .B (n_931), .Y (n_2448));
INVX1 g61083(.A (n_2446), .Y (n_2447));
NAND2X1 g61086(.A (n_991), .B (n_926), .Y (n_2445));
INVX1 g61091(.A (n_2443), .Y (n_2444));
AND2X1 g62569(.A (WX8475), .B (n_2188), .Y (n_2442));
AND2X1 g62572(.A (WX11005), .B (n_2339), .Y (n_2441));
NAND2X1 g61138(.A (n_925), .B (n_922), .Y (n_2440));
NAND2X1 g61140(.A (n_921), .B (n_919), .Y (n_2439));
INVX1 g61151(.A (n_2437), .Y (n_2438));
NAND2X1 g61167(.A (n_963), .B (n_960), .Y (n_2434));
AND2X1 g62573(.A (WX3275), .B (n_2227), .Y (n_2433));
NAND2X1 g61179(.A (n_930), .B (n_916), .Y (n_2431));
NAND2X1 g61185(.A (n_918), .B (n_965), .Y (n_2428));
NAND2X1 g61196(.A (n_1007), .B (n_947), .Y (n_2425));
NAND2X1 g61209(.A (n_914), .B (n_912), .Y (n_2424));
INVX1 g61219(.A (n_2422), .Y (n_2423));
NAND2X1 g61229(.A (n_954), .B (n_909), .Y (n_2421));
AND2X1 g62571(.A (WX5901), .B (n_2298), .Y (n_2420));
NAND2X1 g61233(.A (n_993), .B (n_911), .Y (n_2419));
NAND2X1 g61271(.A (n_959), .B (n_907), .Y (n_2412));
NAND2X1 g61295(.A (n_906), .B (n_902), .Y (n_2409));
AND2X1 g62567(.A (WX2036), .B (n_2188), .Y (n_2408));
NAND2X1 g61307(.A (n_996), .B (n_994), .Y (n_2406));
AND2X1 g55860(.A (WX1780), .B (n_2402), .Y (n_2405));
AND2X1 g61521(.A (WX11059), .B (n_2346), .Y (n_2404));
AND2X1 g61523(.A (WX3271), .B (n_2402), .Y (n_2403));
AND2X1 g61524(.A (WX11033), .B (n_2400), .Y (n_2401));
AND2X1 g61526(.A (WX7252), .B (n_2227), .Y (n_2399));
AND2X1 g61527(.A (WX3257), .B (n_2378), .Y (n_2398));
AND2X1 g61528(.A (WX3403), .B (n_2396), .Y (n_2397));
AND2X1 g61529(.A (WX11115), .B (n_2400), .Y (n_2395));
AND2X1 g61530(.A (WX11049), .B (n_2227), .Y (n_2394));
AND2X1 g61533(.A (WX11037), .B (n_2402), .Y (n_2393));
AND2X1 g61535(.A (WX9852), .B (n_2402), .Y (n_2392));
AND2X1 g61537(.A (WX9702), .B (n_2371), .Y (n_2391));
AND2X1 g61539(.A (WX9876), .B (n_2388), .Y (n_2390));
AND2X1 g61540(.A (WX11121), .B (n_2388), .Y (n_2389));
AND2X1 g61541(.A (WX7114), .B (n_2346), .Y (n_2387));
AND2X1 g61546(.A (WX9802), .B (n_2346), .Y (n_2386));
AND2X1 g61550(.A (WX9824), .B (n_2383), .Y (n_2385));
AND2X1 g61551(.A (WX7220), .B (n_2383), .Y (n_2384));
AND2X1 g61554(.A (WX11073), .B (n_2383), .Y (n_2382));
AND2X1 g61555(.A (WX9878), .B (n_2383), .Y (n_2380));
AND2X1 g61556(.A (WX11111), .B (n_2378), .Y (n_2379));
AND2X1 g61561(.A (WX9850), .B (n_2227), .Y (n_2377));
AND2X1 g61562(.A (WX11079), .B (n_2227), .Y (n_2376));
AND2X1 g61563(.A (WX7110), .B (n_2227), .Y (n_2375));
AND2X1 g61564(.A (WX7240), .B (n_2527), .Y (n_2373));
AND2X1 g61568(.A (WX11083), .B (n_2371), .Y (n_2372));
AND2X1 g61571(.A (WX8491), .B (n_2371), .Y (n_2370));
AND2X1 g62556(.A (WX8473), .B (n_2216), .Y (n_2369));
AND2X1 g61578(.A (WX2068), .B (n_2378), .Y (n_2368));
AND2X1 g61581(.A (WX11093), .B (n_2378), .Y (n_2366));
AND2X1 g61582(.A (WX5919), .B (n_2188), .Y (n_2365));
AND2X1 g61583(.A (WX7160), .B (n_2346), .Y (n_2364));
AND2X1 g62560(.A (WX3421), .B (n_2402), .Y (n_2363));
AND2X1 g61586(.A (WX3349), .B (n_2378), .Y (n_2362));
AND2X1 g61589(.A (WX11153), .B (n_2383), .Y (n_2361));
AND2X1 g61591(.A (WX7182), .B (n_2383), .Y (n_2360));
AND2X1 g61594(.A (WX11103), .B (n_2400), .Y (n_2359));
AND2X1 g61595(.A (WX5925), .B (n_2527), .Y (n_2358));
AND2X1 g61596(.A (WX7196), .B (n_2402), .Y (n_2357));
AND2X1 g61597(.A (WX7204), .B (n_2402), .Y (n_2356));
AND2X1 g61598(.A (WX3279), .B (n_2378), .Y (n_2355));
AND2X1 g61599(.A (WX5953), .B (n_2378), .Y (n_2353));
AND2X1 g61600(.A (WX3285), .B (n_2378), .Y (n_2352));
AND2X1 g61601(.A (WX4594), .B (n_2227), .Y (n_2351));
AND2X1 g61606(.A (WX7164), .B (n_2400), .Y (n_2350));
AND2X1 g61610(.A (WX7294), .B (n_2227), .Y (n_2349));
AND2X1 g61611(.A (WX11113), .B (n_2378), .Y (n_2348));
AND2X1 g61613(.A (WX7234), .B (n_2346), .Y (n_2347));
AND2X1 g61615(.A (WX9712), .B (n_2378), .Y (n_2345));
AND2X1 g61616(.A (WX5929), .B (n_2346), .Y (n_2344));
AND2X1 g61617(.A (WX7244), .B (n_2346), .Y (n_2343));
AND2X1 g61618(.A (WX7248), .B (n_2223), .Y (n_2341));
AND2X1 g61619(.A (WX9882), .B (n_2339), .Y (n_2340));
AND2X1 g61620(.A (WX4550), .B (n_2378), .Y (n_2338));
AND2X1 g61623(.A (WX7232), .B (n_2378), .Y (n_2337));
AND2X1 g61625(.A (WX2064), .B (n_2378), .Y (n_2336));
AND2X1 g61626(.A (WX5927), .B (n_2333), .Y (n_2335));
AND2X1 g61627(.A (WX9822), .B (n_2333), .Y (n_2334));
AND2X1 g61629(.A (WX7276), .B (n_2325), .Y (n_2332));
AND2X1 g61630(.A (WX3277), .B (n_2272), .Y (n_2331));
AND2X1 g62555(.A (WX5851), .B (n_2378), .Y (n_2330));
AND2X1 g61632(.A (WX11177), .B (n_2527), .Y (n_2329));
AND2X1 g61634(.A (WX11133), .B (n_2378), .Y (n_2328));
AND2X1 g61639(.A (WX11137), .B (n_2325), .Y (n_2326));
AND2X1 g61641(.A (WX11161), .B (n_2378), .Y (n_2324));
AND2X1 g61642(.A (WX5933), .B (n_2388), .Y (n_2323));
AND2X1 g61644(.A (WX3379), .B (n_2378), .Y (n_2322));
AND2X1 g61649(.A (WX9750), .B (n_2311), .Y (n_2321));
AND2X1 g61653(.A (WX7230), .B (n_2383), .Y (n_2320));
AND2X1 g61654(.A (WX3237), .B (n_2188), .Y (n_2318));
AND2X1 g61656(.A (WX5939), .B (n_2188), .Y (n_2317));
AND2X1 g61658(.A (WX9716), .B (n_2188), .Y (n_2316));
AND2X1 g61661(.A (WX5871), .B (n_2188), .Y (n_2315));
AND2X1 g61664(.A (WX9744), .B (n_2188), .Y (n_2313));
AND2X1 g61666(.A (WX9762), .B (n_2311), .Y (n_2312));
AND2X1 g61667(.A (WX4558), .B (n_2311), .Y (n_2310));
AND2X1 g61668(.A (WX3273), .B (n_2188), .Y (n_2309));
AND2X1 g61670(.A (WX5945), .B (n_2311), .Y (n_2308));
AND2X1 g61671(.A (WX9860), .B (n_2311), .Y (n_2307));
AND2X1 g61672(.A (WX7228), .B (n_2383), .Y (n_2306));
AND2X1 g61673(.A (WX7226), .B (n_2383), .Y (n_2305));
AND2X1 g61680(.A (WX11109), .B (n_2311), .Y (n_2304));
AND2X1 g61681(.A (WX8423), .B (n_2311), .Y (n_2303));
AND2X1 g61682(.A (WX3327), .B (n_2311), .Y (n_2302));
AND2X1 g62551(.A (WX2042), .B (n_2388), .Y (n_2301));
AND2X1 g61686(.A (WX7222), .B (n_2383), .Y (n_2300));
AND2X1 g61687(.A (WX9856), .B (n_2298), .Y (n_2299));
AND2X1 g61689(.A (WX7118), .B (n_2383), .Y (n_2297));
AND2X1 g61690(.A (WX7218), .B (n_2346), .Y (n_2296));
AND2X1 g61691(.A (WX7224), .B (n_2346), .Y (n_2295));
AND2X1 g61693(.A (WX4544), .B (n_2188), .Y (n_2293));
AND2X1 g61694(.A (WX4560), .B (n_2378), .Y (n_2292));
AND2X1 g62549(.A (WX5819), .B (n_2346), .Y (n_2291));
AND2X1 g61697(.A (WX7214), .B (n_2378), .Y (n_2290));
AND2X1 g61698(.A (WX3319), .B (n_2246), .Y (n_2289));
AND2X1 g61700(.A (WX4598), .B (n_2188), .Y (n_2288));
AND2X1 g61701(.A (WX9820), .B (n_2188), .Y (n_2287));
AND2X1 g61702(.A (WX5979), .B (n_2346), .Y (n_2286));
AND2X1 g61703(.A (WX11107), .B (n_2346), .Y (n_2285));
AND2X1 g61704(.A (WX9698), .B (n_2346), .Y (n_2284));
AND2X1 g61706(.A (WX3365), .B (n_2311), .Y (n_2283));
AND2X1 g61707(.A (WX11131), .B (n_2325), .Y (n_2282));
AND2X1 g61708(.A (WX3361), .B (n_2298), .Y (n_2281));
AND2X1 g61711(.A (WX11163), .B (n_2227), .Y (n_2280));
AND2X1 g61712(.A (WX8517), .B (n_2227), .Y (n_2279));
AND2X1 g61714(.A (WX9772), .B (n_2346), .Y (n_2277));
AND2X1 g61717(.A (WX11123), .B (n_2346), .Y (n_2276));
AND2X1 g61719(.A (WX3351), .B (n_2227), .Y (n_2275));
AND2X1 g61720(.A (WX4562), .B (n_2227), .Y (n_2274));
AND2X1 g61721(.A (WX4540), .B (n_2272), .Y (n_2273));
AND2X1 g61724(.A (WX5879), .B (n_2333), .Y (n_2271));
AND2X1 g61725(.A (WX5875), .B (n_2333), .Y (n_2270));
AND2X1 g61728(.A (WX5991), .B (n_2227), .Y (n_2269));
AND2X1 g61729(.A (WX2056), .B (n_2227), .Y (n_2268));
AND2X1 g61731(.A (WX3263), .B (n_2227), .Y (n_2267));
AND2X1 g61732(.A (WX7166), .B (n_2378), .Y (n_2266));
AND2X1 g61733(.A (WX7190), .B (n_2346), .Y (n_2264));
AND2X1 g62544(.A (WX3381), .B (n_2378), .Y (n_2262));
AND2X1 g61739(.A (WX9774), .B (n_2346), .Y (n_2261));
AND2X1 g61741(.A (WX7256), .B (n_2272), .Y (n_2260));
AND2X1 g62542(.A (WX2084), .B (n_2346), .Y (n_2259));
AND2X1 g61743(.A (WX5985), .B (n_2272), .Y (n_2258));
AND2X1 g61744(.A (WX7192), .B (n_2246), .Y (n_2257));
AND2X1 g61745(.A (WX7194), .B (n_2346), .Y (n_2256));
AND2X1 g61746(.A (WX8445), .B (n_2346), .Y (n_2255));
AND2X1 g61747(.A (WX5999), .B (n_2333), .Y (n_2254));
AND2X1 g61749(.A (WX9726), .B (n_2251), .Y (n_2253));
AND2X1 g61750(.A (WX9704), .B (n_2251), .Y (n_2252));
AND2X1 g61751(.A (WX7186), .B (n_2272), .Y (n_2250));
AND2X1 g61752(.A (WX8441), .B (n_2272), .Y (n_2249));
AND2X1 g61753(.A (WX5923), .B (n_2333), .Y (n_2248));
AND2X1 g61754(.A (WX2128), .B (n_2246), .Y (n_2247));
AND2X1 g61755(.A (WX2126), .B (n_2246), .Y (n_2245));
AND2X1 g61759(.A (WX7278), .B (n_2333), .Y (n_2244));
AND2X1 g61761(.A (WX5997), .B (n_2396), .Y (n_2243));
AND2X1 g61762(.A (WX3363), .B (n_2396), .Y (n_2242));
AND2X1 g61765(.A (WX3259), .B (n_2346), .Y (n_2241));
AND2X1 g61768(.A (WX11099), .B (n_2383), .Y (n_2240));
AND2X1 g61769(.A (WX2088), .B (n_2383), .Y (n_2239));
AND2X1 g61770(.A (WX9800), .B (n_2188), .Y (n_2238));
AND2X1 g61772(.A (WX7280), .B (n_2383), .Y (n_2237));
AND2X1 g61773(.A (WX8519), .B (n_2188), .Y (n_2236));
AND2X1 g62539(.A (WX5831), .B (n_2188), .Y (n_2235));
AND2X1 g61777(.A (WX3289), .B (n_2188), .Y (n_2234));
AND2X1 g61778(.A (WX4638), .B (n_2378), .Y (n_2233));
AND2X1 g61781(.A (WX2112), .B (n_2346), .Y (n_2232));
AND2X1 g61783(.A (WX9730), .B (n_2346), .Y (n_2231));
AND2X1 g61784(.A (WX9754), .B (n_2188), .Y (n_2230));
AND2X1 g61790(.A (WX3415), .B (n_2378), .Y (n_2229));
AND2X1 g61791(.A (WX3255), .B (n_2227), .Y (n_2228));
AND2X1 g58615(.A (WX2066), .B (n_2346), .Y (n_2226));
AND2X1 g61794(.A (WX2122), .B (n_2227), .Y (n_2225));
AND2X1 g61795(.A (WX8529), .B (n_2223), .Y (n_2224));
AND2X1 g61796(.A (WX9832), .B (n_2378), .Y (n_2222));
AND2X1 g61797(.A (WX8449), .B (n_2223), .Y (n_2221));
AND2X1 g61799(.A (WX7158), .B (n_2218), .Y (n_2220));
AND2X1 g61800(.A (WX11011), .B (n_2218), .Y (n_2219));
AND2X1 g61802(.A (WX4676), .B (n_2216), .Y (n_2217));
AND2X1 g61803(.A (WX7156), .B (n_2216), .Y (n_2215));
AND2X1 g61805(.A (WX7154), .B (n_2223), .Y (n_2214));
AND2X1 g61807(.A (WX9816), .B (n_2383), .Y (n_2213));
AND2X1 g61809(.A (WX7134), .B (n_2223), .Y (n_2212));
AND2X1 g61810(.A (WX7246), .B (n_2246), .Y (n_2211));
AND2X1 g61811(.A (WX7144), .B (n_2371), .Y (n_2210));
AND2X1 g61812(.A (WX9736), .B (n_2246), .Y (n_2209));
AND2X1 g61816(.A (WX7150), .B (n_2371), .Y (n_2208));
AND2X1 g61820(.A (WX9842), .B (n_2371), .Y (n_2207));
AND2X1 g61823(.A (WX7148), .B (n_2371), .Y (n_2206));
AND2X1 g61825(.A (WX3321), .B (n_2383), .Y (n_2205));
AND2X1 g61826(.A (WX4634), .B (n_2396), .Y (n_2204));
AND2X1 g61827(.A (WX11087), .B (n_2198), .Y (n_2203));
AND2X1 g61828(.A (WX7124), .B (n_2227), .Y (n_2202));
AND2X1 g61829(.A (WX3301), .B (n_2218), .Y (n_2201));
AND2X1 g61832(.A (WX3409), .B (n_2371), .Y (n_2200));
AND2X1 g61834(.A (WX9778), .B (n_2198), .Y (n_2199));
AND2X1 g61835(.A (WX7272), .B (n_2218), .Y (n_2197));
AND2X1 g61837(.A (WX7138), .B (n_2216), .Y (n_2196));
AND2X1 g61838(.A (WX2118), .B (n_2218), .Y (n_2194));
AND2X1 g61839(.A (WX4626), .B (n_2529), .Y (n_2193));
AND2X1 g61840(.A (WX5949), .B (n_2383), .Y (n_2192));
AND2X1 g61847(.A (WX3265), .B (n_2529), .Y (n_2191));
AND2X1 g61848(.A (WX11141), .B (n_2383), .Y (n_2190));
AND2X1 g61849(.A (WX5947), .B (n_2188), .Y (n_2189));
AND2X1 g62536(.A (WX11025), .B (n_2227), .Y (n_2187));
AND2X1 g61850(.A (WX2114), .B (n_2188), .Y (n_2186));
AND2X1 g61851(.A (WX4584), .B (n_2227), .Y (n_2185));
AND2X1 g61854(.A (WX3267), .B (n_2227), .Y (n_2183));
AND2X1 g61855(.A (WX7120), .B (n_2383), .Y (n_2182));
AND2X1 g61856(.A (WX7132), .B (n_2227), .Y (n_2181));
AND2X1 g61858(.A (WX3357), .B (n_2227), .Y (n_2180));
AND2X1 g61859(.A (WX3281), .B (n_2227), .Y (n_2179));
AND2X1 g61861(.A (WX3247), .B (n_2188), .Y (n_2178));
AND2X1 g61863(.A (WX11119), .B (n_2198), .Y (n_2177));
AND2X1 g61864(.A (WX7126), .B (n_2198), .Y (n_2176));
AND2X1 g61865(.A (WX5937), .B (n_2216), .Y (n_2175));
AND2X1 g61866(.A (WX7128), .B (n_2227), .Y (n_2174));
AND2X1 g61867(.A (WX3347), .B (n_2339), .Y (n_2173));
AND2X1 g61868(.A (WX2060), .B (n_2251), .Y (n_2172));
AND2X1 g61869(.A (WX7130), .B (n_2251), .Y (n_2171));
AND2X1 g61870(.A (WX9742), .B (n_2396), .Y (n_2170));
AND2X1 g61871(.A (WX11085), .B (n_2383), .Y (n_2169));
AND2X1 g61873(.A (WX11043), .B (n_2251), .Y (n_2168));
AND2X1 g61874(.A (WX3283), .B (n_2378), .Y (n_2167));
AND2X1 g61877(.A (WX8447), .B (n_2198), .Y (n_2166));
AND2X1 g61879(.A (WX4564), .B (n_2227), .Y (n_2165));
AND2X1 g61881(.A (WX11067), .B (n_2198), .Y (n_2164));
AND2X1 g61883(.A (WX8453), .B (n_2216), .Y (n_2163));
AND2X1 g61884(.A (WX4538), .B (n_2216), .Y (n_2162));
AND2X1 g61886(.A (WX5959), .B (n_2529), .Y (n_2161));
AND2X1 g61887(.A (WX3355), .B (n_2298), .Y (n_2160));
AND2X1 g61890(.A (WX4588), .B (n_2227), .Y (n_2159));
AND2X1 g61891(.A (WX9724), .B (n_2227), .Y (n_2158));
AND2X1 g61892(.A (WX5965), .B (n_2223), .Y (n_2157));
AND2X1 g61893(.A (WX11147), .B (n_2383), .Y (n_2156));
AND2X1 g61894(.A (WX7122), .B (n_2216), .Y (n_2155));
AND2X1 g61900(.A (WX4636), .B (n_2216), .Y (n_2154));
AND2X1 g61901(.A (WX4628), .B (n_2333), .Y (n_2153));
AND2X1 g61902(.A (WX8551), .B (n_2298), .Y (n_2152));
AND2X1 g61904(.A (WX9872), .B (n_2223), .Y (n_2151));
AND2X1 g61905(.A (WX5861), .B (n_2227), .Y (n_2150));
AND2X1 g61906(.A (WX8407), .B (n_2246), .Y (n_2149));
AND2X1 g61907(.A (WX8547), .B (n_2198), .Y (n_2148));
AND2X1 g61915(.A (WX4570), .B (n_2227), .Y (n_2147));
AND2X1 g61917(.A (WX11027), .B (n_2383), .Y (n_2146));
AND2X1 g61919(.A (WX11139), .B (n_2251), .Y (n_2145));
AND2X1 g61920(.A (WX5683), .B (n_2198), .Y (n_2144));
AND2X1 g61921(.A (WX4652), .B (n_2246), .Y (n_2143));
AND2X1 g61925(.A (WX5957), .B (n_2251), .Y (n_2142));
AND2X1 g61926(.A (WX3287), .B (n_2346), .Y (n_2141));
AND2X1 g61929(.A (WX11149), .B (n_2383), .Y (n_2140));
AND2X1 g61931(.A (WX8557), .B (n_2227), .Y (n_2139));
AND2X1 g61932(.A (WX9722), .B (n_2218), .Y (n_2138));
AND2X1 g61933(.A (WX9840), .B (n_2396), .Y (n_2137));
AND2X1 g62534(.A (WX5867), .B (n_2383), .Y (n_2136));
AND2X1 g61935(.A (WX2076), .B (n_2371), .Y (n_2135));
AND2X1 g61936(.A (WX7116), .B (n_2378), .Y (n_2134));
AND2X1 g61937(.A (WX9796), .B (n_2298), .Y (n_2133));
AND2X1 g61938(.A (WX9776), .B (n_2246), .Y (n_2132));
AND2X1 g61939(.A (WX11071), .B (n_2383), .Y (n_2130));
AND2X1 g61943(.A (WX9760), .B (n_2216), .Y (n_2129));
AND2X1 g61944(.A (WX4576), .B (n_2346), .Y (n_2128));
AND2X1 g61947(.A (WX3395), .B (n_2346), .Y (n_2127));
AND2X1 g61948(.A (WX4526), .B (n_2216), .Y (n_2126));
AND2X1 g61949(.A (WX9790), .B (n_2383), .Y (n_2125));
AND2X1 g61950(.A (WX9768), .B (n_2216), .Y (n_2124));
AND2X1 g61952(.A (WX4662), .B (n_2216), .Y (n_2123));
AND2X1 g61953(.A (WX4580), .B (n_2216), .Y (n_2122));
AND2X1 g61955(.A (WX9728), .B (n_2188), .Y (n_2121));
AND2X1 g61956(.A (WX9718), .B (n_2383), .Y (n_2120));
AND2X1 g61957(.A (WX3405), .B (n_2346), .Y (n_2119));
AND2X1 g61958(.A (WX3245), .B (n_2227), .Y (n_2118));
AND2X1 g61959(.A (WX2010), .B (n_2333), .Y (n_2117));
AND2X1 g61961(.A (WX8589), .B (n_2325), .Y (n_2116));
AND2X1 g61962(.A (WX4688), .B (n_2246), .Y (n_2115));
AND2X1 g61963(.A (WX9706), .B (n_2527), .Y (n_2114));
AND2X1 g61965(.A (WX3243), .B (n_2298), .Y (n_2113));
AND2X1 g61966(.A (WX3241), .B (n_2383), .Y (n_2112));
AND2X1 g61967(.A (WX4698), .B (n_2346), .Y (n_2111));
AND2X1 g61968(.A (WX8591), .B (n_2339), .Y (n_2110));
AND2X1 g61969(.A (WX3239), .B (n_2402), .Y (n_2109));
AND2X1 g61970(.A (WX4704), .B (n_2223), .Y (n_2108));
AND2X1 g61971(.A (WX8583), .B (n_2383), .Y (n_2107));
AND2X1 g61972(.A (WX11029), .B (n_2396), .Y (n_2106));
AND2X1 g61973(.A (WX4712), .B (n_2246), .Y (n_2105));
AND2X1 g61976(.A (WX8565), .B (n_2383), .Y (n_2104));
AND2X1 g61978(.A (WX8579), .B (n_2339), .Y (n_2103));
AND2X1 g61980(.A (WX3383), .B (n_2378), .Y (n_2102));
AND2X1 g61981(.A (WX8559), .B (n_2396), .Y (n_2101));
AND2X1 g61982(.A (WX2104), .B (n_2311), .Y (n_2100));
AND2X1 g61983(.A (WX4678), .B (n_2346), .Y (n_2099));
AND2X1 g61985(.A (WX3233), .B (n_2339), .Y (n_2098));
AND2X1 g61986(.A (WX3393), .B (n_2378), .Y (n_2097));
AND2X1 g61987(.A (WX8455), .B (n_2188), .Y (n_2096));
AND2X1 g61988(.A (WX3235), .B (n_2378), .Y (n_2095));
AND2X1 g61990(.A (WX8567), .B (n_2227), .Y (n_2094));
AND2X1 g61992(.A (WX8573), .B (n_2227), .Y (n_2093));
AND2X1 g61994(.A (WX3391), .B (n_2227), .Y (n_2092));
AND2X1 g61995(.A (WX10995), .B (n_2227), .Y (n_2091));
AND2X1 g61996(.A (WX8571), .B (n_2227), .Y (n_2090));
AND2X1 g61997(.A (WX2108), .B (n_2227), .Y (n_2089));
AND2X1 g61998(.A (WX2008), .B (n_2396), .Y (n_2087));
AND2X1 g62000(.A (WX7242), .B (n_2227), .Y (n_2086));
AND2X1 g62001(.A (WX11015), .B (n_2346), .Y (n_2085));
AND2X1 g62002(.A (WX9864), .B (n_2346), .Y (n_2084));
AND2X1 g62003(.A (WX3385), .B (n_2339), .Y (n_2083));
AND2X1 g62004(.A (WX4710), .B (n_2339), .Y (n_2082));
AND2X1 g62009(.A (WX2012), .B (n_2378), .Y (n_2081));
AND2X1 g62010(.A (WX2086), .B (n_2346), .Y (n_2080));
AND2X1 g62011(.A (WX4680), .B (n_2251), .Y (n_2079));
AND2X1 g62012(.A (WX4696), .B (n_2383), .Y (n_2078));
AND2X1 g62013(.A (WX8561), .B (n_2400), .Y (n_2077));
AND2X1 g62014(.A (WX11077), .B (n_2227), .Y (n_2076));
AND2X1 g62015(.A (WX2106), .B (n_2227), .Y (n_2075));
AND2X1 g62016(.A (WX4686), .B (n_2396), .Y (n_2074));
AND2X1 g62017(.A (WX3335), .B (n_2388), .Y (n_2073));
AND2X1 g62018(.A (WX4666), .B (n_2383), .Y (n_2072));
AND2X1 g62019(.A (WX9830), .B (n_2272), .Y (n_2071));
AND2X1 g62020(.A (WX9788), .B (n_2529), .Y (n_2070));
AND2X1 g62021(.A (WX4674), .B (n_2388), .Y (n_2069));
AND2X1 g62022(.A (WX9838), .B (n_2396), .Y (n_2068));
AND2X1 g62023(.A (WX4670), .B (n_2227), .Y (n_2067));
AND2X1 g62024(.A (WX3253), .B (n_2529), .Y (n_2066));
AND2X1 g62025(.A (WX4664), .B (n_2227), .Y (n_2065));
AND2X1 g62026(.A (WX7296), .B (n_2216), .Y (n_2064));
AND2X1 g62027(.A (WX4660), .B (n_2383), .Y (n_2063));
AND2X1 g62030(.A (WX9696), .B (n_2529), .Y (n_2062));
AND2X1 g62033(.A (WX4566), .B (n_2529), .Y (n_2061));
AND2X1 g62034(.A (WX11001), .B (n_2227), .Y (n_2060));
AND2X1 g62036(.A (WX9812), .B (n_2227), .Y (n_2059));
AND2X1 g62038(.A (WX4620), .B (n_2383), .Y (n_2058));
AND2X1 g62041(.A (WX3407), .B (n_2227), .Y (n_2057));
AND2X1 g62043(.A (WX8531), .B (n_2383), .Y (n_2056));
AND2X1 g62044(.A (WX2102), .B (n_2383), .Y (n_2055));
AND2X1 g62047(.A (WX8555), .B (n_2346), .Y (n_2054));
AND2X1 g62048(.A (WX3295), .B (n_2346), .Y (n_2053));
AND2X1 g62050(.A (WX2100), .B (n_2227), .Y (n_2052));
AND2X1 g62052(.A (WX11017), .B (n_2346), .Y (n_2051));
AND2X1 g62055(.A (WX5951), .B (n_2378), .Y (n_2050));
AND2X1 g62057(.A (WX2098), .B (n_2396), .Y (n_2049));
AND2X1 g62058(.A (WX3297), .B (n_2188), .Y (n_2048));
AND2X1 g62059(.A (WX5849), .B (n_2198), .Y (n_2047));
AND2X1 g62060(.A (WX8553), .B (n_2529), .Y (n_2046));
AND2X1 g62529(.A (WX3401), .B (n_2298), .Y (n_2045));
AND2X1 g62061(.A (WX2016), .B (n_2529), .Y (n_2044));
AND2X1 g62062(.A (WX11063), .B (n_2188), .Y (n_2043));
AND2X1 g62064(.A (WX9700), .B (n_2216), .Y (n_2042));
AND2X1 g62065(.A (WX8463), .B (n_2227), .Y (n_2041));
AND2X1 g62066(.A (WX2096), .B (n_2325), .Y (n_2040));
AND2X1 g62067(.A (WX3331), .B (n_2188), .Y (n_2039));
AND2X1 g62068(.A (WX3299), .B (n_2371), .Y (n_2038));
AND2X1 g62072(.A (WX8549), .B (n_2378), .Y (n_2037));
AND2X1 g62075(.A (WX5859), .B (n_2400), .Y (n_2036));
AND2X1 g62076(.A (WX4548), .B (n_2346), .Y (n_2035));
AND2X1 g62077(.A (WX3419), .B (n_2378), .Y (n_2034));
AND2X1 g62078(.A (WX8545), .B (n_2383), .Y (n_2033));
AND2X1 g62080(.A (WX4622), .B (n_2272), .Y (n_2032));
AND2X1 g62081(.A (WX8539), .B (n_2378), .Y (n_2031));
AND2X1 g62082(.A (WX2094), .B (n_2402), .Y (n_2030));
AND2X1 g62084(.A (WX2048), .B (n_2396), .Y (n_2029));
AND2X1 g62086(.A (WX4600), .B (n_2346), .Y (n_2028));
AND2X1 g62087(.A (WX4602), .B (n_2251), .Y (n_2027));
AND2X1 g62088(.A (WX8405), .B (n_2400), .Y (n_2026));
AND2X1 g62089(.A (WX4650), .B (n_2218), .Y (n_2025));
AND2X1 g62090(.A (WX8543), .B (n_2223), .Y (n_2024));
AND2X1 g62091(.A (WX10997), .B (n_2383), .Y (n_2023));
AND2X1 g62092(.A (WX7282), .B (n_2216), .Y (n_2022));
AND2X1 g62094(.A (WX9884), .B (n_2346), .Y (n_2021));
AND2X1 g62096(.A (WX5899), .B (n_2223), .Y (n_2020));
AND2X1 g62098(.A (WX4616), .B (n_2346), .Y (n_2019));
AND2X1 g62099(.A (WX8457), .B (n_2402), .Y (n_2018));
AND2X1 g62100(.A (WX5855), .B (n_2339), .Y (n_2017));
AND2X1 g62101(.A (WX8435), .B (n_2388), .Y (n_2016));
AND2X1 g62104(.A (WX8537), .B (n_2402), .Y (n_2015));
AND2X1 g62106(.A (WX9854), .B (n_2188), .Y (n_2014));
AND2X1 g62107(.A (WX10999), .B (n_2388), .Y (n_2013));
AND2X1 g62108(.A (WX7250), .B (n_2383), .Y (n_2012));
AND2X1 g62531(.A (WX2006), .B (n_2188), .Y (n_2011));
AND2X1 g62113(.A (WX3387), .B (n_2527), .Y (n_2010));
AND2X1 g62116(.A (WX8535), .B (n_2272), .Y (n_2009));
AND2X1 g62117(.A (WX7212), .B (n_2402), .Y (n_2008));
AND2X1 g62118(.A (WX5981), .B (n_2378), .Y (n_2007));
AND2X1 g62119(.A (WX4586), .B (n_2272), .Y (n_2006));
AND2X1 g62120(.A (WX4656), .B (n_2383), .Y (n_2005));
AND2X1 g62121(.A (WX3333), .B (n_2188), .Y (n_2004));
AND2X1 g62122(.A (WX9826), .B (n_2383), .Y (n_2003));
AND2X1 g62124(.A (WX2092), .B (n_2311), .Y (n_2002));
AND2X1 g62126(.A (WX4624), .B (n_2388), .Y (n_2001));
AND2X1 g62127(.A (WX7136), .B (n_2388), .Y (n_2000));
AND2X1 g62128(.A (WX7268), .B (n_2346), .Y (n_1999));
AND2X1 g62129(.A (WX4642), .B (n_2527), .Y (n_1998));
AND2X1 g62130(.A (WX8409), .B (n_2346), .Y (n_1997));
AND2X1 g62131(.A (WX4618), .B (n_2246), .Y (n_1996));
AND2X1 g62132(.A (WX4612), .B (n_2298), .Y (n_1995));
AND2X1 g62133(.A (WX7292), .B (n_2378), .Y (n_1994));
AND2X1 g62135(.A (WX3231), .B (n_2378), .Y (n_1993));
AND2X1 g62136(.A (WX8489), .B (n_2346), .Y (n_1992));
AND2X1 g62138(.A (WX8525), .B (n_2325), .Y (n_1991));
AND2X1 g62140(.A (WX11159), .B (n_2346), .Y (n_1990));
AND2X1 g62143(.A (WX3367), .B (n_2383), .Y (n_1989));
AND2X1 g62144(.A (WX11061), .B (n_2227), .Y (n_1988));
AND2X1 g62148(.A (WX4392), .B (n_2227), .Y (n_1987));
AND2X1 g62149(.A (WX8569), .B (n_2188), .Y (n_1986));
AND2X1 g62150(.A (WX11125), .B (n_2246), .Y (n_1985));
AND2X1 g62155(.A (WX8413), .B (n_2246), .Y (n_1984));
AND2X1 g62156(.A (WX2062), .B (n_2272), .Y (n_1983));
AND2X1 g62158(.A (WX9758), .B (n_2251), .Y (n_1982));
AND2X1 g62160(.A (WX3397), .B (n_2346), .Y (n_1981));
AND2X1 g62161(.A (WX7300), .B (n_2346), .Y (n_1980));
AND2X1 g62162(.A (WX6003), .B (n_2333), .Y (n_1979));
AND2X1 g62164(.A (WX4646), .B (n_2333), .Y (n_1978));
AND2X1 g62165(.A (WX9880), .B (n_2346), .Y (n_1977));
AND2X1 g62166(.A (WX7258), .B (n_2325), .Y (n_1976));
AND2X1 g62167(.A (WX8593), .B (n_2227), .Y (n_1975));
AND2X1 g62168(.A (WX11057), .B (n_2227), .Y (n_1974));
AND2X1 g62172(.A (WX3371), .B (n_2346), .Y (n_1973));
AND2X1 g62175(.A (WX8411), .B (n_2227), .Y (n_1972));
AND2X1 g62176(.A (WX9836), .B (n_2227), .Y (n_1971));
AND2X1 g62177(.A (WX11055), .B (n_2378), .Y (n_1970));
AND2X1 g62178(.A (WX8467), .B (n_2227), .Y (n_1969));
AND2X1 g62180(.A (WX9870), .B (n_2378), .Y (n_1968));
AND2X1 g62182(.A (WX7264), .B (n_2227), .Y (n_1967));
AND2X1 g62183(.A (WX4604), .B (n_2223), .Y (n_1966));
AND2X1 g62184(.A (WX9804), .B (n_2218), .Y (n_1965));
AND2X1 g62185(.A (WX8429), .B (n_2527), .Y (n_1964));
AND2X1 g62188(.A (WX5877), .B (n_2188), .Y (n_1963));
AND2X1 g62189(.A (WX6001), .B (n_2378), .Y (n_1962));
AND2X1 g62190(.A (WX8521), .B (n_2378), .Y (n_1961));
AND2X1 g62191(.A (WX7270), .B (n_2216), .Y (n_1960));
AND2X1 g62194(.A (WX5989), .B (n_2218), .Y (n_1959));
AND2X1 g62195(.A (WX5993), .B (n_2383), .Y (n_1958));
AND2X1 g62196(.A (WX3303), .B (n_2198), .Y (n_1957));
AND2X1 g62197(.A (WX7142), .B (n_2216), .Y (n_1956));
AND2X1 g62201(.A (WX9756), .B (n_2383), .Y (n_1955));
AND2X1 g62202(.A (WX7260), .B (n_2216), .Y (n_1954));
AND2X1 g62203(.A (WX5903), .B (n_2383), .Y (n_1953));
AND2X1 g62205(.A (WX11065), .B (n_2223), .Y (n_1951));
AND2X1 g62206(.A (WX4534), .B (n_2223), .Y (n_1950));
AND2X1 g62207(.A (WX4546), .B (n_2383), .Y (n_1949));
AND2X1 g62208(.A (WX2074), .B (n_2346), .Y (n_1948));
AND2X1 g62209(.A (WX8483), .B (n_2383), .Y (n_1947));
AND2X1 g62210(.A (WX3307), .B (n_2227), .Y (n_1946));
AND2X1 g62211(.A (WX9866), .B (n_2378), .Y (n_1945));
AND2X1 g62218(.A (WX4582), .B (n_2216), .Y (n_1944));
AND2X1 g62222(.A (WX4640), .B (n_2383), .Y (n_1943));
AND2X1 g62224(.A (WX4596), .B (n_2383), .Y (n_1942));
AND2X1 g62229(.A (WX7298), .B (n_2227), .Y (n_1941));
AND2X1 g62230(.A (WX2078), .B (n_2227), .Y (n_1940));
AND2X1 g62231(.A (WX2038), .B (n_2227), .Y (n_1939));
AND2X1 g62233(.A (WX11003), .B (n_2378), .Y (n_1938));
AND2X1 g62236(.A (WX5881), .B (n_2346), .Y (n_1937));
AND2X1 g62237(.A (WX4644), .B (n_2383), .Y (n_1936));
AND2X1 g62238(.A (WX2120), .B (n_2378), .Y (n_1935));
AND2X1 g62240(.A (WX4654), .B (n_2371), .Y (n_1934));
AND2X1 g62241(.A (WX3353), .B (n_2383), .Y (n_1933));
AND2X1 g62243(.A (WX5983), .B (n_2383), .Y (n_1932));
AND2X1 g62244(.A (WX4572), .B (n_2383), .Y (n_1931));
AND2X1 g62245(.A (WX8427), .B (n_2346), .Y (n_1930));
AND2X1 g62247(.A (WX4684), .B (n_2339), .Y (n_1929));
AND2X1 g62248(.A (WX4694), .B (n_2346), .Y (n_1928));
AND2X1 g62252(.A (WX9886), .B (n_2227), .Y (n_1927));
AND2X1 g62253(.A (WX4552), .B (n_2227), .Y (n_1926));
AND2X1 g62255(.A (WX4606), .B (n_2378), .Y (n_1925));
AND2X1 g62256(.A (WX4536), .B (n_2227), .Y (n_1924));
AND2X1 g62258(.A (WX5975), .B (n_2188), .Y (n_1923));
AND2X1 g62259(.A (WX2110), .B (n_2402), .Y (n_1922));
AND2X1 g62260(.A (WX7274), .B (n_2346), .Y (n_1921));
AND2X1 g62261(.A (WX5977), .B (n_2272), .Y (n_1920));
AND2X1 g62262(.A (WX3417), .B (n_2378), .Y (n_1919));
AND2X1 g62263(.A (WX8507), .B (n_2371), .Y (n_1918));
AND2X1 g62264(.A (WX9720), .B (n_2383), .Y (n_1917));
AND2X1 g62265(.A (WX5971), .B (n_2346), .Y (n_1916));
AND2X1 g62267(.A (WX5967), .B (n_2227), .Y (n_1915));
AND2X1 g62269(.A (WX7146), .B (n_2383), .Y (n_1914));
AND2X1 g62270(.A (WX8541), .B (n_2198), .Y (n_1913));
AND2X1 g62272(.A (WX5969), .B (n_2346), .Y (n_1912));
AND2X1 g62274(.A (WX3373), .B (n_2371), .Y (n_1911));
AND2X1 g62277(.A (WX5963), .B (n_2333), .Y (n_1910));
AND2X1 g62279(.A (WX8513), .B (n_2346), .Y (n_1909));
AND2X1 g62280(.A (WX8509), .B (n_2383), .Y (n_1908));
AND2X1 g62281(.A (WX8433), .B (n_2383), .Y (n_1907));
AND2X1 g62283(.A (WX11047), .B (n_2346), .Y (n_1906));
AND2X1 g62285(.A (WX5961), .B (n_2198), .Y (n_1905));
AND2X1 g62286(.A (WX8511), .B (n_2298), .Y (n_1904));
AND2X1 g62288(.A (WX8431), .B (n_2198), .Y (n_1903));
AND2X1 g62289(.A (WX7286), .B (n_2216), .Y (n_1902));
AND2X1 g62290(.A (WX7288), .B (n_2216), .Y (n_1901));
AND2X1 g62291(.A (WX3101), .B (n_2216), .Y (n_1900));
AND2X1 g62294(.A (WX3343), .B (n_2227), .Y (n_1899));
AND2X1 g62295(.A (WX7112), .B (n_2371), .Y (n_1898));
AND2X1 g62296(.A (WX9766), .B (n_2227), .Y (n_1897));
AND2X1 g62297(.A (WX3315), .B (n_2383), .Y (n_1896));
AND2X1 g62298(.A (WX2070), .B (n_2198), .Y (n_1895));
AND2X1 g62299(.A (WX11091), .B (n_2339), .Y (n_1894));
AND2X1 g62303(.A (WX3377), .B (n_2218), .Y (n_1893));
AND2X1 g62305(.A (WX5943), .B (n_2227), .Y (n_1892));
AND2X1 g62306(.A (WX8479), .B (n_2227), .Y (n_1891));
AND2X1 g62311(.A (WX8439), .B (n_2346), .Y (n_1890));
AND2X1 g62312(.A (WX9738), .B (n_2251), .Y (n_1889));
AND2X1 g62313(.A (WX9858), .B (n_2383), .Y (n_1888));
AND2X1 g62528(.A (WX9834), .B (n_2527), .Y (n_1887));
AND2X1 g62314(.A (WX7216), .B (n_2325), .Y (n_1886));
AND2X1 g62315(.A (WX2022), .B (n_2246), .Y (n_1885));
AND2X1 g62316(.A (WX4702), .B (n_2527), .Y (n_1884));
AND2X1 g62317(.A (WX4524), .B (n_2527), .Y (n_1883));
AND2X1 g62318(.A (WX5853), .B (n_2529), .Y (n_1882));
AND2X1 g62319(.A (WX5889), .B (n_2227), .Y (n_1881));
AND2X1 g62320(.A (WX8477), .B (n_2378), .Y (n_1880));
AND2X1 g62322(.A (WX4608), .B (n_2227), .Y (n_1879));
AND2X1 g62324(.A (WX5915), .B (n_2216), .Y (n_1878));
AND2X1 g62325(.A (WX8495), .B (n_2371), .Y (n_1877));
AND2X1 g62326(.A (WX3313), .B (n_2198), .Y (n_1876));
AND2X1 g62327(.A (WX8437), .B (n_2216), .Y (n_1875));
AND2X1 g62329(.A (WX5935), .B (n_2246), .Y (n_1874));
AND2X1 g62331(.A (WX8501), .B (n_2246), .Y (n_1873));
AND2X1 g62332(.A (WX11009), .B (n_2218), .Y (n_1872));
AND2X1 g62333(.A (WX5931), .B (n_2218), .Y (n_1871));
AND2X1 g62335(.A (WX4590), .B (n_2246), .Y (n_1870));
AND2X1 g62336(.A (WX2124), .B (n_2378), .Y (n_1869));
AND2X1 g62341(.A (WX9792), .B (n_2216), .Y (n_1868));
AND2X1 g62344(.A (WX8499), .B (n_2378), .Y (n_1867));
AND2X1 g62345(.A (WX10991), .B (n_2383), .Y (n_1866));
AND2X1 g62348(.A (WX7162), .B (n_2227), .Y (n_1865));
AND2X1 g62349(.A (WX3411), .B (n_2188), .Y (n_1864));
AND2X1 g62350(.A (WX8497), .B (n_2246), .Y (n_1863));
AND2X1 g62354(.A (WX5917), .B (n_2246), .Y (n_1862));
AND2X1 g62355(.A (WX11157), .B (n_2383), .Y (n_1861));
AND2X1 g62362(.A (WX8493), .B (n_2227), .Y (n_1860));
AND2X1 g62363(.A (WX9828), .B (n_2227), .Y (n_1859));
AND2X1 g62364(.A (WX5911), .B (n_2378), .Y (n_1858));
AND2X1 g62367(.A (WX2040), .B (n_2346), .Y (n_1857));
AND2X1 g62369(.A (WX8487), .B (n_2251), .Y (n_1856));
AND2X1 g62370(.A (WX5913), .B (n_2333), .Y (n_1855));
AND2X1 g62372(.A (WX5905), .B (n_2325), .Y (n_1854));
AND2X1 g62373(.A (WX3345), .B (n_2188), .Y (n_1853));
AND2X1 g62374(.A (WX9748), .B (n_2346), .Y (n_1852));
AND2X1 g62376(.A (WX2058), .B (n_2227), .Y (n_1851));
AND2X1 g62518(.A (WX8461), .B (n_2378), .Y (n_1850));
AND2X1 g62519(.A (WX3329), .B (n_2400), .Y (n_1849));
AND2X1 g62521(.A (WX9734), .B (n_2383), .Y (n_1848));
AND2X1 g62515(.A (WX5883), .B (n_2396), .Y (n_1847));
AND2X1 g62517(.A (WX9868), .B (n_2400), .Y (n_1846));
AND2X1 g62513(.A (WX8417), .B (n_2333), .Y (n_1845));
AND2X1 g62510(.A (WX4714), .B (n_2346), .Y (n_1844));
AND2X1 g62504(.A (WX2090), .B (n_2346), .Y (n_1843));
AND2X1 g62503(.A (WX8421), .B (n_2346), .Y (n_1842));
AND2X1 g62502(.A (WX4554), .B (n_2346), .Y (n_1841));
AND2X1 g62501(.A (WX7168), .B (n_2378), .Y (n_1840));
AND2X1 g62467(.A (WX5907), .B (n_2378), .Y (n_1838));
AND2X1 g62468(.A (WX3249), .B (n_2227), .Y (n_1837));
AND2X1 g62470(.A (WX4630), .B (n_2378), .Y (n_1836));
AND2X1 g62471(.A (WX5895), .B (n_2246), .Y (n_1835));
AND2X1 g62472(.A (WX5887), .B (n_2346), .Y (n_1834));
AND2X1 g62475(.A (WX8403), .B (n_2298), .Y (n_1833));
AND2X1 g62499(.A (WX2024), .B (n_2388), .Y (n_1832));
AND2X1 g62480(.A (WX5897), .B (n_2325), .Y (n_1831));
AND2X1 g62481(.A (WX11173), .B (n_2246), .Y (n_1830));
AND2X1 g62482(.A (WX8425), .B (n_2383), .Y (n_1829));
AND2X1 g62483(.A (WX7170), .B (n_2378), .Y (n_1828));
AND2X1 g62484(.A (WX8465), .B (n_2298), .Y (n_1827));
AND2X1 g62485(.A (WX4530), .B (n_2311), .Y (n_1826));
AND2X1 g62492(.A (WX5891), .B (n_2339), .Y (n_1825));
AND2X1 g62495(.A (WX11097), .B (n_2325), .Y (n_1824));
AND2X1 g62496(.A (WX2116), .B (n_2402), .Y (n_1823));
AND2X1 g62497(.A (WX11151), .B (n_2339), .Y (n_1822));
AND2X1 g62500(.A (WX4706), .B (n_2402), .Y (n_1821));
AND2X1 g62509(.A (WX9784), .B (n_2188), .Y (n_1820));
AND2X1 g62511(.A (WX11013), .B (n_2346), .Y (n_1819));
AND2X1 g62512(.A (WX2052), .B (n_2378), .Y (n_1818));
AND2X1 g62514(.A (WX3341), .B (n_2227), .Y (n_1817));
AND2X1 g62516(.A (WX3323), .B (n_2298), .Y (n_1816));
AND2X1 g62523(.A (WX7176), .B (n_2227), .Y (n_1815));
AND2X1 g62526(.A (WX2018), .B (n_2378), .Y (n_1814));
AND2X1 g62533(.A (WX8503), .B (n_2346), .Y (n_1813));
AND2X1 g62535(.A (WX6005), .B (n_2188), .Y (n_1812));
AND2X1 g62540(.A (WX5955), .B (n_2346), .Y (n_1811));
AND2X1 g62541(.A (WX8523), .B (n_2383), .Y (n_1810));
AND2X1 g62545(.A (WX5865), .B (n_2378), .Y (n_1809));
AND2X1 g62547(.A (WX5885), .B (n_2188), .Y (n_1808));
AND2X1 g62552(.A (WX7178), .B (n_2388), .Y (n_1807));
AND2X1 g62557(.A (WX4578), .B (n_2223), .Y (n_1806));
AND2X1 g62562(.A (WX9732), .B (n_2218), .Y (n_1805));
AND2X1 g62563(.A (WX11127), .B (n_2246), .Y (n_1804));
AND2X1 g62564(.A (WX5847), .B (n_2227), .Y (n_1803));
AND2X1 g62565(.A (WX8469), .B (n_2223), .Y (n_1802));
AND2X1 g62494(.A (WX2028), .B (n_2388), .Y (n_1801));
AND2X1 g62570(.A (WX11021), .B (n_2378), .Y (n_1800));
AND2X1 g62574(.A (WX4632), .B (n_2378), .Y (n_1799));
AND2X1 g62576(.A (WX5841), .B (n_2188), .Y (n_1798));
AND2X1 g62577(.A (WX5973), .B (n_2346), .Y (n_1797));
AND2X1 g62581(.A (WX11019), .B (n_2227), .Y (n_1796));
AND2X1 g62585(.A (WX5833), .B (n_2251), .Y (n_1795));
AND2X1 g62586(.A (WX5995), .B (n_2383), .Y (n_1794));
AND2X1 g62588(.A (WX3261), .B (n_2378), .Y (n_1793));
AND2X1 g62589(.A (WX7184), .B (n_2227), .Y (n_1792));
AND2X1 g62593(.A (WX11165), .B (n_2298), .Y (n_1791));
AND2X1 g62594(.A (WX8419), .B (n_2298), .Y (n_1790));
AND2X1 g62597(.A (WX5857), .B (n_2383), .Y (n_1789));
AND2X1 g62599(.A (WX4528), .B (n_2218), .Y (n_1788));
AND2X1 g62600(.A (WX5843), .B (n_2388), .Y (n_1787));
AND2X1 g62601(.A (WX5827), .B (n_2400), .Y (n_1786));
AND2X1 g62602(.A (WX7254), .B (n_2188), .Y (n_1785));
AND2X1 g62603(.A (WX5835), .B (n_2272), .Y (n_1784));
AND2X1 g62605(.A (WX3293), .B (n_2400), .Y (n_1783));
AND2X1 g62606(.A (WX9846), .B (n_2333), .Y (n_1782));
AND2X1 g62487(.A (WX5893), .B (n_2325), .Y (n_1781));
AND2X1 g62608(.A (WX9814), .B (n_2216), .Y (n_1780));
AND2X1 g62489(.A (WX2050), .B (n_2388), .Y (n_1779));
AND2X1 g62610(.A (WX4658), .B (n_2402), .Y (n_1778));
AND2X1 g62612(.A (WX5825), .B (n_2388), .Y (n_1777));
AND2X1 g62614(.A (WX3399), .B (n_2246), .Y (n_1776));
AND2X1 g62617(.A (WX8471), .B (n_2378), .Y (n_1775));
AND2X1 g62620(.A (WX7290), .B (n_2227), .Y (n_1774));
AND2X1 g62621(.A (WX11101), .B (n_2227), .Y (n_1773));
AND2X1 g62624(.A (WX8459), .B (n_2378), .Y (n_1772));
AND2X1 g62626(.A (WX4668), .B (n_2383), .Y (n_1771));
AND2X1 g62627(.A (WX4614), .B (n_2246), .Y (n_1770));
AND2X1 g62629(.A (WX4672), .B (n_2216), .Y (n_1769));
AND2X1 g62630(.A (WX9844), .B (n_2227), .Y (n_1768));
AND2X1 g62633(.A (WX3325), .B (n_2227), .Y (n_1767));
AND2X1 g62637(.A (WX9746), .B (n_2346), .Y (n_1766));
AND2X1 g62486(.A (WX7172), .B (n_2246), .Y (n_1765));
AND2X1 g62640(.A (WX8451), .B (n_2529), .Y (n_1764));
AND2X1 g62642(.A (WX5909), .B (n_2246), .Y (n_1763));
AND2X1 g62643(.A (WX8515), .B (n_2378), .Y (n_1762));
AND2X1 g62646(.A (WX7236), .B (n_2251), .Y (n_1761));
AND2X1 g62647(.A (WX4700), .B (n_2188), .Y (n_1760));
AND2X1 g62649(.A (WX4692), .B (n_2378), .Y (n_1759));
AND2X1 g62653(.A (WX8443), .B (n_2298), .Y (n_1758));
AND2X1 g62656(.A (WX2032), .B (n_2227), .Y (n_1757));
AND2X1 g62658(.A (WX11023), .B (n_2378), .Y (n_1756));
AND2X1 g62660(.A (WX3317), .B (n_2346), .Y (n_1755));
AND2X1 g62662(.A (WX2014), .B (n_2227), .Y (n_1754));
AND2X1 g62664(.A (WX2020), .B (n_2378), .Y (n_1753));
AND2X1 g62665(.A (WX6007), .B (n_2218), .Y (n_1752));
AND2X1 g62667(.A (WX4708), .B (n_2378), .Y (n_1751));
AND2X1 g62669(.A (WX2044), .B (n_2383), .Y (n_1750));
AND2X1 g62670(.A (WX2046), .B (n_2346), .Y (n_1749));
AND2X1 g62672(.A (WX2054), .B (n_2246), .Y (n_1748));
AND2X1 g62674(.A (WX5869), .B (n_2272), .Y (n_1747));
AND2X1 g62675(.A (WX11179), .B (n_2346), .Y (n_1746));
AND2X1 g62677(.A (WX11145), .B (n_2272), .Y (n_1745));
AND2X1 g62679(.A (WX2080), .B (n_2246), .Y (n_1744));
AND2X1 g62681(.A (WX2030), .B (n_2346), .Y (n_1743));
AND2X1 g62682(.A (WX11075), .B (n_2325), .Y (n_1742));
AND2X1 g62684(.A (WX3311), .B (n_2188), .Y (n_1741));
AND2X1 g62685(.A (WX9818), .B (n_2311), .Y (n_1740));
AND2X1 g62687(.A (WX2026), .B (n_2188), .Y (n_1739));
AND2X1 g62690(.A (WX5839), .B (n_2378), .Y (n_1738));
AND2X1 g62693(.A (WX11007), .B (n_2339), .Y (n_1737));
AND2X1 g62698(.A (WX8563), .B (n_2383), .Y (n_1736));
AND2X1 g62699(.A (WX3309), .B (n_2339), .Y (n_1735));
AND2X1 g62703(.A (WX8415), .B (n_2339), .Y (n_1734));
AND2X1 g62704(.A (WX9810), .B (n_2378), .Y (n_1733));
AND2X1 g62709(.A (WX3269), .B (n_2188), .Y (n_1732));
AND2X1 g62710(.A (WX7200), .B (n_2346), .Y (n_1731));
AND2X1 g62714(.A (WX7174), .B (n_2400), .Y (n_1730));
AND2X1 g62717(.A (WX8581), .B (n_2400), .Y (n_1729));
AND2X1 g62718(.A (WX5845), .B (n_2227), .Y (n_1728));
AND2X1 g62720(.A (WX9782), .B (n_2188), .Y (n_1727));
AND2X1 g62723(.A (WX8485), .B (n_2216), .Y (n_1726));
AND2X1 g62725(.A (WX8575), .B (n_2383), .Y (n_1725));
AND2X1 g62726(.A (WX8481), .B (n_2188), .Y (n_1724));
AND2X1 g62729(.A (WX4532), .B (n_2378), .Y (n_1723));
AND2X1 g62731(.A (WX11031), .B (n_2188), .Y (n_1722));
AND2X1 g62733(.A (WX7210), .B (n_2227), .Y (n_1721));
AND2X1 g62737(.A (WX6974), .B (n_2529), .Y (n_1720));
AND2X1 g62738(.A (WX7206), .B (n_2311), .Y (n_1719));
AND2X1 g62748(.A (WX3413), .B (n_2529), .Y (n_1718));
AND2X1 g62753(.A (WX3291), .B (n_2383), .Y (n_1717));
AND2X1 g62759(.A (WX4568), .B (n_2383), .Y (n_1716));
AND2X1 g62763(.A (WX11035), .B (n_2216), .Y (n_1715));
AND2X1 g62767(.A (WX3251), .B (n_2227), .Y (n_1714));
AND2X1 g62613(.A (WX7188), .B (n_2378), .Y (n_1713));
AND2X1 g61862(.A (WX9798), .B (n_2188), .Y (n_1712));
AND2X1 g62766(.A (WX11039), .B (n_2396), .Y (n_1711));
AND2X1 g62760(.A (WX8527), .B (n_2218), .Y (n_1710));
AND2X1 g62758(.A (WX7266), .B (n_2227), .Y (n_1709));
AND2X1 g62749(.A (WX8577), .B (n_2529), .Y (n_1708));
AND2X1 g62747(.A (WX10993), .B (n_2227), .Y (n_1707));
NOR2X1 g57543(.A (n_847), .B (n_1648), .Y (n_1706));
AND2X1 g62719(.A (WX5873), .B (n_2400), .Y (n_1702));
AND2X1 g61763(.A (WX5921), .B (n_2188), .Y (n_1701));
AND2X1 g61766(.A (WX9780), .B (n_2188), .Y (n_1700));
AND2X1 g62257(.A (WX7140), .B (n_2251), .Y (n_1699));
AND2X1 g62715(.A (WX3389), .B (n_2246), .Y (n_1698));
NOR2X1 g59240(.A (n_1190), .B (n_5712), .Y (n_1697));
NOR2X1 g59241(.A (n_1172), .B (n_5181), .Y (n_1696));
NOR2X1 g59243(.A (n_1077), .B (n_1425), .Y (n_1694));
NOR2X1 g59245(.A (n_1149), .B (n_1425), .Y (n_1693));
NOR2X1 g59246(.A (n_1185), .B (n_1425), .Y (n_1691));
NOR2X1 g59252(.A (n_1118), .B (n_1425), .Y (n_1690));
NOR2X1 g59253(.A (n_1049), .B (n_1425), .Y (n_1688));
NOR2X1 g59254(.A (n_1147), .B (n_5712), .Y (n_1687));
NOR2X1 g59255(.A (n_1109), .B (n_5712), .Y (n_1685));
NOR2X1 g59256(.A (n_1216), .B (n_1648), .Y (n_1684));
NOR2X1 g59259(.A (n_1194), .B (n_5181), .Y (n_1682));
NOR2X1 g59260(.A (n_1218), .B (n_5181), .Y (n_1681));
NOR2X1 g59261(.A (n_1267), .B (n_5181), .Y (n_1679));
AND2X1 g62711(.A (WX9752), .B (n_2227), .Y (n_1678));
NOR2X1 g59263(.A (n_1239), .B (n_1648), .Y (n_1677));
NOR2X1 g59264(.A (n_1229), .B (n_1425), .Y (n_1676));
NOR2X1 g59265(.A (n_1123), .B (n_5181), .Y (n_1675));
NOR2X1 g59267(.A (n_1217), .B (n_1648), .Y (n_1673));
AND2X1 g61757(.A (WX7180), .B (n_2246), .Y (n_1672));
AND2X1 g62700(.A (WX9710), .B (n_2378), .Y (n_1671));
NOR2X1 g59287(.A (n_1022), .B (n_5181), .Y (n_1670));
NOR2X1 g59288(.A (n_1209), .B (n_5181), .Y (n_1669));
NOR2X1 g59289(.A (n_1059), .B (n_5712), .Y (n_1668));
NOR2X1 g59290(.A (n_1208), .B (n_5712), .Y (n_1666));
NOR2X1 g59291(.A (n_1058), .B (n_5712), .Y (n_1665));
NOR2X1 g59292(.A (n_1207), .B (n_1425), .Y (n_1664));
NOR2X1 g59295(.A (n_1204), .B (n_1648), .Y (n_1662));
NOR2X1 g59296(.A (n_1060), .B (n_1648), .Y (n_1661));
NOR2X1 g59297(.A (n_1203), .B (n_1648), .Y (n_1660));
NOR2X1 g59298(.A (n_1202), .B (n_5712), .Y (n_1659));
NOR2X1 g59299(.A (n_1201), .B (n_5712), .Y (n_1658));
NOR2X1 g59300(.A (n_1045), .B (n_5181), .Y (n_1656));
NOR2X1 g59301(.A (n_1030), .B (n_5181), .Y (n_1655));
NOR2X1 g59302(.A (n_1199), .B (n_1425), .Y (n_1654));
NOR2X1 g59303(.A (n_1014), .B (n_1425), .Y (n_1652));
NOR2X1 g59304(.A (n_1250), .B (n_1648), .Y (n_1651));
NOR2X1 g59305(.A (n_1196), .B (n_1648), .Y (n_1650));
NOR2X1 g59306(.A (n_1062), .B (n_1648), .Y (n_1649));
NOR2X1 g59307(.A (n_1193), .B (n_1648), .Y (n_1647));
NOR2X1 g59308(.A (n_1192), .B (n_5181), .Y (n_1646));
NOR2X1 g59309(.A (n_1191), .B (n_5712), .Y (n_1645));
NOR2X1 g59310(.A (n_1188), .B (n_1648), .Y (n_1644));
NOR2X1 g59311(.A (n_1187), .B (n_1648), .Y (n_1642));
NOR2X1 g59312(.A (n_1251), .B (n_5712), .Y (n_1641));
NOR2X1 g59313(.A (n_1213), .B (n_5712), .Y (n_1640));
NOR2X1 g59314(.A (n_1184), .B (n_1425), .Y (n_1639));
NOR2X1 g59315(.A (n_1183), .B (n_1425), .Y (n_1638));
NOR2X1 g59316(.A (n_1098), .B (n_5181), .Y (n_1637));
NOR2X1 g59317(.A (n_1180), .B (n_5712), .Y (n_1636));
NOR2X1 g59318(.A (n_1179), .B (n_5712), .Y (n_1635));
NOR2X1 g59319(.A (n_1177), .B (n_5712), .Y (n_1633));
AND2X1 g62702(.A (WX7202), .B (n_2378), .Y (n_1632));
NOR2X1 g59322(.A (n_1175), .B (n_1648), .Y (n_1631));
NOR2X1 g59323(.A (n_1256), .B (n_5712), .Y (n_1629));
NOR2X1 g59324(.A (n_1260), .B (n_1648), .Y (n_1628));
NOR2X1 g59325(.A (n_1056), .B (n_1648), .Y (n_1627));
NOR2X1 g59326(.A (n_1057), .B (n_1425), .Y (n_1626));
NOR2X1 g59327(.A (n_1173), .B (n_1425), .Y (n_1625));
NOR2X1 g59328(.A (n_1171), .B (n_5712), .Y (n_1624));
NOR2X1 g59329(.A (n_1017), .B (n_5181), .Y (n_1623));
NOR2X1 g59332(.A (n_1169), .B (n_1648), .Y (n_1622));
NOR2X1 g59333(.A (n_1126), .B (n_1648), .Y (n_1620));
NOR2X1 g59334(.A (n_1253), .B (n_1425), .Y (n_1619));
NOR2X1 g59335(.A (n_1259), .B (n_1425), .Y (n_1618));
NOR2X1 g59336(.A (n_1225), .B (n_1425), .Y (n_1617));
NOR2X1 g59337(.A (n_1105), .B (n_1425), .Y (n_1615));
NOR2X1 g59340(.A (n_1166), .B (n_5712), .Y (n_1614));
NOR2X1 g59341(.A (n_1252), .B (n_5712), .Y (n_1613));
NOR2X1 g59342(.A (n_1164), .B (n_5181), .Y (n_1612));
NOR2X1 g59343(.A (n_1240), .B (n_5181), .Y (n_1611));
NOR2X1 g59344(.A (n_1163), .B (n_5712), .Y (n_1609));
NOR2X1 g59345(.A (n_1162), .B (n_5712), .Y (n_1608));
NOR2X1 g59346(.A (n_1161), .B (n_5181), .Y (n_1607));
NOR2X1 g59348(.A (n_1095), .B (n_5181), .Y (n_1606));
NOR2X1 g59349(.A (n_1262), .B (n_5181), .Y (n_1605));
NOR2X1 g59350(.A (n_1160), .B (n_1425), .Y (n_1604));
NOR2X1 g59351(.A (n_1024), .B (n_1425), .Y (n_1603));
NOR2X1 g59354(.A (n_1157), .B (n_1425), .Y (n_1601));
NOR2X1 g59355(.A (n_1156), .B (n_1425), .Y (n_1600));
NOR2X1 g59358(.A (n_1037), .B (n_1648), .Y (n_1599));
NOR2X1 g59359(.A (n_1258), .B (n_5712), .Y (n_1598));
NOR2X1 g59360(.A (n_1153), .B (n_5712), .Y (n_1597));
NOR2X1 g59361(.A (n_1025), .B (n_5712), .Y (n_1595));
NOR2X1 g59362(.A (n_1151), .B (n_1648), .Y (n_1594));
NOR2X1 g59363(.A (n_1215), .B (n_1648), .Y (n_1593));
NOR2X1 g59364(.A (n_1243), .B (n_5712), .Y (n_1592));
NOR2X1 g59366(.A (n_1146), .B (n_1648), .Y (n_1591));
NOR2X1 g59368(.A (n_1018), .B (n_5181), .Y (n_1590));
NOR2X1 g59369(.A (n_1144), .B (n_5181), .Y (n_1588));
NOR2X1 g59370(.A (n_1214), .B (n_5712), .Y (n_1587));
NOR2X1 g59371(.A (n_1143), .B (n_5712), .Y (n_1585));
NOR2X1 g59372(.A (n_1036), .B (n_5181), .Y (n_1584));
NOR2X1 g59373(.A (n_1034), .B (n_5181), .Y (n_1583));
NOR2X1 g59374(.A (n_1139), .B (n_1648), .Y (n_1582));
NOR2X1 g59375(.A (n_1138), .B (n_1648), .Y (n_1581));
NOR2X1 g59377(.A (n_1137), .B (n_5712), .Y (n_1580));
NOR2X1 g59380(.A (n_1134), .B (n_1648), .Y (n_1579));
NOR2X1 g59381(.A (n_1212), .B (n_1425), .Y (n_1577));
NOR2X1 g59382(.A (n_1117), .B (n_5712), .Y (n_1576));
NOR2X1 g59383(.A (n_1046), .B (n_5181), .Y (n_1575));
NOR2X1 g59384(.A (n_1140), .B (n_1648), .Y (n_1574));
NOR2X1 g59385(.A (n_1255), .B (n_1648), .Y (n_1573));
NOR2X1 g59387(.A (n_1127), .B (n_1425), .Y (n_1572));
NOR2X1 g59388(.A (n_1053), .B (n_5712), .Y (n_1571));
NOR2X1 g59389(.A (n_1261), .B (n_5712), .Y (n_1570));
NOR2X1 g59392(.A (n_1061), .B (n_5712), .Y (n_1568));
NOR2X1 g59393(.A (n_1125), .B (n_5712), .Y (n_1567));
AND2X1 g62226(.A (WX4592), .B (n_2383), .Y (n_1566));
NOR2X1 g59395(.A (n_1122), .B (n_5712), .Y (n_1565));
NOR2X1 g59398(.A (n_1220), .B (n_1425), .Y (n_1564));
NOR2X1 g59399(.A (n_1219), .B (n_1425), .Y (n_1563));
NOR2X1 g59400(.A (n_1152), .B (n_5712), .Y (n_1561));
NOR2X1 g59401(.A (n_1249), .B (n_5712), .Y (n_1560));
NOR2X1 g59402(.A (n_1112), .B (n_1425), .Y (n_1559));
NOR2X1 g59403(.A (n_1211), .B (n_1425), .Y (n_1558));
NOR2X1 g59404(.A (n_1241), .B (n_5712), .Y (n_1557));
NOR2X1 g59406(.A (n_1107), .B (n_5712), .Y (n_1555));
NOR2X1 g59407(.A (n_1040), .B (n_5712), .Y (n_1554));
NOR2X1 g59410(.A (n_1039), .B (n_5181), .Y (n_1553));
NOR2X1 g59411(.A (n_1103), .B (n_5181), .Y (n_1552));
NOR2X1 g59417(.A (n_1096), .B (n_5181), .Y (n_1551));
NOR2X1 g59418(.A (n_1021), .B (n_5712), .Y (n_1550));
NOR2X1 g59419(.A (n_1246), .B (n_5712), .Y (n_1548));
NOR2X1 g59420(.A (n_1092), .B (n_5712), .Y (n_1547));
NOR2X1 g59421(.A (n_1063), .B (n_5181), .Y (n_1546));
NOR2X1 g59423(.A (n_1090), .B (n_1648), .Y (n_1545));
NOR2X1 g59424(.A (n_1089), .B (n_5712), .Y (n_1544));
NOR2X1 g59425(.A (n_1050), .B (n_5712), .Y (n_1542));
NOR2X1 g59426(.A (n_1088), .B (n_5712), .Y (n_1541));
NOR2X1 g59427(.A (n_1165), .B (n_5181), .Y (n_1540));
NOR2X1 g59428(.A (n_1087), .B (n_1425), .Y (n_1539));
NOR2X1 g59429(.A (n_1189), .B (n_1425), .Y (n_1537));
NOR2X1 g59432(.A (n_1085), .B (n_1648), .Y (n_1536));
NOR2X1 g59433(.A (n_1013), .B (n_1425), .Y (n_1535));
NOR2X1 g59438(.A (n_1041), .B (n_5181), .Y (n_1534));
NOR2X1 g59439(.A (n_1081), .B (n_5181), .Y (n_1533));
NOR2X1 g59440(.A (n_1174), .B (n_1648), .Y (n_1531));
NOR2X1 g59441(.A (n_1224), .B (n_5181), .Y (n_1530));
NOR2X1 g59442(.A (n_1052), .B (n_5181), .Y (n_1529));
NOR2X1 g59443(.A (n_1080), .B (n_5181), .Y (n_1528));
NOR2X1 g59444(.A (n_1028), .B (n_5712), .Y (n_1527));
AND2X1 g61735(.A (WX9556), .B (n_2246), .Y (n_1526));
NOR2X1 g59445(.A (n_1078), .B (n_1648), .Y (n_1525));
NOR2X1 g59446(.A (n_1223), .B (n_1648), .Y (n_1524));
NOR2X1 g59454(.A (n_1071), .B (n_1648), .Y (n_1523));
NOR2X1 g59455(.A (n_1236), .B (n_1648), .Y (n_1522));
NOR2X1 g59456(.A (n_1070), .B (n_5181), .Y (n_1521));
NOR2X1 g59457(.A (n_1016), .B (n_5181), .Y (n_1519));
NOR2X1 g59458(.A (n_1069), .B (n_5712), .Y (n_1518));
NOR2X1 g59459(.A (n_1232), .B (n_5712), .Y (n_1517));
NOR2X1 g59461(.A (n_1067), .B (n_1648), .Y (n_1516));
NOR2X1 g59462(.A (n_1124), .B (n_5712), .Y (n_1515));
NOR2X1 g59463(.A (n_1197), .B (n_1648), .Y (n_1514));
NOR2X1 g59471(.A (n_1198), .B (n_5181), .Y (n_1513));
NOR2X1 g59472(.A (n_1031), .B (n_5181), .Y (n_1512));
NOR2X1 g59473(.A (n_1110), .B (n_1425), .Y (n_1511));
NOR2X1 g59474(.A (n_1206), .B (n_1425), .Y (n_1510));
NOR2X1 g59483(.A (n_1100), .B (n_1425), .Y (n_1509));
NOR2X1 g59484(.A (n_1133), .B (n_5712), .Y (n_1508));
NOR2X1 g59485(.A (n_1129), .B (n_5712), .Y (n_1507));
NOR2X1 g59486(.A (n_1141), .B (n_5712), .Y (n_1506));
NOR2X1 g59487(.A (n_1200), .B (n_5712), .Y (n_1504));
NOR2X1 g59489(.A (n_1178), .B (n_5712), .Y (n_1503));
NOR2X1 g59490(.A (n_1093), .B (n_5712), .Y (n_1502));
NOR2X1 g59492(.A (n_1115), .B (n_5712), .Y (n_1500));
NOR2X1 g59493(.A (n_1012), .B (n_5712), .Y (n_1499));
NOR2X1 g59495(.A (n_1130), .B (n_5712), .Y (n_1498));
NOR2X1 g59496(.A (n_1248), .B (n_1648), .Y (n_1497));
NOR2X1 g59497(.A (n_1159), .B (n_5712), .Y (n_1496));
AND2X1 g59498(.A (WX11053), .B (n_2325), .Y (n_1495));
AND2X1 g62676(.A (WX11129), .B (n_2346), .Y (n_1494));
AND2X1 g59512(.A (WX2002), .B (n_2346), .Y (n_1493));
AND2X1 g62671(.A (WX3359), .B (n_2333), .Y (n_1492));
AND2X1 g61705(.A (WX7198), .B (n_2311), .Y (n_1491));
AND2X1 g62663(.A (WX11155), .B (n_2251), .Y (n_1490));
AND2X1 g62181(.A (WX7262), .B (n_2223), .Y (n_1489));
AND2X1 g62548(.A (WX9794), .B (n_2383), .Y (n_1488));
AND2X1 g62659(.A (WX8265), .B (n_2198), .Y (n_1487));
AND2X1 g62657(.A (WX9848), .B (n_2272), .Y (n_1486));
AND2X1 g61684(.A (WX8533), .B (n_2325), .Y (n_1485));
AND2X1 g62638(.A (WX9874), .B (n_2383), .Y (n_1484));
AND2X1 g61663(.A (WX11045), .B (n_2311), .Y (n_1483));
AND2X1 g62636(.A (WX11069), .B (n_2371), .Y (n_1482));
AND2X1 g61655(.A (WX11041), .B (n_2527), .Y (n_1481));
AND2X1 g61650(.A (WX9786), .B (n_2383), .Y (n_1480));
AND2X1 g61640(.A (WX2072), .B (n_2325), .Y (n_1479));
AND2X1 g62632(.A (WX4648), .B (n_2227), .Y (n_1478));
AND2X1 g62625(.A (WX5817), .B (n_2527), .Y (n_1477));
AND2X1 g62622(.A (WX5837), .B (n_2400), .Y (n_1476));
AOI21X1 g57873(.A0 (_2107_), .A1 (WX837), .B0 (n_1038), .Y (n_1473));
AND2X1 g61631(.A (WX7284), .B (n_2527), .Y (n_1472));
AND2X1 g62554(.A (WX5821), .B (n_2227), .Y (n_1471));
AND2X1 g61607(.A (WX11167), .B (n_2227), .Y (n_1470));
INVX4 g63523(.A (n_2227), .Y (n_3690));
NOR2X1 g61584(.A (n_5181), .B (n_35), .Y (n_1465));
NOR2X1 g56990(.A (WX5659), .B (n_1648), .Y (n_1464));
NOR2X1 g62598(.A (n_1425), .B (n_2), .Y (n_1462));
NOR2X1 g62595(.A (n_5181), .B (n_970), .Y (n_1461));
NAND2X1 g60725(.A (n_597), .B (n_596), .Y (n_2511));
NAND2X1 g60796(.A (n_568), .B (n_590), .Y (n_2498));
NAND2X1 g60808(.A (n_582), .B (n_583), .Y (n_2494));
NOR2X1 g57058(.A (WX6952), .B (n_1648), .Y (n_1459));
NOR2X1 g62566(.A (n_5181), .B (n_112), .Y (n_1458));
NOR2X1 g55933(.A (n_1425), .B (n_3685), .Y (n_1456));
NAND2X1 g60903(.A (n_578), .B (n_576), .Y (n_2472));
NAND2X1 g60951(.A (n_548), .B (n_771), .Y (n_2468));
NOR2X1 g57096(.A (WX8245), .B (n_1648), .Y (n_1454));
NAND2X1 g60965(.A (n_570), .B (n_569), .Y (n_2466));
NAND2X1 g61011(.A (n_564), .B (n_563), .Y (n_2458));
NAND2X1 g61058(.A (n_593), .B (n_573), .Y (n_2453));
NAND2X1 g61092(.A (n_559), .B (n_547), .Y (n_2443));
NAND2X1 g61152(.A (n_557), .B (n_555), .Y (n_2437));
NOR2X1 g57161(.A (WX9538), .B (n_1425), .Y (n_1453));
NAND2X1 g61220(.A (n_545), .B (n_544), .Y (n_2422));
NOR2X1 g61559(.A (n_1451), .B (n_1425), .Y (n_1452));
NOR2X1 g61565(.A (n_1449), .B (n_5181), .Y (n_1450));
NOR2X1 g61579(.A (n_5181), .B (n_69), .Y (n_1448));
NOR2X1 g61588(.A (n_5181), .B (n_87), .Y (n_1447));
NOR2X1 g61605(.A (n_1425), .B (n_81), .Y (n_1446));
NOR2X1 g61608(.A (n_1425), .B (n_4), .Y (n_1444));
NOR2X1 g61612(.A (n_1442), .B (n_1425), .Y (n_1443));
NOR2X1 g61624(.A (n_1425), .B (n_951), .Y (n_1441));
NOR2X1 g61633(.A (n_1425), .B (n_1006), .Y (n_1440));
NOR2X1 g61636(.A (n_1437), .B (n_1425), .Y (n_1438));
NOR2X1 g61662(.A (n_5181), .B (n_67), .Y (n_1436));
NOR2X1 g61683(.A (n_1425), .B (n_119), .Y (n_1435));
NOR2X1 g61696(.A (n_5181), .B (n_1001), .Y (n_1433));
NOR2X1 g61736(.A (n_1431), .B (n_5712), .Y (n_1432));
NOR2X1 g61740(.A (n_1429), .B (n_5712), .Y (n_1430));
NOR2X1 g61748(.A (n_1427), .B (n_5181), .Y (n_1428));
NOR2X1 g61758(.A (n_1425), .B (n_12), .Y (n_1426));
NOR2X1 g58602(.A (n_5181), .B (n_0), .Y (n_1424));
NOR2X1 g61764(.A (n_1425), .B (n_940), .Y (n_1423));
NOR2X1 g61767(.A (n_1421), .B (n_1425), .Y (n_1422));
NOR2X1 g61776(.A (n_1419), .B (n_1425), .Y (n_1420));
NOR2X1 g61780(.A (n_1425), .B (n_958), .Y (n_1418));
NOR2X1 g61786(.A (n_1425), .B (n_56), .Y (n_1417));
NOR2X1 g61787(.A (n_1425), .B (n_109), .Y (n_1415));
NOR2X1 g61798(.A (n_5181), .B (n_52), .Y (n_1414));
NOR2X1 g61813(.A (n_1412), .B (n_1648), .Y (n_1413));
NOR2X1 g61818(.A (n_5181), .B (n_32), .Y (n_1411));
NOR2X1 g61822(.A (n_1425), .B (n_96), .Y (n_1410));
NOR2X1 g61844(.A (n_1425), .B (n_985), .Y (n_1409));
NOR2X1 g61853(.A (n_5181), .B (n_14), .Y (n_1407));
NOR2X1 g61875(.A (n_1425), .B (n_19), .Y (n_1405));
NOR2X1 g61878(.A (n_1425), .B (n_981), .Y (n_1404));
NOR2X1 g61880(.A (n_1425), .B (n_913), .Y (n_1403));
NOR2X1 g61895(.A (n_1425), .B (n_975), .Y (n_1402));
NOR2X1 g61924(.A (n_1425), .B (n_101), .Y (n_1400));
NOR2X1 g61927(.A (n_5181), .B (n_28), .Y (n_1399));
NOR2X1 g61928(.A (n_5181), .B (n_118), .Y (n_1398));
NOR2X1 g61930(.A (n_5181), .B (n_995), .Y (n_1396));
NOR2X1 g61945(.A (n_5181), .B (n_117), .Y (n_1395));
NOR2X1 g61951(.A (n_1425), .B (n_990), .Y (n_1393));
NOR2X1 g61974(.A (n_5181), .B (n_16), .Y (n_1391));
NOR2X1 g61984(.A (n_5181), .B (n_1004), .Y (n_1389));
NOR2X1 g61989(.A (n_1425), .B (n_46), .Y (n_1388));
NOR2X1 g62005(.A (n_5181), .B (n_41), .Y (n_1387));
NOR2X1 g62007(.A (n_1425), .B (n_18), .Y (n_1386));
NOR2X1 g62008(.A (n_5181), .B (n_51), .Y (n_1385));
NOR2X1 g62042(.A (n_5181), .B (n_130), .Y (n_1384));
NOR2X1 g62045(.A (n_5181), .B (n_929), .Y (n_1382));
NOR2X1 g62046(.A (n_5181), .B (n_68), .Y (n_1381));
NOR2X1 g62051(.A (n_5181), .B (n_3), .Y (n_1380));
NOR2X1 g62073(.A (n_1425), .B (n_79), .Y (n_1379));
NOR2X1 g62085(.A (n_1425), .B (n_105), .Y (n_1378));
NOR2X1 g62102(.A (n_1425), .B (n_111), .Y (n_1377));
NOR2X1 g62110(.A (n_1374), .B (n_1648), .Y (n_1375));
NOR2X1 g62153(.A (n_1425), .B (n_964), .Y (n_1373));
NOR2X1 g62169(.A (n_1425), .B (n_948), .Y (n_1372));
NOR2X1 g62173(.A (n_1425), .B (n_24), .Y (n_1371));
NOR2X1 g62179(.A (n_1425), .B (n_70), .Y (n_1370));
NOR2X1 g62186(.A (n_1425), .B (n_73), .Y (n_1369));
NOR2X1 g62193(.A (n_1425), .B (n_938), .Y (n_1367));
NOR2X1 g62200(.A (n_5181), .B (n_38), .Y (n_1366));
NOR2X1 g62223(.A (n_1425), .B (n_905), .Y (n_1365));
NOR2X1 g62225(.A (n_5181), .B (n_987), .Y (n_1364));
NOR2X1 g62250(.A (n_1425), .B (n_129), .Y (n_1362));
NOR2X1 g62284(.A (n_1359), .B (n_1425), .Y (n_1360));
NOR2X1 g62307(.A (n_1357), .B (n_5181), .Y (n_1358));
NOR2X1 g62309(.A (n_1425), .B (n_43), .Y (n_1356));
NOR2X1 g62330(.A (n_1425), .B (n_71), .Y (n_1355));
NOR2X1 g62338(.A (n_1425), .B (n_83), .Y (n_1354));
NOR2X1 g62342(.A (n_5181), .B (n_21), .Y (n_1353));
NOR2X1 g62353(.A (n_1425), .B (n_956), .Y (n_1352));
NOR2X1 g62356(.A (n_1350), .B (n_1425), .Y (n_1351));
NOR2X1 g62359(.A (n_1348), .B (n_1425), .Y (n_1349));
NOR2X1 g62365(.A (n_1425), .B (n_89), .Y (n_1347));
NOR2X1 g62366(.A (n_1345), .B (n_5181), .Y (n_1346));
NOR2X1 g62368(.A (n_1425), .B (n_58), .Y (n_1344));
NOR2X1 g62371(.A (n_1341), .B (n_5181), .Y (n_1342));
NOR2X1 g62469(.A (n_1339), .B (n_5181), .Y (n_1340));
NOR2X1 g62473(.A (n_1337), .B (n_1425), .Y (n_1338));
NOR2X1 g62474(.A (n_1335), .B (n_1425), .Y (n_1336));
NOR2X1 g62478(.A (n_5181), .B (n_104), .Y (n_1334));
NOR2X1 g62488(.A (n_1425), .B (n_98), .Y (n_1333));
NOR2X1 g62493(.A (n_5181), .B (n_992), .Y (n_1332));
NOR2X1 g62498(.A (n_1425), .B (n_932), .Y (n_1330));
NOR2X1 g62537(.A (n_1328), .B (n_1425), .Y (n_1329));
NOR2X1 g62543(.A (n_5181), .B (n_27), .Y (n_1327));
NOR2X1 g62584(.A (n_5181), .B (n_997), .Y (n_1326));
NOR2X1 g62604(.A (n_5181), .B (n_48), .Y (n_1325));
NOR2X1 g62607(.A (n_1323), .B (n_1425), .Y (n_1324));
NOR2X1 g62635(.A (n_1425), .B (n_63), .Y (n_1322));
NOR2X1 g62644(.A (n_1320), .B (n_1648), .Y (n_1321));
NOR2X1 g62655(.A (n_1318), .B (n_5181), .Y (n_1319));
NOR2X1 g62678(.A (n_5181), .B (n_973), .Y (n_1317));
NOR2X1 g62741(.A (n_1315), .B (n_5712), .Y (n_1316));
NOR2X1 g62742(.A (n_5181), .B (n_113), .Y (n_1314));
NOR2X1 g62744(.A (n_5181), .B (n_36), .Y (n_1313));
NOR2X1 g62755(.A (n_1425), .B (n_20), .Y (n_1312));
NOR2X1 g62756(.A (n_1425), .B (n_106), .Y (n_1311));
NOR2X1 g62761(.A (n_1309), .B (n_1425), .Y (n_1310));
NOR2X1 g62768(.A (n_1425), .B (n_44), .Y (n_1308));
NOR2X1 g62746(.A (n_1425), .B (n_100), .Y (n_1307));
NOR2X1 g62745(.A (n_5181), .B (n_65), .Y (n_1306));
INVX4 g63039(.A (n_1460), .Y (n_3058));
INVX4 g63043(.A (n_1305), .Y (n_3106));
INVX1 g63227(.A (n_1278), .Y (n_2993));
INVX1 g63230(.A (n_1278), .Y (n_3044));
INVX1 g63231(.A (n_1278), .Y (n_2996));
INVX1 g63233(.A (n_1278), .Y (n_2976));
INVX4 g63503(.A (n_2378), .Y (n_2605));
INVX8 g63530(.A (n_2227), .Y (n_2851));
INVX8 g63543(.A (n_1297), .Y (n_3188));
INVX8 g63554(.A (n_2227), .Y (n_2620));
INVX4 g63584(.A (n_6428), .Y (n_2938));
INVX8 g63599(.A (n_1294), .Y (n_3072));
NOR2X1 g62686(.A (n_5181), .B (n_962), .Y (n_1291));
NOR2X1 g59500(.A (n_1425), .B (n_95), .Y (n_1290));
NOR2X1 g62651(.A (n_1288), .B (n_5712), .Y (n_1289));
NOR2X1 g62650(.A (n_1286), .B (n_1648), .Y (n_1287));
NOR2X1 g62641(.A (n_1284), .B (n_5712), .Y (n_1285));
NOR2X1 g61688(.A (n_1282), .B (n_5712), .Y (n_1283));
INVX4 g63665(.A (n_1281), .Y (n_2945));
INVX4 g63659(.A (n_3120), .Y (n_3086));
NOR2X1 g62553(.A (n_5181), .B (n_49), .Y (n_1280));
NAND2X1 g61084(.A (n_551), .B (n_566), .Y (n_2446));
NOR2X1 g56884(.A (WX3073), .B (n_1648), .Y (n_1279));
INVX1 g63232(.A (n_1278), .Y (n_3004));
INVX1 g63228(.A (n_1278), .Y (n_3056));
INVX1 g63226(.A (n_1278), .Y (n_3105));
INVX1 g63225(.A (n_1278), .Y (n_3103));
NOR2X1 g61621(.A (n_1425), .B (n_953), .Y (n_1277));
INVX4 g63591(.A (n_1276), .Y (n_3041));
NOR2X1 g61609(.A (n_1425), .B (n_944), .Y (n_1275));
NOR2X1 g61593(.A (_2078_), .B (WX895), .Y (n_1272));
AOI21X1 g60389(.A0 (WX9936), .A1 (_2307_), .B0 (n_412), .Y (n_1268));
AOI21X1 g60390(.A0 (WX9930), .A1 (_2310_), .B0 (n_302), .Y (n_1267));
AOI21X1 g60391(.A0 (WX7302), .A1 (_2267_), .B0 (n_419), .Y (n_1265));
AOI21X1 g60392(.A0 (WX11213), .A1 (_2347_), .B0 (n_285), .Y (n_1264));
AOI21X1 g60393(.A0 (WX6041), .A1 (_2219_), .B0 (n_324), .Y (n_1263));
BUFX3 g63475(.A (n_2298), .Y (n_2216));
AOI21X1 g60394(.A0 (WX4732), .A1 (_2195_), .B0 (n_332), .Y (n_1262));
AOI21X1 g60395(.A0 (WX6069), .A1 (_2205_), .B0 (n_328), .Y (n_1261));
AOI21X1 g60396(.A0 (WX3435), .A1 (_2165_), .B0 (n_427), .Y (n_1260));
AOI21X1 g60397(.A0 (WX4766), .A1 (_2178_), .B0 (n_145), .Y (n_1259));
AOI21X1 g60398(.A0 (WX6059), .A1 (_2210_), .B0 (n_200), .Y (n_1258));
AOI21X1 g60400(.A0 (WX4746), .A1 (_2204_), .B0 (n_422), .Y (n_1257));
BUFX3 g63477(.A (n_2298), .Y (n_2188));
AOI21X1 g60401(.A0 (WX3437), .A1 (_2164_), .B0 (n_232), .Y (n_1256));
AOI21X1 g60403(.A0 (WX7326), .A1 (_2255_), .B0 (n_148), .Y (n_1255));
AOI21X1 g60404(.A0 (WX2184), .A1 (_2140_), .B0 (n_469), .Y (n_1254));
AOI21X1 g60406(.A0 (WX4768), .A1 (_2177_), .B0 (n_198), .Y (n_1253));
AOI21X1 g60407(.A0 (WX4750), .A1 (_2186_), .B0 (n_254), .Y (n_1252));
AOI21X1 g60408(.A0 (WX3469), .A1 (_2148_), .B0 (n_377), .Y (n_1251));
AOI21X1 g60409(.A0 (WX2138), .A1 (_2135_), .B0 (n_136), .Y (n_1250));
AOI21X1 g60410(.A0 (WX8631), .A1 (_2281_), .B0 (n_181), .Y (n_1249));
AOI21X1 g60411(.A0 (WX8643), .A1 (_2275_), .B0 (n_415), .Y (n_1248));
AOI21X1 g60412(.A0 (WX11203), .A1 (_2352_), .B0 (n_151), .Y (n_1247));
AOI21X1 g60413(.A0 (WX9922), .A1 (_2314_), .B0 (n_428), .Y (n_1246));
AOI21X1 g60414(.A0 (WX8605), .A1 (_2294_), .B0 (n_317), .Y (n_1245));
AOI21X1 g60415(.A0 (WX9946), .A1 (_2302_), .B0 (n_407), .Y (n_1244));
AOI21X1 g60416(.A0 (WX6047), .A1 (_2216_), .B0 (n_453), .Y (n_1243));
AOI21X1 g60417(.A0 (WX7310), .A1 (_2263_), .B0 (n_433), .Y (n_1242));
AOI21X1 g60418(.A0 (WX8621), .A1 (_2286_), .B0 (n_461), .Y (n_1241));
AOI21X1 g60419(.A0 (WX4744), .A1 (_2189_), .B0 (n_199), .Y (n_1240));
AOI21X1 g60420(.A0 (WX7340), .A1 (_2248_), .B0 (n_157), .Y (n_1239));
INVX4 g63466(.A (n_2298), .Y (n_2849));
AOI21X1 g60421(.A0 (WX7342), .A1 (_2268_), .B0 (n_150), .Y (n_1237));
AOI21X1 g60422(.A0 (WX11195), .A1 (_2356_), .B0 (n_349), .Y (n_1236));
AOI21X1 g60423(.A0 (WX4728), .A1 (_2197_), .B0 (n_479), .Y (n_1235));
AOI21X1 g60424(.A0 (WX4754), .A1 (_2184_), .B0 (n_192), .Y (n_1234));
AOI21X1 g60425(.A0 (WX3425), .A1 (_2170_), .B0 (n_176), .Y (n_1233));
AOI21X1 g60426(.A0 (WX11187), .A1 (_2360_), .B0 (n_405), .Y (n_1232));
AOI21X1 g60427(.A0 (WX2160), .A1 (_2140_), .B0 (n_306), .Y (n_1231));
AOI21X1 g60429(.A0 (WX11241), .A1 (_2333_), .B0 (n_153), .Y (n_1230));
AOI21X1 g60430(.A0 (WX6061), .A1 (_2209_), .B0 (n_178), .Y (n_1229));
AOI21X1 g60432(.A0 (WX8609), .A1 (_2292_), .B0 (n_410), .Y (n_1228));
AOI21X1 g60433(.A0 (WX3441), .A1 (_2162_), .B0 (n_341), .Y (n_1227));
AOI21X1 g60434(.A0 (WX7354), .A1 (_2241_), .B0 (n_316), .Y (n_1226));
AOI21X1 g60435(.A0 (WX4764), .A1 (_2179_), .B0 (n_142), .Y (n_1225));
AOI21X1 g60436(.A0 (WX11229), .A1 (_2339_), .B0 (n_386), .Y (n_1224));
AOI21X1 g60437(.A0 (WX11217), .A1 (_2345_), .B0 (n_194), .Y (n_1223));
AOI21X1 g60438(.A0 (WX8651), .A1 (_2271_), .B0 (n_382), .Y (n_1222));
AOI21X1 g60439(.A0 (WX2170), .A1 (_2140_), .B0 (n_228), .Y (n_1221));
AOI21X1 g60441(.A0 (WX8645), .A1 (_2274_), .B0 (n_440), .Y (n_1220));
AOI21X1 g60442(.A0 (WX8641), .A1 (_2276_), .B0 (n_213), .Y (n_1219));
AOI21X1 g60443(.A0 (WX7328), .A1 (_2254_), .B0 (n_468), .Y (n_1218));
AOI21X1 g60444(.A0 (WX8607), .A1 (_2293_), .B0 (n_362), .Y (n_1217));
AOI21X1 g60445(.A0 (WX7362), .A1 (_2237_), .B0 (n_227), .Y (n_1216));
AOI21X1 g60446(.A0 (WX6051), .A1 (_2214_), .B0 (n_172), .Y (n_1215));
AOI21X1 g60447(.A0 (WX6023), .A1 (_2228_), .B0 (n_295), .Y (n_1214));
AOI21X1 g60448(.A0 (WX3465), .A1 (_2150_), .B0 (n_374), .Y (n_1213));
AOI21X1 g60450(.A0 (WX6025), .A1 (_2227_), .B0 (n_408), .Y (n_1212));
AOI21X1 g60454(.A0 (WX8627), .A1 (_2283_), .B0 (n_318), .Y (n_1211));
AOI21X1 g60467(.A0 (WX4770), .A1 (_2204_), .B0 (n_169), .Y (n_1210));
AOI21X1 g60468(.A0 (WX2190), .A1 (_2109_), .B0 (n_376), .Y (n_1209));
AOI21X1 g60469(.A0 (WX2186), .A1 (_2111_), .B0 (n_291), .Y (n_1208));
AOI21X1 g60470(.A0 (WX2180), .A1 (_2114_), .B0 (n_399), .Y (n_1207));
AOI21X1 g60471(.A0 (WX2176), .A1 (_2116_), .B0 (n_385), .Y (n_1206));
AOI21X1 g60472(.A0 (WX2172), .A1 (_2118_), .B0 (n_185), .Y (n_1205));
AOI21X1 g60473(.A0 (WX2166), .A1 (_2121_), .B0 (n_326), .Y (n_1204));
AOI21X1 g60474(.A0 (WX2162), .A1 (_2123_), .B0 (n_209), .Y (n_1203));
AOI21X1 g60475(.A0 (WX2158), .A1 (_2125_), .B0 (n_235), .Y (n_1202));
AOI21X1 g60476(.A0 (WX2156), .A1 (_2126_), .B0 (n_365), .Y (n_1201));
AOI21X1 g60477(.A0 (WX2152), .A1 (_2128_), .B0 (n_325), .Y (n_1200));
AOI21X1 g60478(.A0 (WX2144), .A1 (_2132_), .B0 (n_205), .Y (n_1199));
AOI21X1 g60479(.A0 (WX2140), .A1 (_2134_), .B0 (n_304), .Y (n_1198));
AOI21X1 g60480(.A0 (WX2136), .A1 (_2136_), .B0 (n_373), .Y (n_1197));
AOI21X1 g60481(.A0 (WX2134), .A1 (_2137_), .B0 (n_247), .Y (n_1196));
AOI21X1 g60482(.A0 (WX2132), .A1 (_2138_), .B0 (n_229), .Y (n_1195));
AOI21X1 g60483(.A0 (WX3485), .A1 (_2172_), .B0 (n_171), .Y (n_1194));
AOI21X1 g60484(.A0 (WX3483), .A1 (_2141_), .B0 (n_402), .Y (n_1193));
AOI21X1 g60485(.A0 (WX3481), .A1 (_2142_), .B0 (n_401), .Y (n_1192));
AOI21X1 g60486(.A0 (WX3479), .A1 (_2143_), .B0 (n_314), .Y (n_1191));
AOI21X1 g60487(.A0 (WX3475), .A1 (_2145_), .B0 (n_464), .Y (n_1190));
AOI21X1 g60488(.A0 (WX9900), .A1 (_2325_), .B0 (n_135), .Y (n_1189));
AOI21X1 g60489(.A0 (WX3473), .A1 (_2146_), .B0 (n_489), .Y (n_1188));
AOI21X1 g60490(.A0 (WX3471), .A1 (_2147_), .B0 (n_313), .Y (n_1187));
AOI21X1 g60491(.A0 (WX3463), .A1 (_2172_), .B0 (n_457), .Y (n_1186));
AOI21X1 g60492(.A0 (WX3461), .A1 (_2152_), .B0 (n_423), .Y (n_1185));
AOI21X1 g60493(.A0 (WX3459), .A1 (_2153_), .B0 (n_488), .Y (n_1184));
AOI21X1 g60494(.A0 (WX3457), .A1 (_2154_), .B0 (n_414), .Y (n_1183));
AOI21X1 g60495(.A0 (WX9940), .A1 (_2305_), .B0 (n_131), .Y (n_1182));
AOI21X1 g60496(.A0 (WX3453), .A1 (_2172_), .B0 (n_356), .Y (n_1181));
AOI21X1 g60497(.A0 (WX3451), .A1 (_2157_), .B0 (n_206), .Y (n_1180));
AOI21X1 g60498(.A0 (WX3449), .A1 (_2158_), .B0 (n_396), .Y (n_1179));
AOI21X1 g60499(.A0 (WX3447), .A1 (_2159_), .B0 (n_170), .Y (n_1178));
AOI21X1 g60500(.A0 (WX3445), .A1 (_2160_), .B0 (n_389), .Y (n_1177));
AOI21X1 g60501(.A0 (WX3443), .A1 (_2161_), .B0 (n_299), .Y (n_1176));
AOI21X1 g60502(.A0 (WX3439), .A1 (_2163_), .B0 (n_395), .Y (n_1175));
AOI21X1 g60503(.A0 (WX11231), .A1 (_2338_), .B0 (n_257), .Y (n_1174));
AOI21X1 g60504(.A0 (WX3429), .A1 (_2168_), .B0 (n_460), .Y (n_1173));
AOI21X1 g60505(.A0 (WX3427), .A1 (_2169_), .B0 (n_387), .Y (n_1172));
AOI21X1 g60506(.A0 (WX3423), .A1 (_2171_), .B0 (n_394), .Y (n_1171));
AOI21X1 g60507(.A0 (WX4776), .A1 (_2173_), .B0 (n_184), .Y (n_1170));
AOI21X1 g60508(.A0 (WX4772), .A1 (_2175_), .B0 (n_391), .Y (n_1169));
AOI21X1 g60509(.A0 (WX4762), .A1 (_2180_), .B0 (n_141), .Y (n_1168));
AOI21X1 g60510(.A0 (WX4758), .A1 (_2182_), .B0 (n_163), .Y (n_1167));
AOI21X1 g60511(.A0 (WX4752), .A1 (_2185_), .B0 (n_322), .Y (n_1166));
AOI21X1 g60512(.A0 (WX9904), .A1 (_2323_), .B0 (n_329), .Y (n_1165));
AOI21X1 g60513(.A0 (WX4748), .A1 (_2187_), .B0 (n_154), .Y (n_1164));
AOI21X1 g60514(.A0 (WX4742), .A1 (_2190_), .B0 (n_189), .Y (n_1163));
AOI21X1 g60515(.A0 (WX4740), .A1 (_2191_), .B0 (n_179), .Y (n_1162));
AOI21X1 g60516(.A0 (WX4738), .A1 (_2192_), .B0 (n_173), .Y (n_1161));
AOI21X1 g60517(.A0 (WX4730), .A1 (_2196_), .B0 (n_353), .Y (n_1160));
AOI21X1 g60518(.A0 (WX4726), .A1 (_2198_), .B0 (n_357), .Y (n_1159));
AOI21X1 g60519(.A0 (WX4722), .A1 (_2200_), .B0 (n_331), .Y (n_1158));
AOI21X1 g60520(.A0 (WX4718), .A1 (_2202_), .B0 (n_162), .Y (n_1157));
AOI21X1 g60521(.A0 (WX4716), .A1 (_2203_), .B0 (n_300), .Y (n_1156));
AOI21X1 g60522(.A0 (WX6067), .A1 (_2206_), .B0 (n_315), .Y (n_1155));
AOI21X1 g60523(.A0 (WX6063), .A1 (_2236_), .B0 (n_212), .Y (n_1154));
AOI21X1 g60524(.A0 (WX6057), .A1 (_2211_), .B0 (n_406), .Y (n_1153));
AOI21X1 g60525(.A0 (WX8637), .A1 (_2278_), .B0 (n_366), .Y (n_1152));
AOI21X1 g60526(.A0 (WX6053), .A1 (_2213_), .B0 (n_397), .Y (n_1151));
AOI21X1 g60527(.A0 (WX6049), .A1 (_2236_), .B0 (n_307), .Y (n_1150));
AOI21X1 g60528(.A0 (WX6043), .A1 (_2218_), .B0 (n_470), .Y (n_1149));
AOI21X1 g60529(.A0 (WX6039), .A1 (_2236_), .B0 (n_347), .Y (n_1148));
AOI21X1 g60530(.A0 (WX6037), .A1 (_2221_), .B0 (n_301), .Y (n_1147));
AOI21X1 g60531(.A0 (WX6035), .A1 (_2222_), .B0 (n_392), .Y (n_1146));
AOI21X1 g60532(.A0 (WX6033), .A1 (_2223_), .B0 (n_164), .Y (n_1145));
AOI21X1 g60533(.A0 (WX6029), .A1 (_2225_), .B0 (n_372), .Y (n_1144));
AOI21X1 g60534(.A0 (WX6021), .A1 (_2229_), .B0 (n_156), .Y (n_1143));
AOI21X1 g60535(.A0 (WX6017), .A1 (_2231_), .B0 (n_418), .Y (n_1142));
AOI21X1 g60536(.A0 (WX6013), .A1 (_2233_), .B0 (n_133), .Y (n_1141));
AOI21X1 g60537(.A0 (WX7330), .A1 (_2253_), .B0 (n_256), .Y (n_1140));
AOI21X1 g60538(.A0 (WX6011), .A1 (_2234_), .B0 (n_339), .Y (n_1139));
AOI21X1 g60539(.A0 (WX6009), .A1 (_2235_), .B0 (n_166), .Y (n_1138));
AOI21X1 g60540(.A0 (WX7360), .A1 (_2238_), .B0 (n_177), .Y (n_1137));
AOI21X1 g60541(.A0 (WX7358), .A1 (_2239_), .B0 (n_211), .Y (n_1136));
AOI21X1 g60542(.A0 (WX7356), .A1 (_2268_), .B0 (n_180), .Y (n_1135));
AOI21X1 g60543(.A0 (WX7352), .A1 (_2242_), .B0 (n_231), .Y (n_1134));
AOI21X1 g60544(.A0 (WX7344), .A1 (_2246_), .B0 (n_350), .Y (n_1133));
AOI21X1 g60545(.A0 (WX11183), .A1 (_2362_), .B0 (n_409), .Y (n_1132));
AOI21X1 g60546(.A0 (WX7338), .A1 (_2249_), .B0 (n_384), .Y (n_1131));
AOI21X1 g60547(.A0 (WX7334), .A1 (_2251_), .B0 (n_167), .Y (n_1130));
AOI21X1 g60548(.A0 (WX7324), .A1 (_2256_), .B0 (n_230), .Y (n_1129));
AOI21X1 g60549(.A0 (WX7322), .A1 (_2257_), .B0 (n_416), .Y (n_1128));
AOI21X1 g60550(.A0 (WX7320), .A1 (_2258_), .B0 (n_233), .Y (n_1127));
AOI21X1 g60551(.A0 (WX7316), .A1 (_2260_), .B0 (n_195), .Y (n_1126));
AOI21X1 g60552(.A0 (WX7306), .A1 (_2265_), .B0 (n_380), .Y (n_1125));
AOI21X1 g60553(.A0 (WX7304), .A1 (_2266_), .B0 (n_334), .Y (n_1124));
AOI21X1 g60554(.A0 (WX8657), .A1 (_2300_), .B0 (n_447), .Y (n_1123));
AOI21X1 g60555(.A0 (WX8655), .A1 (_2269_), .B0 (n_289), .Y (n_1122));
AOI21X1 g60556(.A0 (WX8653), .A1 (_2270_), .B0 (n_146), .Y (n_1121));
AOI21X1 g60557(.A0 (WX8649), .A1 (_2300_), .B0 (n_369), .Y (n_1120));
AOI21X1 g60558(.A0 (WX4720), .A1 (_2201_), .B0 (n_465), .Y (n_1119));
AOI21X1 g60559(.A0 (WX8601), .A1 (_2296_), .B0 (n_147), .Y (n_1118));
AOI21X1 g60560(.A0 (WX8647), .A1 (_2273_), .B0 (n_417), .Y (n_1117));
AOI21X1 g60561(.A0 (WX7332), .A1 (_2268_), .B0 (n_393), .Y (n_1116));
AOI21X1 g60562(.A0 (WX8639), .A1 (_2277_), .B0 (n_288), .Y (n_1115));
AOI21X1 g60563(.A0 (WX8635), .A1 (_2300_), .B0 (n_426), .Y (n_1114));
AOI21X1 g60564(.A0 (WX8633), .A1 (_2280_), .B0 (n_225), .Y (n_1113));
AOI21X1 g60565(.A0 (WX8629), .A1 (_2282_), .B0 (n_187), .Y (n_1112));
AOI21X1 g60566(.A0 (WX8625), .A1 (_2300_), .B0 (n_188), .Y (n_1111));
AOI21X1 g60567(.A0 (WX8623), .A1 (_2285_), .B0 (n_358), .Y (n_1110));
AOI21X1 g60568(.A0 (WX8619), .A1 (_2287_), .B0 (n_197), .Y (n_1109));
AOI21X1 g60569(.A0 (WX8617), .A1 (_2288_), .B0 (n_298), .Y (n_1108));
AOI21X1 g60570(.A0 (WX8615), .A1 (_2289_), .B0 (n_226), .Y (n_1107));
AOI21X1 g60571(.A0 (WX8611), .A1 (_2291_), .B0 (n_403), .Y (n_1106));
AOI21X1 g60572(.A0 (WX4760), .A1 (_2181_), .B0 (n_258), .Y (n_1105));
AOI21X1 g60573(.A0 (WX8599), .A1 (_2297_), .B0 (n_293), .Y (n_1104));
AOI21X1 g60574(.A0 (WX8595), .A1 (_2299_), .B0 (n_330), .Y (n_1103));
AOI21X1 g60575(.A0 (WX9950), .A1 (_2332_), .B0 (n_241), .Y (n_1102));
AOI21X1 g60576(.A0 (WX9948), .A1 (_2301_), .B0 (n_333), .Y (n_1101));
AOI21X1 g60577(.A0 (WX9944), .A1 (_2303_), .B0 (n_207), .Y (n_1100));
AOI21X1 g60578(.A0 (WX9938), .A1 (_2306_), .B0 (n_375), .Y (n_1099));
AOI21X1 g60579(.A0 (WX3455), .A1 (_2155_), .B0 (n_175), .Y (n_1098));
AOI21X1 g60580(.A0 (WX9934), .A1 (_2308_), .B0 (n_337), .Y (n_1097));
AOI21X1 g60581(.A0 (WX9932), .A1 (_2309_), .B0 (n_411), .Y (n_1096));
AOI21X1 g60582(.A0 (WX4734), .A1 (_2194_), .B0 (n_327), .Y (n_1095));
AOI21X1 g60583(.A0 (WX9928), .A1 (_2332_), .B0 (n_305), .Y (n_1094));
AOI21X1 g60584(.A0 (WX9924), .A1 (_2313_), .B0 (n_342), .Y (n_1093));
AOI21X1 g60585(.A0 (WX9920), .A1 (_2315_), .B0 (n_378), .Y (n_1092));
AOI21X1 g60586(.A0 (WX9918), .A1 (_2332_), .B0 (n_282), .Y (n_1091));
AOI21X1 g60587(.A0 (WX9912), .A1 (_2319_), .B0 (n_236), .Y (n_1090));
AOI21X1 g60588(.A0 (WX9910), .A1 (_2320_), .B0 (n_204), .Y (n_1089));
AOI21X1 g60589(.A0 (WX9906), .A1 (_2322_), .B0 (n_361), .Y (n_1088));
AOI21X1 g60590(.A0 (WX9902), .A1 (_2324_), .B0 (n_390), .Y (n_1087));
AOI21X1 g60591(.A0 (WX9898), .A1 (_2326_), .B0 (n_193), .Y (n_1086));
AOI21X1 g60592(.A0 (WX9894), .A1 (_2328_), .B0 (n_379), .Y (n_1085));
AOI21X1 g60593(.A0 (WX11243), .A1 (_2364_), .B0 (n_158), .Y (n_1084));
AOI21X1 g60594(.A0 (WX11239), .A1 (_2334_), .B0 (n_310), .Y (n_1083));
AOI21X1 g60595(.A0 (WX11235), .A1 (_2364_), .B0 (n_294), .Y (n_1082));
AOI21X1 g60596(.A0 (WX11233), .A1 (_2337_), .B0 (n_303), .Y (n_1081));
AOI21X1 g60597(.A0 (WX11225), .A1 (_2341_), .B0 (n_296), .Y (n_1080));
AOI21X1 g60598(.A0 (WX11221), .A1 (_2364_), .B0 (n_208), .Y (n_1079));
AOI21X1 g60599(.A0 (WX11219), .A1 (_2344_), .B0 (n_467), .Y (n_1078));
AOI21X1 g60600(.A0 (WX11215), .A1 (_2346_), .B0 (n_343), .Y (n_1077));
AOI21X1 g60601(.A0 (WX11211), .A1 (_2364_), .B0 (n_371), .Y (n_1076));
AOI21X1 g60602(.A0 (WX11209), .A1 (_2349_), .B0 (n_160), .Y (n_1075));
AOI21X1 g60603(.A0 (WX11205), .A1 (_2351_), .B0 (n_174), .Y (n_1074));
AOI21X1 g60604(.A0 (WX11201), .A1 (_2353_), .B0 (n_260), .Y (n_1073));
AOI21X1 g60605(.A0 (WX11199), .A1 (_2354_), .B0 (n_320), .Y (n_1072));
AOI21X1 g60606(.A0 (WX11197), .A1 (_2355_), .B0 (n_346), .Y (n_1071));
AOI21X1 g60607(.A0 (WX11193), .A1 (_2357_), .B0 (n_442), .Y (n_1070));
AOI21X1 g60608(.A0 (WX11189), .A1 (_2359_), .B0 (n_352), .Y (n_1069));
AOI21X1 g60609(.A0 (WX3467), .A1 (_2149_), .B0 (n_155), .Y (n_1068));
AOI21X1 g60610(.A0 (WX2150), .A1 (_2129_), .B0 (n_360), .Y (n_1067));
AOI21X1 g60611(.A0 (WX4774), .A1 (_2174_), .B0 (n_381), .Y (n_1066));
AOI21X1 g60612(.A0 (WX7312), .A1 (_2262_), .B0 (n_165), .Y (n_1065));
AOI21X1 g60613(.A0 (WX9888), .A1 (_2331_), .B0 (n_413), .Y (n_1064));
AOI21X1 g60614(.A0 (WX9916), .A1 (_2317_), .B0 (n_259), .Y (n_1063));
AOI21X1 g60615(.A0 (WX7348), .A1 (_2244_), .B0 (n_348), .Y (n_1062));
AOI21X1 g60616(.A0 (WX6027), .A1 (_2226_), .B0 (n_335), .Y (n_1061));
AOI21X1 g60617(.A0 (WX2164), .A1 (_2122_), .B0 (n_383), .Y (n_1060));
AOI21X1 g60618(.A0 (WX2188), .A1 (_2110_), .B0 (n_152), .Y (n_1059));
AOI21X1 g60619(.A0 (WX2182), .A1 (_2113_), .B0 (n_149), .Y (n_1058));
AOI21X1 g60620(.A0 (WX3431), .A1 (_2167_), .B0 (n_364), .Y (n_1057));
AOI21X1 g60621(.A0 (WX3433), .A1 (_2166_), .B0 (n_368), .Y (n_1056));
AOI21X1 g60622(.A0 (WX7314), .A1 (_2261_), .B0 (n_159), .Y (n_1055));
AOI21X1 g60624(.A0 (WX7364), .A1 (_2268_), .B0 (n_186), .Y (n_1054));
AOI21X1 g60625(.A0 (WX7318), .A1 (_2259_), .B0 (n_351), .Y (n_1053));
AOI21X1 g60626(.A0 (WX11227), .A1 (_2340_), .B0 (n_363), .Y (n_1052));
AOI21X1 g60627(.A0 (WX9942), .A1 (_2332_), .B0 (n_287), .Y (n_1051));
AOI21X1 g60628(.A0 (WX9908), .A1 (_2321_), .B0 (n_336), .Y (n_1050));
AOI21X1 g60629(.A0 (WX8603), .A1 (_2295_), .B0 (n_292), .Y (n_1049));
AOI21X1 g60630(.A0 (WX9914), .A1 (_2318_), .B0 (n_312), .Y (n_1048));
AOI21X1 g60631(.A0 (WX3477), .A1 (_2172_), .B0 (n_201), .Y (n_1047));
AOI21X1 g60632(.A0 (WX7336), .A1 (_2250_), .B0 (n_191), .Y (n_1046));
AOI21X1 g60633(.A0 (WX2154), .A1 (_2127_), .B0 (n_297), .Y (n_1045));
AOI21X1 g60634(.A0 (WX4756), .A1 (_2204_), .B0 (n_478), .Y (n_1044));
AOI21X1 g60636(.A0 (WX11185), .A1 (_2361_), .B0 (n_168), .Y (n_1043));
AOI21X1 g60637(.A0 (WX9890), .A1 (_2330_), .B0 (n_404), .Y (n_1042));
AOI21X1 g60638(.A0 (WX11237), .A1 (_2335_), .B0 (n_143), .Y (n_1041));
AOI21X1 g60639(.A0 (WX8613), .A1 (_2290_), .B0 (n_319), .Y (n_1040));
AOI21X1 g60640(.A0 (WX8597), .A1 (_2298_), .B0 (n_345), .Y (n_1039));
NOR2X1 g58167(.A (_2107_), .B (WX837), .Y (n_1038));
AOI21X1 g60641(.A0 (WX6065), .A1 (_2207_), .B0 (n_398), .Y (n_1037));
AOI21X1 g60642(.A0 (WX6019), .A1 (_2230_), .B0 (n_137), .Y (n_1036));
AOI21X1 g60643(.A0 (WX7346), .A1 (_2245_), .B0 (n_323), .Y (n_1035));
AOI21X1 g60644(.A0 (WX6015), .A1 (_2232_), .B0 (n_424), .Y (n_1034));
AOI21X1 g60645(.A0 (WX6071), .A1 (_2236_), .B0 (n_344), .Y (n_1033));
AOI21X1 g60646(.A0 (WX4736), .A1 (_2193_), .B0 (n_367), .Y (n_1032));
AOI21X1 g60647(.A0 (WX2178), .A1 (_2115_), .B0 (n_466), .Y (n_1031));
AOI21X1 g60648(.A0 (WX2146), .A1 (_2131_), .B0 (n_255), .Y (n_1030));
AOI21X1 g60651(.A0 (WX2174), .A1 (_2117_), .B0 (n_219), .Y (n_1029));
AOI21X1 g60652(.A0 (WX11223), .A1 (_2342_), .B0 (n_311), .Y (n_1028));
AOI21X1 g60653(.A0 (WX7350), .A1 (_2243_), .B0 (n_290), .Y (n_1027));
AOI21X1 g60654(.A0 (WX2148), .A1 (_2130_), .B0 (n_214), .Y (n_1026));
AOI21X1 g60655(.A0 (WX6055), .A1 (_2212_), .B0 (n_490), .Y (n_1025));
AOI21X1 g60656(.A0 (WX4724), .A1 (_2199_), .B0 (n_190), .Y (n_1024));
AOI21X1 g60659(.A0 (WX2168), .A1 (_2120_), .B0 (n_183), .Y (n_1023));
AOI21X1 g60660(.A0 (WX2192), .A1 (_2140_), .B0 (n_161), .Y (n_1022));
AOI21X1 g60661(.A0 (WX9926), .A1 (_2312_), .B0 (n_370), .Y (n_1021));
AOI21X1 g60663(.A0 (WX9896), .A1 (_2327_), .B0 (n_458), .Y (n_1020));
AOI21X1 g60664(.A0 (WX6045), .A1 (_2217_), .B0 (n_388), .Y (n_1019));
AOI21X1 g60665(.A0 (WX6031), .A1 (_2224_), .B0 (n_321), .Y (n_1018));
AOI21X1 g60666(.A0 (WX4778), .A1 (_2204_), .B0 (n_340), .Y (n_1017));
AOI21X1 g60667(.A0 (WX11191), .A1 (_2358_), .B0 (n_144), .Y (n_1016));
AOI21X1 g60668(.A0 (WX11207), .A1 (_2350_), .B0 (n_210), .Y (n_1015));
AOI21X1 g60669(.A0 (WX2142), .A1 (_2133_), .B0 (n_338), .Y (n_1014));
AOI21X1 g60670(.A0 (WX9892), .A1 (_2329_), .B0 (n_359), .Y (n_1013));
AOI21X1 g60671(.A0 (WX7308), .A1 (_2264_), .B0 (n_286), .Y (n_1012));
CLKBUFX3 g63046(.A (n_1011), .Y (n_1305));
CLKBUFX3 g63041(.A (n_1011), .Y (n_1460));
INVX2 g63023(.A (n_1009), .Y (n_2988));
INVX2 g63024(.A (n_1009), .Y (n_2953));
INVX2 g63018(.A (n_1009), .Y (n_2775));
INVX2 g63012(.A (n_1009), .Y (n_2755));
OR2X1 g61310(.A (n_1006), .B (n_1000), .Y (n_1007));
OR2X1 g61311(.A (n_1004), .B (n_943), .Y (n_1005));
NAND2X1 g61312(.A (n_983), .B (n_1004), .Y (n_1003));
OR2X1 g61315(.A (n_1001), .B (n_1000), .Y (n_1002));
NAND2X1 g61316(.A (n_1001), .B (n_979), .Y (n_999));
OR2X1 g61318(.A (n_997), .B (n_1000), .Y (n_998));
OR2X1 g61320(.A (n_995), .B (n_972), .Y (n_996));
NAND2X1 g61321(.A (n_6511), .B (n_995), .Y (n_994));
OR2X1 g61324(.A (n_992), .B (n_7490), .Y (n_993));
OR2X1 g61325(.A (n_990), .B (n_7490), .Y (n_991));
OR2X1 g61326(.A (n_987), .B (n_7490), .Y (n_988));
OR2X1 g61327(.A (n_985), .B (n_966), .Y (n_986));
NAND2X1 g61328(.A (n_985), .B (n_983), .Y (n_984));
OR2X1 g61331(.A (n_981), .B (n_1000), .Y (n_982));
NAND2X1 g61332(.A (n_981), .B (n_979), .Y (n_980));
OR2X1 g61337(.A (n_977), .B (n_7490), .Y (n_6697));
OR2X1 g61340(.A (n_975), .B (n_943), .Y (n_976));
OR2X1 g61347(.A (n_973), .B (n_972), .Y (n_974));
NAND2X1 g61349(.A (n_970), .B (n_966), .Y (n_971));
OR2X1 g61351(.A (n_970), .B (n_943), .Y (n_969));
NAND2X1 g61352(.A (n_973), .B (n_966), .Y (n_967));
NAND2X1 g61358(.A (n_964), .B (n_966), .Y (n_965));
OR2X1 g61359(.A (n_962), .B (n_966), .Y (n_963));
NAND2X1 g61360(.A (n_962), .B (n_983), .Y (n_960));
OR2X1 g61363(.A (n_958), .B (n_966), .Y (n_959));
OR2X1 g61365(.A (n_956), .B (n_943), .Y (n_957));
NAND2X1 g61370(.A (n_975), .B (n_983), .Y (n_955));
OR2X1 g61371(.A (n_953), .B (n_6432), .Y (n_954));
OR2X1 g61373(.A (n_951), .B (n_943), .Y (n_952));
NAND2X1 g61374(.A (n_951), .B (n_983), .Y (n_950));
OR2X1 g61458(.A (n_948), .B (n_7490), .Y (n_949));
NAND2X1 g61459(.A (n_1006), .B (n_6432), .Y (n_947));
OR2X1 g61460(.A (n_944), .B (n_943), .Y (n_945));
NAND2X1 g61461(.A (n_944), .B (n_966), .Y (n_942));
NAND2X1 g61462(.A (n_940), .B (n_979), .Y (n_941));
OR2X1 g61464(.A (n_938), .B (n_972), .Y (n_939));
NAND2X1 g61465(.A (n_938), .B (n_966), .Y (n_937));
OR2X1 g61469(.A (n_935), .B (n_7490), .Y (n_6699));
NAND2X1 g61470(.A (n_935), .B (n_6433), .Y (n_6698));
OR2X1 g61473(.A (n_932), .B (n_943), .Y (n_933));
NAND2X1 g61474(.A (n_983), .B (n_932), .Y (n_931));
OR2X1 g61477(.A (n_929), .B (n_7490), .Y (n_930));
NAND2X1 g61478(.A (n_927), .B (n_979), .Y (n_928));
NAND2X1 g61479(.A (n_990), .B (n_979), .Y (n_926));
OR2X1 g61480(.A (n_924), .B (n_943), .Y (n_925));
OR2X1 g61481(.A (n_940), .B (n_7490), .Y (n_923));
NAND2X1 g61482(.A (n_924), .B (n_983), .Y (n_922));
OR2X1 g61486(.A (n_920), .B (n_7490), .Y (n_921));
NAND2X1 g61487(.A (n_920), .B (n_6433), .Y (n_919));
OR2X1 g61490(.A (n_964), .B (n_966), .Y (n_918));
NAND2X1 g61492(.A (n_977), .B (n_6433), .Y (n_6696));
NAND2X1 g61499(.A (n_929), .B (n_6433), .Y (n_916));
NAND2X1 g61500(.A (n_956), .B (n_966), .Y (n_915));
OR2X1 g61501(.A (n_913), .B (n_972), .Y (n_914));
NAND2X1 g61503(.A (n_913), .B (n_966), .Y (n_912));
NAND2X1 g61506(.A (n_992), .B (n_6433), .Y (n_911));
NAND2X1 g61508(.A (n_987), .B (n_979), .Y (n_910));
NAND2X1 g61509(.A (n_953), .B (n_6433), .Y (n_909));
NAND2X1 g61511(.A (n_997), .B (n_979), .Y (n_908));
NAND2X1 g61513(.A (n_958), .B (n_966), .Y (n_907));
OR2X1 g61516(.A (n_905), .B (n_7490), .Y (n_906));
NAND2X1 g61517(.A (n_948), .B (n_6433), .Y (n_904));
OR2X1 g61518(.A (n_927), .B (n_7490), .Y (n_903));
NAND2X1 g61519(.A (n_905), .B (n_6433), .Y (n_902));
NOR2X1 g61522(.A (_2083_), .B (WX885), .Y (n_901));
NOR2X1 g61543(.A (_2086_), .B (WX879), .Y (n_900));
NOR2X1 g61547(.A (_2089_), .B (WX873), .Y (n_899));
NOR2X1 g61549(.A (_2108_), .B (WX877), .Y (n_898));
NOR2X1 g61603(.A (_2100_), .B (WX851), .Y (n_897));
INVX2 g63013(.A (n_1009), .Y (n_2770));
NOR2X1 g61831(.A (_2077_), .B (WX897), .Y (n_896));
NOR2X1 g61940(.A (_2096_), .B (WX859), .Y (n_895));
NOR2X1 g61946(.A (_2090_), .B (WX871), .Y (n_894));
NOR2X1 g61979(.A (_2097_), .B (WX857), .Y (n_893));
NOR2X1 g62069(.A (_2088_), .B (WX875), .Y (n_892));
NOR2X1 g62083(.A (_2081_), .B (WX889), .Y (n_891));
NOR2X1 g62103(.A (_2093_), .B (WX865), .Y (n_890));
NOR2X1 g62146(.A (_2105_), .B (WX841), .Y (n_889));
NOR2X1 g62187(.A (_2102_), .B (WX847), .Y (n_888));
NOR2X1 g62214(.A (_2108_), .B (WX891), .Y (n_887));
NOR2X1 g62275(.A (_2103_), .B (WX845), .Y (n_886));
NOR2X1 g62282(.A (_2104_), .B (WX843), .Y (n_885));
NOR2X1 g62301(.A (_2082_), .B (WX887), .Y (n_884));
NOR2X1 g62304(.A (_2106_), .B (WX839), .Y (n_883));
NOR2X1 g62321(.A (_2108_), .B (WX899), .Y (n_882));
NOR2X1 g62337(.A (_2079_), .B (WX893), .Y (n_881));
NOR2X1 g62587(.A (_2099_), .B (WX853), .Y (n_879));
NOR2X1 g62623(.A (_2108_), .B (WX867), .Y (n_878));
NOR2X1 g62689(.A (_2091_), .B (WX869), .Y (n_877));
NOR2X1 g62707(.A (_2094_), .B (WX863), .Y (n_876));
NOR2X1 g62735(.A (_2098_), .B (WX855), .Y (n_875));
NOR2X1 g62751(.A (_2095_), .B (WX861), .Y (n_874));
NOR2X1 g62762(.A (_2101_), .B (WX849), .Y (n_873));
INVX2 g63011(.A (n_1009), .Y (n_2817));
INVX2 g63021(.A (n_1009), .Y (n_3089));
INVX2 g63027(.A (n_1009), .Y (n_2837));
INVX4 g63032(.A (n_880), .Y (n_2744));
INVX2 g63240(.A (n_6512), .Y (n_2986));
INVX1 g63241(.A (n_6512), .Y (n_2838));
INVX4 g63247(.A (n_9424), .Y (n_2795));
INVX4 g63252(.A (n_869), .Y (n_2813));
INVX4 g63253(.A (n_869), .Y (n_2815));
INVX4 g63259(.A (n_868), .Y (n_2716));
INVX4 g63261(.A (n_867), .Y (n_2829));
INVX4 g63263(.A (n_867), .Y (n_2798));
INVX4 g63266(.A (n_866), .Y (n_2935));
INVX4 g63267(.A (n_866), .Y (n_2776));
BUFX3 g63480(.A (n_2298), .Y (n_2246));
BUFX3 g63488(.A (n_2346), .Y (n_2198));
BUFX3 g63489(.A (n_2346), .Y (n_2333));
BUFX3 g63490(.A (n_2346), .Y (n_2223));
BUFX3 g63493(.A (n_2383), .Y (n_2251));
BUFX3 g63494(.A (n_2383), .Y (n_2400));
BUFX3 g63498(.A (n_2383), .Y (n_2218));
BUFX3 g63572(.A (n_2227), .Y (n_2371));
BUFX3 g63574(.A (n_2227), .Y (n_2527));
INVX2 g63592(.A (n_6429), .Y (n_1276));
INVX4 g63612(.A (n_2826), .Y (n_860));
INVX4 g63616(.A (n_2826), .Y (n_858));
INVX2 g63618(.A (n_2826), .Y (n_3031));
INVX8 g63632(.A (n_857), .Y (n_3021));
INVX4 g63646(.A (n_7482), .Y (n_3120));
INVX2 g63652(.A (n_853), .Y (n_3027));
INVX2 g63666(.A (n_7482), .Y (n_1281));
NOR2X1 g61730(.A (_2084_), .B (WX883), .Y (n_852));
INVX4 g63258(.A (n_868), .Y (n_2809));
INVX2 g63248(.A (n_9425), .Y (n_2828));
AOI21X1 g57864(.A0 (WX2066), .A1 (WX2130), .B0 (n_472), .Y (n_850));
AOI21X1 g57865(.A0 (WX11117), .A1 (WX11181), .B0 (n_473), .Y (n_849));
XOR2X1 g57866(.A (n_108), .B (WX2130), .Y (n_848));
XOR2X1 g57870(.A (n_124), .B (WX11181), .Y (n_847));
NOR2X1 g62111(.A (_2085_), .B (WX881), .Y (n_846));
INVX8 g63621(.A (n_857), .Y (n_3137));
INVX4 g63229(.A (n_842), .Y (n_1278));
INVX4 g63222(.A (n_6623), .Y (n_2757));
INVX4 g63598(.A (n_836), .Y (n_1294));
BUFX3 g63571(.A (n_2227), .Y (n_2272));
INVX4 g63581(.A (n_836), .Y (n_3140));
BUFX3 g63573(.A (n_2227), .Y (n_2325));
BUFX3 g63575(.A (n_2227), .Y (n_2529));
BUFX3 g63569(.A (n_2227), .Y (n_2339));
BUFX3 g63570(.A (n_2227), .Y (n_2388));
BUFX3 g63563(.A (n_2227), .Y (n_2396));
BUFX3 g63560(.A (n_2227), .Y (n_2311));
BUFX3 g63561(.A (n_2227), .Y (n_2402));
INVX4 g63516(.A (n_3188), .Y (n_2378));
INVX4 g63501(.A (n_3188), .Y (n_2383));
XOR2X1 g60976(.A (WX8543), .B (WX8607), .Y (n_831));
NAND2X1 g58180(.A (n_0), .B (WX837), .Y (n_830));
INVX8 g63359(.A (n_823), .Y (n_1648));
NAND2X1 g58181(.A (WX773), .B (n_139), .Y (n_817));
INVX2 g63270(.A (n_517), .Y (n_866));
XOR2X1 g60706(.A (WX8583), .B (WX8647), .Y (n_816));
XOR2X1 g60708(.A (WX4668), .B (WX4732), .Y (n_815));
XOR2X1 g60713(.A (WX8587), .B (WX8651), .Y (n_814));
XOR2X1 g60714(.A (WX2068), .B (WX2132), .Y (n_813));
XOR2X1 g60715(.A (WX4670), .B (WX4734), .Y (n_812));
XOR2X1 g60717(.A (WX8589), .B (WX8653), .Y (n_811));
XOR2X1 g60721(.A (WX4672), .B (WX4736), .Y (n_810));
XOR2X1 g60723(.A (WX8593), .B (WX8657), .Y (n_809));
XOR2X1 g60732(.A (WX8541), .B (WX8605), .Y (n_808));
XOR2X1 g60736(.A (WX4680), .B (WX4744), .Y (n_807));
XOR2X1 g60740(.A (WX4684), .B (WX4748), .Y (n_806));
XOR2X1 g60742(.A (WX4686), .B (WX4750), .Y (n_805));
XOR2X1 g60749(.A (WX9824), .B (WX9888), .Y (n_804));
XOR2X1 g60750(.A (WX4682), .B (WX4746), .Y (n_803));
XOR2X1 g60752(.A (WX4714), .B (WX4778), .Y (n_802));
XOR2X1 g60753(.A (WX9826), .B (WX9890), .Y (n_801));
XOR2X1 g60756(.A (WX4690), .B (WX4754), .Y (n_800));
XOR2X1 g60759(.A (WX9828), .B (WX9892), .Y (n_799));
XOR2X1 g60762(.A (WX9830), .B (WX9894), .Y (n_798));
XOR2X1 g60763(.A (WX5999), .B (WX6063), .Y (n_797));
INVX2 g63047(.A (n_520), .Y (n_1011));
XOR2X1 g60767(.A (WX4692), .B (WX4756), .Y (n_796));
XOR2X1 g60768(.A (WX9832), .B (WX9896), .Y (n_795));
XOR2X1 g60771(.A (WX9834), .B (WX9898), .Y (n_794));
XOR2X1 g60772(.A (WX9858), .B (WX9922), .Y (n_793));
XOR2X1 g60775(.A (WX4694), .B (WX4758), .Y (n_792));
XOR2X1 g60777(.A (WX9836), .B (WX9900), .Y (n_791));
XOR2X1 g60783(.A (WX9840), .B (WX9904), .Y (n_790));
XOR2X1 g60790(.A (WX9848), .B (WX9912), .Y (n_789));
XOR2X1 g60791(.A (WX3387), .B (WX3451), .Y (n_788));
XOR2X1 g60792(.A (WX3359), .B (WX3423), .Y (n_787));
XOR2X1 g60794(.A (WX9850), .B (WX9914), .Y (n_786));
XOR2X1 g60798(.A (WX4702), .B (WX4766), .Y (n_785));
XOR2X1 g60799(.A (WX9852), .B (WX9916), .Y (n_784));
XOR2X1 g60806(.A (WX9856), .B (WX9920), .Y (n_783));
XOR2X1 g60809(.A (WX5955), .B (WX6019), .Y (n_782));
XOR2X1 g60812(.A (WX4706), .B (WX4770), .Y (n_781));
XOR2X1 g60814(.A (WX9860), .B (WX9924), .Y (n_780));
XOR2X1 g60815(.A (WX4708), .B (WX4772), .Y (n_779));
XOR2X1 g60817(.A (WX9864), .B (WX9928), .Y (n_778));
XOR2X1 g60824(.A (WX9868), .B (WX9932), .Y (n_777));
XOR2X1 g60836(.A (WX9874), .B (WX9938), .Y (n_776));
XOR2X1 g60839(.A (WX3363), .B (WX3427), .Y (n_775));
XOR2X1 g60841(.A (WX9876), .B (WX9940), .Y (n_774));
XOR2X1 g60844(.A (WX4704), .B (WX4768), .Y (n_773));
XOR2X1 g60845(.A (WX11119), .B (WX11183), .Y (n_772));
NAND2X1 g61520(.A (n_129), .B (WX897), .Y (n_771));
XOR2X1 g60847(.A (WX4674), .B (WX4738), .Y (n_770));
XOR2X1 g60851(.A (WX9880), .B (WX9944), .Y (n_768));
XOR2X1 g60852(.A (WX2070), .B (WX2134), .Y (n_767));
XOR2X1 g60855(.A (WX11131), .B (WX11195), .Y (n_766));
XOR2X1 g60858(.A (WX9884), .B (WX9948), .Y (n_765));
XOR2X1 g60859(.A (WX8537), .B (WX8601), .Y (n_764));
XOR2X1 g61033(.A (WX7248), .B (WX7312), .Y (n_763));
XOR2X1 g60869(.A (WX3367), .B (WX3431), .Y (n_762));
XOR2X1 g60870(.A (WX2096), .B (WX2160), .Y (n_761));
XOR2X1 g60871(.A (WX6005), .B (WX6069), .Y (n_760));
XOR2X1 g60873(.A (WX5977), .B (WX6041), .Y (n_759));
XOR2X1 g60876(.A (WX3369), .B (WX3433), .Y (n_758));
XOR2X1 g60878(.A (WX9854), .B (WX9918), .Y (n_757));
XOR2X1 g60879(.A (WX5945), .B (WX6009), .Y (n_756));
XOR2X1 g60881(.A (WX9878), .B (WX9942), .Y (n_755));
XOR2X1 g60882(.A (WX2074), .B (WX2138), .Y (n_754));
XOR2X1 g60883(.A (WX2076), .B (WX2140), .Y (n_753));
XOR2X1 g60886(.A (WX5947), .B (WX6011), .Y (n_752));
XOR2X1 g60887(.A (WX6001), .B (WX6065), .Y (n_751));
XOR2X1 g60892(.A (WX11125), .B (WX11189), .Y (n_750));
XOR2X1 g60893(.A (WX5949), .B (WX6013), .Y (n_749));
XOR2X1 g60894(.A (WX3371), .B (WX3435), .Y (n_748));
XOR2X1 g60895(.A (WX2088), .B (WX2152), .Y (n_747));
XOR2X1 g60898(.A (WX5951), .B (WX6015), .Y (n_746));
XOR2X1 g60901(.A (WX2078), .B (WX2142), .Y (n_745));
INVX4 g63020(.A (n_769), .Y (n_1009));
XOR2X1 g60913(.A (WX9862), .B (WX9926), .Y (n_744));
XOR2X1 g60914(.A (WX5959), .B (WX6023), .Y (n_743));
XOR2X1 g60915(.A (WX3373), .B (WX3437), .Y (n_742));
XOR2X1 g60917(.A (WX5965), .B (WX6029), .Y (n_741));
XOR2X1 g60919(.A (WX5993), .B (WX6057), .Y (n_740));
XOR2X1 g60921(.A (WX5967), .B (WX6031), .Y (n_739));
XOR2X1 g60927(.A (WX3377), .B (WX3441), .Y (n_738));
XOR2X1 g60928(.A (WX5973), .B (WX6037), .Y (n_737));
XOR2X1 g60930(.A (WX4696), .B (WX4760), .Y (n_736));
XOR2X1 g60931(.A (WX8533), .B (WX8597), .Y (n_735));
XOR2X1 g60934(.A (WX3389), .B (WX3453), .Y (n_734));
XOR2X1 g60935(.A (WX3379), .B (WX3443), .Y (n_733));
XOR2X1 g60937(.A (WX5981), .B (WX6045), .Y (n_732));
XOR2X1 g60939(.A (WX5971), .B (WX6035), .Y (n_731));
XOR2X1 g60940(.A (WX11133), .B (WX11197), .Y (n_730));
XOR2X1 g60941(.A (WX5983), .B (WX6047), .Y (n_729));
XOR2X1 g60942(.A (WX7284), .B (WX7348), .Y (n_728));
XOR2X1 g60943(.A (WX3381), .B (WX3445), .Y (n_727));
XOR2X1 g60947(.A (WX2090), .B (WX2154), .Y (n_726));
XOR2X1 g60949(.A (WX5991), .B (WX6055), .Y (n_725));
XOR2X1 g60956(.A (WX3385), .B (WX3449), .Y (n_724));
XOR2X1 g60961(.A (WX11123), .B (WX11187), .Y (n_723));
XOR2X1 g60963(.A (WX11135), .B (WX11199), .Y (n_722));
XOR2X1 g60969(.A (WX6003), .B (WX6067), .Y (n_721));
XOR2X1 g60977(.A (WX5985), .B (WX6049), .Y (n_720));
XOR2X1 g60979(.A (WX11141), .B (WX11205), .Y (n_719));
XOR2X1 g60982(.A (WX2098), .B (WX2162), .Y (n_718));
XOR2X1 g60984(.A (WX2100), .B (WX2164), .Y (n_717));
XOR2X1 g60985(.A (WX11171), .B (WX11235), .Y (n_716));
XOR2X1 g60986(.A (WX5961), .B (WX6025), .Y (n_715));
XOR2X1 g60987(.A (WX11143), .B (WX11207), .Y (n_714));
XOR2X1 g60990(.A (WX3393), .B (WX3457), .Y (n_713));
XOR2X1 g60997(.A (WX2102), .B (WX2166), .Y (n_712));
XOR2X1 g61005(.A (WX7238), .B (WX7302), .Y (n_711));
XOR2X1 g61006(.A (WX11145), .B (WX11209), .Y (n_710));
XOR2X1 g61007(.A (WX3395), .B (WX3459), .Y (n_709));
XOR2X1 g61015(.A (WX7242), .B (WX7306), .Y (n_708));
XOR2X1 g61016(.A (WX3397), .B (WX3461), .Y (n_707));
XOR2X1 g61017(.A (WX3375), .B (WX3439), .Y (n_706));
XOR2X1 g61019(.A (WX7244), .B (WX7308), .Y (n_705));
XOR2X1 g61025(.A (WX2104), .B (WX2168), .Y (n_704));
XOR2X1 g61027(.A (WX7246), .B (WX7310), .Y (n_703));
XOR2X1 g61028(.A (WX5957), .B (WX6021), .Y (n_702));
XOR2X1 g61029(.A (WX11147), .B (WX11211), .Y (n_701));
XOR2X1 g61030(.A (WX11129), .B (WX11193), .Y (n_700));
XOR2X1 g61036(.A (WX3399), .B (WX3463), .Y (n_699));
XOR2X1 g61038(.A (WX7250), .B (WX7314), .Y (n_698));
XOR2X1 g61042(.A (WX2106), .B (WX2170), .Y (n_697));
XOR2X1 g61043(.A (WX7252), .B (WX7316), .Y (n_696));
XOR2X1 g61047(.A (WX7254), .B (WX7318), .Y (n_695));
XOR2X1 g61050(.A (WX11149), .B (WX11213), .Y (n_693));
XOR2X1 g61052(.A (WX2108), .B (WX2172), .Y (n_692));
XOR2X1 g61054(.A (WX2072), .B (WX2136), .Y (n_691));
XOR2X1 g61055(.A (WX7256), .B (WX7320), .Y (n_690));
XOR2X1 g61064(.A (WX3401), .B (WX3465), .Y (n_689));
XOR2X1 g61065(.A (WX4712), .B (WX4776), .Y (n_688));
XOR2X1 g61066(.A (WX3417), .B (WX3481), .Y (n_687));
XOR2X1 g61074(.A (WX7262), .B (WX7326), .Y (n_686));
XOR2X1 g61075(.A (WX11151), .B (WX11215), .Y (n_685));
XOR2X1 g61078(.A (WX7264), .B (WX7328), .Y (n_684));
XOR2X1 g61079(.A (WX4666), .B (WX4730), .Y (n_683));
XOR2X1 g61081(.A (WX2110), .B (WX2174), .Y (n_682));
XOR2X1 g61085(.A (WX7266), .B (WX7330), .Y (n_681));
XOR2X1 g61090(.A (WX2112), .B (WX2176), .Y (n_680));
XOR2X1 g61093(.A (WX8579), .B (WX8643), .Y (n_679));
XOR2X1 g61096(.A (WX7270), .B (WX7334), .Y (n_678));
XOR2X1 g61098(.A (WX11153), .B (WX11217), .Y (n_677));
XOR2X1 g61100(.A (WX3405), .B (WX3469), .Y (n_676));
XOR2X1 g61101(.A (WX7272), .B (WX7336), .Y (n_675));
XOR2X1 g61102(.A (WX9870), .B (WX9934), .Y (n_674));
XOR2X1 g61107(.A (WX3407), .B (WX3471), .Y (n_673));
XOR2X1 g61109(.A (WX7276), .B (WX7340), .Y (n_672));
XOR2X1 g61110(.A (WX5953), .B (WX6017), .Y (n_671));
XOR2X1 g61111(.A (WX9846), .B (WX9910), .Y (n_670));
XOR2X1 g61114(.A (WX7278), .B (WX7342), .Y (n_669));
XOR2X1 g61116(.A (WX2114), .B (WX2178), .Y (n_668));
XOR2X1 g61118(.A (WX2084), .B (WX2148), .Y (n_667));
XOR2X1 g61119(.A (WX7280), .B (WX7344), .Y (n_666));
XOR2X1 g61120(.A (WX11155), .B (WX11219), .Y (n_665));
XOR2X1 g61124(.A (WX2116), .B (WX2180), .Y (n_664));
XOR2X1 g61125(.A (WX7282), .B (WX7346), .Y (n_663));
XOR2X1 g61128(.A (WX3409), .B (WX3473), .Y (n_662));
XOR2X1 g61130(.A (WX7286), .B (WX7350), .Y (n_661));
XOR2X1 g61135(.A (WX7288), .B (WX7352), .Y (n_660));
XOR2X1 g61136(.A (WX11157), .B (WX11221), .Y (n_659));
XOR2X1 g61137(.A (WX2118), .B (WX2182), .Y (n_658));
XOR2X1 g61141(.A (WX7290), .B (WX7354), .Y (n_657));
XOR2X1 g61000(.A (WX2124), .B (WX2188), .Y (n_656));
XOR2X1 g61143(.A (WX3411), .B (WX3475), .Y (n_655));
XOR2X1 g61148(.A (WX7294), .B (WX7358), .Y (n_654));
XOR2X1 g61153(.A (WX3413), .B (WX3477), .Y (n_653));
XOR2X1 g61155(.A (WX7296), .B (WX7360), .Y (n_652));
XOR2X1 g61158(.A (WX11159), .B (WX11223), .Y (n_651));
XOR2X1 g61159(.A (WX11127), .B (WX11191), .Y (n_650));
XOR2X1 g61162(.A (WX7298), .B (WX7362), .Y (n_649));
XOR2X1 g61163(.A (WX2120), .B (WX2184), .Y (n_648));
XOR2X1 g61164(.A (WX5975), .B (WX6039), .Y (n_647));
XOR2X1 g61165(.A (WX8575), .B (WX8639), .Y (n_646));
XOR2X1 g61168(.A (WX7300), .B (WX7364), .Y (n_645));
XOR2X1 g61172(.A (WX2122), .B (WX2186), .Y (n_644));
XOR2X1 g61174(.A (WX9844), .B (WX9908), .Y (n_643));
XOR2X1 g61175(.A (WX3415), .B (WX3479), .Y (n_642));
XOR2X1 g61176(.A (WX11161), .B (WX11225), .Y (n_641));
XOR2X1 g61181(.A (WX2126), .B (WX2190), .Y (n_640));
XOR2X1 g61186(.A (WX3419), .B (WX3483), .Y (n_639));
XOR2X1 g61191(.A (WX3421), .B (WX3485), .Y (n_638));
XOR2X1 g61198(.A (WX4710), .B (WX4774), .Y (n_637));
XOR2X1 g61199(.A (WX11167), .B (WX11231), .Y (n_636));
XOR2X1 g61203(.A (WX11169), .B (WX11233), .Y (n_635));
XOR2X1 g61204(.A (WX4662), .B (WX4726), .Y (n_634));
XOR2X1 g61205(.A (WX5979), .B (WX6043), .Y (n_633));
XOR2X1 g61207(.A (WX2086), .B (WX2150), .Y (n_632));
XOR2X1 g61210(.A (WX9866), .B (WX9930), .Y (n_631));
XOR2X1 g61211(.A (WX8531), .B (WX8595), .Y (n_630));
XOR2X1 g61216(.A (WX8535), .B (WX8599), .Y (n_629));
XOR2X1 g61217(.A (WX2082), .B (WX2146), .Y (n_628));
XOR2X1 g61222(.A (WX8539), .B (WX8603), .Y (n_627));
XOR2X1 g61223(.A (WX11173), .B (WX11237), .Y (n_626));
XOR2X1 g61224(.A (WX6007), .B (WX6071), .Y (n_625));
XOR2X1 g61231(.A (WX8571), .B (WX8635), .Y (n_624));
XOR2X1 g61232(.A (WX9842), .B (WX9906), .Y (n_623));
XOR2X1 g61235(.A (WX2094), .B (WX2158), .Y (n_622));
XOR2X1 g61236(.A (WX8545), .B (WX8609), .Y (n_621));
XOR2X1 g61241(.A (WX8547), .B (WX8611), .Y (n_620));
XOR2X1 g61242(.A (WX9838), .B (WX9902), .Y (n_619));
XOR2X1 g61243(.A (WX11175), .B (WX11239), .Y (n_618));
XOR2X1 g61245(.A (WX8549), .B (WX8613), .Y (n_617));
XOR2X1 g61250(.A (WX8551), .B (WX8615), .Y (n_616));
XOR2X1 g61251(.A (WX4652), .B (WX4716), .Y (n_615));
XOR2X1 g61260(.A (WX8555), .B (WX8619), .Y (n_614));
XOR2X1 g61264(.A (WX11177), .B (WX11241), .Y (n_613));
XOR2X1 g61267(.A (WX8557), .B (WX8621), .Y (n_612));
XOR2X1 g61268(.A (WX3391), .B (WX3455), .Y (n_611));
XOR2X1 g61273(.A (WX4656), .B (WX4720), .Y (n_610));
XOR2X1 g61275(.A (WX8561), .B (WX8625), .Y (n_609));
XOR2X1 g61280(.A (WX8563), .B (WX8627), .Y (n_608));
XOR2X1 g61281(.A (WX4658), .B (WX4722), .Y (n_607));
XOR2X1 g61282(.A (WX11179), .B (WX11243), .Y (n_606));
XOR2X1 g61289(.A (WX8567), .B (WX8631), .Y (n_605));
XOR2X1 g61290(.A (WX4660), .B (WX4724), .Y (n_604));
XOR2X1 g61297(.A (WX8573), .B (WX8637), .Y (n_603));
XOR2X1 g61298(.A (WX3383), .B (WX3447), .Y (n_602));
XOR2X1 g61301(.A (WX4664), .B (WX4728), .Y (n_601));
XOR2X1 g61302(.A (WX8577), .B (WX8641), .Y (n_600));
XOR2X1 g61303(.A (WX9886), .B (WX9950), .Y (n_599));
XOR2X1 g61309(.A (WX8581), .B (WX8645), .Y (n_598));
NAND2X1 g61313(.A (WX817), .B (n_261), .Y (n_597));
NAND2X1 g61314(.A (n_70), .B (WX881), .Y (n_596));
NAND2X1 g61317(.A (n_69), .B (WX887), .Y (n_595));
NAND2X1 g61319(.A (n_24), .B (WX847), .Y (n_594));
NAND2X1 g61322(.A (WX819), .B (n_484), .Y (n_593));
NAND2X1 g61323(.A (n_79), .B (WX859), .Y (n_592));
NAND2X1 g61329(.A (WX801), .B (n_462), .Y (n_591));
NAND2X1 g61330(.A (n_130), .B (WX885), .Y (n_590));
NAND2X1 g61333(.A (WX795), .B (n_280), .Y (n_589));
NAND2X1 g61334(.A (WX783), .B (n_252), .Y (n_588));
NAND2X1 g61335(.A (WX823), .B (n_266), .Y (n_587));
NAND2X1 g61338(.A (n_117), .B (WX867), .Y (n_586));
NAND2X1 g61339(.A (WX829), .B (n_451), .Y (n_585));
NAND2X1 g61342(.A (WX825), .B (n_268), .Y (n_584));
NAND2X1 g61343(.A (n_98), .B (WX849), .Y (n_583));
NAND2X1 g61344(.A (WX785), .B (n_420), .Y (n_582));
NAND2X1 g61345(.A (WX799), .B (n_438), .Y (n_581));
NAND2X1 g61346(.A (n_3), .B (WX889), .Y (n_580));
NAND2X1 g61348(.A (n_89), .B (WX861), .Y (n_579));
NAND2X1 g61354(.A (WX827), .B (n_448), .Y (n_578));
NAND2X1 g61355(.A (n_81), .B (WX841), .Y (n_577));
NAND2X1 g61356(.A (n_58), .B (WX891), .Y (n_576));
NAND2X1 g61357(.A (WX777), .B (n_273), .Y (n_575));
NAND2X1 g61361(.A (n_68), .B (WX893), .Y (n_574));
NAND2X1 g61362(.A (n_96), .B (WX883), .Y (n_573));
NAND2X1 g61364(.A (WX835), .B (n_480), .Y (n_572));
NAND2X1 g61366(.A (n_28), .B (WX865), .Y (n_571));
NAND2X1 g61367(.A (WX831), .B (n_278), .Y (n_570));
NAND2X1 g61368(.A (n_5), .B (WX895), .Y (n_569));
NAND2X1 g61369(.A (WX821), .B (n_482), .Y (n_568));
NAND2X1 g61372(.A (n_83), .B (WX839), .Y (n_567));
NAND2X1 g61375(.A (n_41), .B (WX843), .Y (n_566));
NAND2X1 g61463(.A (WX787), .B (n_454), .Y (n_565));
NAND2X1 g61466(.A (WX805), .B (n_474), .Y (n_564));
NAND2X1 g61467(.A (n_118), .B (WX869), .Y (n_563));
NAND2X1 g61471(.A (WX789), .B (n_264), .Y (n_562));
NAND2X1 g61472(.A (WX797), .B (n_244), .Y (n_561));
NAND2X1 g61475(.A (n_27), .B (WX853), .Y (n_560));
NAND2X1 g61476(.A (WX807), .B (n_283), .Y (n_559));
NAND2X1 g61483(.A (WX809), .B (n_486), .Y (n_558));
NAND2X1 g61484(.A (WX781), .B (n_308), .Y (n_557));
NAND2X1 g61485(.A (n_33), .B (WX873), .Y (n_556));
NAND2X1 g61488(.A (n_40), .B (WX845), .Y (n_555));
NAND2X1 g61489(.A (WX791), .B (n_434), .Y (n_554));
NAND2X1 g61491(.A (n_35), .B (WX855), .Y (n_553));
NAND2X1 g61493(.A (WX811), .B (n_429), .Y (n_552));
NAND2X1 g61494(.A (WX779), .B (n_436), .Y (n_551));
NAND2X1 g61495(.A (n_126), .B (WX899), .Y (n_550));
NAND2X1 g61496(.A (n_21), .B (WX875), .Y (n_549));
NAND2X1 g61497(.A (WX833), .B (n_443), .Y (n_548));
NAND2X1 g61498(.A (n_119), .B (WX871), .Y (n_547));
NAND2X1 g61502(.A (WX803), .B (n_476), .Y (n_546));
NAND2X1 g61504(.A (WX813), .B (n_271), .Y (n_545));
NAND2X1 g61505(.A (n_49), .B (WX877), .Y (n_544));
NAND2X1 g61507(.A (n_73), .B (WX879), .Y (n_543));
NAND2X1 g61510(.A (n_56), .B (WX851), .Y (n_542));
NAND2X1 g61512(.A (WX793), .B (n_354), .Y (n_541));
NAND2X1 g61514(.A (WX815), .B (n_431), .Y (n_540));
NAND2X1 g61515(.A (n_38), .B (WX857), .Y (n_539));
XOR2X1 g60972(.A (WX8585), .B (WX8649), .Y (n_538));
XOR2X1 g60959(.A (WX2092), .B (WX2156), .Y (n_537));
XOR2X1 g60955(.A (WX5995), .B (WX6059), .Y (n_536));
XOR2X1 g60923(.A (WX5969), .B (WX6033), .Y (n_535));
INVX4 g63483(.A (n_3188), .Y (n_2298));
XOR2X1 g60908(.A (WX2080), .B (WX2144), .Y (n_532));
XOR2X1 g60904(.A (WX5963), .B (WX6027), .Y (n_531));
XOR2X1 g60862(.A (WX11121), .B (WX11185), .Y (n_530));
XOR2X1 g60854(.A (WX9882), .B (WX9946), .Y (n_529));
XOR2X1 g60831(.A (WX9872), .B (WX9936), .Y (n_527));
XOR2X1 g60829(.A (WX5989), .B (WX6053), .Y (n_526));
XOR2X1 g60823(.A (WX3361), .B (WX3425), .Y (n_525));
NAND2X1 g61353(.A (n_36), .B (WX863), .Y (n_524));
NAND2X1 g61350(.A (WX775), .B (n_276), .Y (n_523));
XOR2X1 g60789(.A (WX4700), .B (WX4764), .Y (n_522));
XOR2X1 g60786(.A (WX4698), .B (WX4762), .Y (n_521));
CLKBUFX3 g63036(.A (n_520), .Y (n_880));
XOR2X1 g60760(.A (WX11139), .B (WX11203), .Y (n_519));
XOR2X1 g61306(.A (WX5987), .B (WX6051), .Y (n_518));
INVX2 g63255(.A (n_517), .Y (n_869));
XOR2X1 g61292(.A (WX8569), .B (WX8633), .Y (n_516));
XOR2X1 g60748(.A (WX4688), .B (WX4752), .Y (n_515));
XOR2X1 g61284(.A (WX8565), .B (WX8629), .Y (n_514));
INVX2 g63235(.A (n_943), .Y (n_842));
INVX2 g63260(.A (n_517), .Y (n_868));
INVX2 g63265(.A (n_517), .Y (n_867));
INVX8 g63418(.A (n_471), .Y (n_5712));
INVX4 g63492(.A (n_3188), .Y (n_2346));
XOR2X1 g61270(.A (WX8559), .B (WX8623), .Y (n_510));
XOR2X1 g61263(.A (WX4654), .B (WX4718), .Y (n_509));
XOR2X1 g60734(.A (WX4678), .B (WX4742), .Y (n_508));
XOR2X1 g60720(.A (WX8591), .B (WX8655), .Y (n_507));
XOR2X1 g61253(.A (WX8553), .B (WX8617), .Y (n_506));
INVX8 g63319(.A (n_471), .Y (n_5181));
XOR2X1 g61247(.A (WX5997), .B (WX6061), .Y (n_505));
XOR2X1 g61240(.A (WX11137), .B (WX11201), .Y (n_504));
INVX8 g63447(.A (n_471), .Y (n_1425));
XOR2X1 g61214(.A (WX3365), .B (WX3429), .Y (n_503));
XOR2X1 g61193(.A (WX2128), .B (WX2192), .Y (n_502));
XOR2X1 g61190(.A (WX11165), .B (WX11229), .Y (n_501));
XOR2X1 g61180(.A (WX11163), .B (WX11227), .Y (n_500));
XOR2X1 g61145(.A (WX7292), .B (WX7356), .Y (n_499));
INVX2 g63653(.A (n_7487), .Y (n_853));
XOR2X1 g61105(.A (WX7274), .B (WX7338), .Y (n_497));
INVX1 g63643(.A (n_7487), .Y (n_2800));
XOR2X1 g61089(.A (WX7268), .B (WX7332), .Y (n_496));
XOR2X1 g61073(.A (WX3403), .B (WX3467), .Y (n_495));
INVX4 g63630(.A (n_1000), .Y (n_857));
INVX4 g63604(.A (n_6431), .Y (n_836));
INVX8 g63619(.A (n_6432), .Y (n_2826));
XOR2X1 g61068(.A (WX7260), .B (WX7324), .Y (n_492));
INVX8 g63567(.A (n_3188), .Y (n_2227));
XOR2X1 g61061(.A (WX7258), .B (WX7322), .Y (n_491));
NOR2X1 g62558(.A (WX6055), .B (_2212_), .Y (n_490));
NOR2X1 g62559(.A (WX3473), .B (_2146_), .Y (n_489));
NOR2X1 g62095(.A (WX3459), .B (_2153_), .Y (n_488));
NOR2X1 g61590(.A (WX4728), .B (_2197_), .Y (n_479));
NOR2X1 g61538(.A (WX4756), .B (_2204_), .Y (n_478));
NOR2X1 g58179(.A (WX11117), .B (WX11181), .Y (n_473));
NOR2X1 g58178(.A (WX2066), .B (WX2130), .Y (n_472));
NOR2X1 g62750(.A (WX6043), .B (_2218_), .Y (n_470));
NOR2X1 g61574(.A (WX2184), .B (_2140_), .Y (n_469));
NOR2X1 g61575(.A (WX7328), .B (_2254_), .Y (n_468));
NOR2X1 g61576(.A (WX11219), .B (_2344_), .Y (n_467));
NOR2X1 g62049(.A (WX2178), .B (_2115_), .Y (n_466));
NOR2X1 g61569(.A (WX4720), .B (_2201_), .Y (n_465));
NOR2X1 g61560(.A (WX3475), .B (_2145_), .Y (n_464));
NOR2X1 g62029(.A (WX8621), .B (_2286_), .Y (n_461));
NOR2X1 g62591(.A (WX3429), .B (_2168_), .Y (n_460));
INVX2 g63048(.A (n_456), .Y (n_520));
NOR2X1 g61544(.A (WX9896), .B (_2327_), .Y (n_458));
NOR2X1 g61545(.A (WX3463), .B (_2172_), .Y (n_457));
CLKBUFX3 g63031(.A (n_456), .Y (n_769));
NOR2X1 g62040(.A (WX6047), .B (_2216_), .Y (n_453));
INVX4 g63009(.A (n_450), .Y (n_966));
NOR2X1 g62578(.A (WX8657), .B (_2300_), .Y (n_447));
NOR2X1 g62579(.A (WX11193), .B (_2357_), .Y (n_442));
NOR2X1 g62580(.A (WX8645), .B (_2274_), .Y (n_440));
NOR2X1 g62357(.A (WX7310), .B (_2263_), .Y (n_433));
NOR2X1 g61913(.A (WX9922), .B (_2314_), .Y (n_428));
NOR2X1 g62568(.A (WX3435), .B (_2165_), .Y (n_427));
NOR2X1 g61897(.A (WX8635), .B (_2300_), .Y (n_426));
NOR2X1 g62522(.A (WX6015), .B (_2232_), .Y (n_424));
NOR2X1 g61534(.A (WX3461), .B (_2152_), .Y (n_423));
NOR2X1 g61536(.A (WX4746), .B (_2204_), .Y (n_422));
NOR2X1 g61567(.A (WX7302), .B (_2267_), .Y (n_419));
NOR2X1 g62561(.A (WX6017), .B (_2231_), .Y (n_418));
NOR2X1 g62071(.A (WX8647), .B (_2273_), .Y (n_417));
NOR2X1 g61602(.A (WX7322), .B (_2257_), .Y (n_416));
NOR2X1 g61525(.A (WX8643), .B (_2275_), .Y (n_415));
NOR2X1 g61635(.A (WX3457), .B (_2154_), .Y (n_414));
NOR2X1 g61637(.A (WX9888), .B (_2331_), .Y (n_413));
NOR2X1 g61645(.A (WX9936), .B (_2307_), .Y (n_412));
NOR2X1 g61651(.A (WX9932), .B (_2309_), .Y (n_411));
NOR2X1 g61659(.A (WX8609), .B (_2292_), .Y (n_410));
NOR2X1 g61669(.A (WX11183), .B (_2362_), .Y (n_409));
NOR2X1 g61674(.A (WX6025), .B (_2227_), .Y (n_408));
NOR2X1 g61695(.A (WX9946), .B (_2302_), .Y (n_407));
NOR2X1 g61709(.A (WX6057), .B (_2211_), .Y (n_406));
NOR2X1 g61710(.A (WX11187), .B (_2360_), .Y (n_405));
NOR2X1 g61713(.A (WX9890), .B (_2330_), .Y (n_404));
NOR2X1 g61722(.A (WX8611), .B (_2291_), .Y (n_403));
NOR2X1 g61726(.A (WX3483), .B (_2141_), .Y (n_402));
NOR2X1 g61742(.A (WX3481), .B (_2142_), .Y (n_401));
NOR2X1 g62538(.A (WX2180), .B (_2114_), .Y (n_399));
NOR2X1 g61782(.A (WX6065), .B (_2207_), .Y (n_398));
NOR2X1 g61785(.A (WX6053), .B (_2213_), .Y (n_397));
NOR2X1 g61788(.A (WX3449), .B (_2158_), .Y (n_396));
NOR2X1 g61789(.A (WX3439), .B (_2163_), .Y (n_395));
NOR2X1 g61792(.A (WX3423), .B (_2171_), .Y (n_394));
NOR2X1 g61804(.A (WX7332), .B (_2268_), .Y (n_393));
NOR2X1 g61824(.A (WX6035), .B (_2222_), .Y (n_392));
NOR2X1 g61830(.A (WX4772), .B (_2175_), .Y (n_391));
NOR2X1 g61836(.A (WX9902), .B (_2324_), .Y (n_390));
NOR2X1 g61842(.A (WX3445), .B (_2160_), .Y (n_389));
NOR2X1 g61845(.A (WX6045), .B (_2217_), .Y (n_388));
NOR2X1 g61860(.A (WX3427), .B (_2169_), .Y (n_387));
NOR2X1 g61876(.A (WX11229), .B (_2339_), .Y (n_386));
NOR2X1 g61882(.A (WX2176), .B (_2116_), .Y (n_385));
NOR2X1 g61885(.A (WX7338), .B (_2249_), .Y (n_384));
NOR2X1 g61888(.A (WX2164), .B (_2122_), .Y (n_383));
NOR2X1 g61896(.A (WX8651), .B (_2271_), .Y (n_382));
NOR2X1 g61903(.A (WX4774), .B (_2174_), .Y (n_381));
NOR2X1 g61909(.A (WX7306), .B (_2265_), .Y (n_380));
NOR2X1 g61911(.A (WX9894), .B (_2328_), .Y (n_379));
NOR2X1 g61916(.A (WX9920), .B (_2315_), .Y (n_378));
NOR2X1 g61918(.A (WX3469), .B (_2148_), .Y (n_377));
NOR2X1 g61922(.A (WX2190), .B (_2109_), .Y (n_376));
NOR2X1 g61923(.A (WX9938), .B (_2306_), .Y (n_375));
NOR2X1 g61679(.A (WX3465), .B (_2150_), .Y (n_374));
NOR2X1 g61942(.A (WX2136), .B (_2136_), .Y (n_373));
NOR2X1 g61954(.A (WX6029), .B (_2225_), .Y (n_372));
NOR2X1 g61975(.A (WX11211), .B (_2364_), .Y (n_371));
NOR2X1 g61977(.A (WX9926), .B (_2312_), .Y (n_370));
NOR2X1 g62006(.A (WX8649), .B (_2300_), .Y (n_369));
NOR2X1 g62028(.A (WX3433), .B (_2166_), .Y (n_368));
NOR2X1 g62031(.A (WX4736), .B (_2193_), .Y (n_367));
NOR2X1 g62032(.A (WX8637), .B (_2278_), .Y (n_366));
NOR2X1 g62035(.A (WX2156), .B (_2126_), .Y (n_365));
NOR2X1 g62037(.A (WX3431), .B (_2167_), .Y (n_364));
NOR2X1 g62039(.A (WX11227), .B (_2340_), .Y (n_363));
NOR2X1 g62053(.A (WX8607), .B (_2293_), .Y (n_362));
NOR2X1 g62054(.A (WX9906), .B (_2322_), .Y (n_361));
NOR2X1 g62056(.A (WX2150), .B (_2129_), .Y (n_360));
NOR2X1 g62070(.A (WX9892), .B (_2329_), .Y (n_359));
NOR2X1 g62079(.A (WX8623), .B (_2285_), .Y (n_358));
NOR2X1 g62093(.A (WX4726), .B (_2198_), .Y (n_357));
NOR2X1 g62105(.A (WX3453), .B (_2172_), .Y (n_356));
NOR2X1 g62109(.A (WX4730), .B (_2196_), .Y (n_353));
NOR2X1 g62115(.A (WX11189), .B (_2359_), .Y (n_352));
NOR2X1 g62125(.A (WX7318), .B (_2259_), .Y (n_351));
NOR2X1 g62134(.A (WX7344), .B (_2246_), .Y (n_350));
NOR2X1 g62141(.A (WX11195), .B (_2356_), .Y (n_349));
NOR2X1 g62147(.A (WX7348), .B (_2244_), .Y (n_348));
NOR2X1 g62152(.A (WX6039), .B (_2236_), .Y (n_347));
NOR2X1 g62154(.A (WX11197), .B (_2355_), .Y (n_346));
NOR2X1 g62157(.A (WX8597), .B (_2298_), .Y (n_345));
NOR2X1 g62159(.A (WX6071), .B (_2236_), .Y (n_344));
NOR2X1 g62170(.A (WX11215), .B (_2346_), .Y (n_343));
NOR2X1 g62192(.A (WX9924), .B (_2313_), .Y (n_342));
NOR2X1 g62198(.A (WX3441), .B (_2162_), .Y (n_341));
NOR2X1 g62204(.A (WX4778), .B (_2204_), .Y (n_340));
NOR2X1 g62212(.A (WX6011), .B (_2234_), .Y (n_339));
NOR2X1 g62216(.A (WX2142), .B (_2133_), .Y (n_338));
NOR2X1 g62217(.A (WX9934), .B (_2308_), .Y (n_337));
NOR2X1 g62227(.A (WX9908), .B (_2321_), .Y (n_336));
NOR2X1 g62232(.A (WX6027), .B (_2226_), .Y (n_335));
NOR2X1 g62234(.A (WX7304), .B (_2266_), .Y (n_334));
NOR2X1 g62239(.A (WX9948), .B (_2301_), .Y (n_333));
NOR2X1 g62242(.A (WX4732), .B (_2195_), .Y (n_332));
NOR2X1 g62246(.A (WX4722), .B (_2200_), .Y (n_331));
NOR2X1 g62251(.A (WX8595), .B (_2299_), .Y (n_330));
NOR2X1 g62254(.A (WX9904), .B (_2323_), .Y (n_329));
NOR2X1 g62266(.A (WX6069), .B (_2205_), .Y (n_328));
NOR2X1 g62271(.A (WX4734), .B (_2194_), .Y (n_327));
NOR2X1 g62273(.A (WX2166), .B (_2121_), .Y (n_326));
NOR2X1 g62278(.A (WX2152), .B (_2128_), .Y (n_325));
NOR2X1 g62292(.A (WX6041), .B (_2219_), .Y (n_324));
NOR2X1 g62300(.A (WX7346), .B (_2245_), .Y (n_323));
NOR2X1 g62302(.A (WX4752), .B (_2185_), .Y (n_322));
NOR2X1 g62310(.A (WX6031), .B (_2224_), .Y (n_321));
NOR2X1 g62323(.A (WX11199), .B (_2354_), .Y (n_320));
NOR2X1 g62328(.A (WX8613), .B (_2290_), .Y (n_319));
NOR2X1 g62339(.A (WX8627), .B (_2283_), .Y (n_318));
NOR2X1 g62343(.A (WX8605), .B (_2294_), .Y (n_317));
NOR2X1 g62346(.A (WX7354), .B (_2241_), .Y (n_316));
NOR2X1 g62351(.A (WX6067), .B (_2206_), .Y (n_315));
NOR2X1 g62352(.A (WX3479), .B (_2143_), .Y (n_314));
NOR2X1 g62358(.A (WX3471), .B (_2147_), .Y (n_313));
NOR2X1 g62360(.A (WX9914), .B (_2318_), .Y (n_312));
NOR2X1 g62361(.A (WX11223), .B (_2342_), .Y (n_311));
NOR2X1 g62525(.A (WX11239), .B (_2334_), .Y (n_310));
NOR2X1 g62508(.A (WX6049), .B (_2236_), .Y (n_307));
NOR2X1 g62507(.A (WX2160), .B (_2140_), .Y (n_306));
NOR2X1 g62505(.A (WX9928), .B (_2332_), .Y (n_305));
NOR2X1 g62476(.A (WX2140), .B (_2134_), .Y (n_304));
NOR2X1 g62479(.A (WX11233), .B (_2337_), .Y (n_303));
NOR2X1 g62506(.A (WX9930), .B (_2310_), .Y (n_302));
NOR2X1 g62575(.A (WX6037), .B (_2221_), .Y (n_301));
NOR2X1 g62583(.A (WX4716), .B (_2203_), .Y (n_300));
NOR2X1 g62590(.A (WX3443), .B (_2161_), .Y (n_299));
NOR2X1 g62592(.A (WX8617), .B (_2288_), .Y (n_298));
NOR2X1 g62611(.A (WX2154), .B (_2127_), .Y (n_297));
NOR2X1 g61548(.A (WX11225), .B (_2341_), .Y (n_296));
NOR2X1 g62631(.A (WX6023), .B (_2228_), .Y (n_295));
NOR2X1 g62634(.A (WX11235), .B (_2364_), .Y (n_294));
NOR2X1 g62654(.A (WX8599), .B (_2297_), .Y (n_293));
NOR2X1 g62691(.A (WX8603), .B (_2295_), .Y (n_292));
NOR2X1 g62695(.A (WX2186), .B (_2111_), .Y (n_291));
NOR2X1 g62477(.A (WX7350), .B (_2243_), .Y (n_290));
NOR2X1 g62705(.A (WX8655), .B (_2269_), .Y (n_289));
NOR2X1 g61941(.A (WX8639), .B (_2277_), .Y (n_288));
NOR2X1 g62712(.A (WX9942), .B (_2332_), .Y (n_287));
NOR2X1 g62727(.A (WX7308), .B (_2264_), .Y (n_286));
NOR2X1 g62739(.A (WX11213), .B (_2347_), .Y (n_285));
NOR2X1 g62754(.A (WX9918), .B (_2332_), .Y (n_282));
NOR2X1 g61910(.A (WX11201), .B (_2353_), .Y (n_260));
NOR2X1 g61912(.A (WX9916), .B (_2317_), .Y (n_259));
NOR2X1 g61908(.A (WX4760), .B (_2181_), .Y (n_258));
NOR2X1 g62375(.A (WX11231), .B (_2338_), .Y (n_257));
NOR2X1 g62524(.A (WX7330), .B (_2253_), .Y (n_256));
NOR2X1 g61899(.A (WX2146), .B (_2131_), .Y (n_255));
NOR2X1 g61898(.A (WX4750), .B (_2186_), .Y (n_254));
NOR2X1 g61889(.A (WX2134), .B (_2137_), .Y (n_247));
NOR2X1 g61872(.A (WX9950), .B (_2332_), .Y (n_241));
NOR2X1 g61857(.A (WX9912), .B (_2319_), .Y (n_236));
NOR2X1 g62347(.A (WX2158), .B (_2125_), .Y (n_235));
INVX2 g63272(.A (n_6510), .Y (n_983));
NOR2X1 g62764(.A (WX7320), .B (_2258_), .Y (n_233));
NOR2X1 g62340(.A (WX3437), .B (_2164_), .Y (n_232));
NOR2X1 g62765(.A (WX7352), .B (_2242_), .Y (n_231));
NOR2X1 g61852(.A (WX7324), .B (_2256_), .Y (n_230));
NOR2X1 g62757(.A (WX2132), .B (_2138_), .Y (n_229));
NOR2X1 g61846(.A (WX2170), .B (_2140_), .Y (n_228));
NOR2X1 g61841(.A (WX7362), .B (_2237_), .Y (n_227));
NOR2X1 g62752(.A (WX8615), .B (_2289_), .Y (n_226));
INVX2 g63271(.A (n_6510), .Y (n_517));
NOR2X1 g61833(.A (WX8633), .B (_2280_), .Y (n_225));
NOR2X1 g62527(.A (WX2174), .B (_2117_), .Y (n_219));
NOR2X1 g61821(.A (WX2148), .B (_2130_), .Y (n_214));
NOR2X1 g62743(.A (WX8641), .B (_2276_), .Y (n_213));
NOR2X1 g61815(.A (WX6063), .B (_2236_), .Y (n_212));
NOR2X1 g61814(.A (WX7358), .B (_2239_), .Y (n_211));
NOR2X1 g61991(.A (WX11207), .B (_2350_), .Y (n_210));
NOR2X1 g62293(.A (WX2162), .B (_2123_), .Y (n_209));
NOR2X1 g61793(.A (WX11221), .B (_2364_), .Y (n_208));
NOR2X1 g62740(.A (WX9944), .B (_2303_), .Y (n_207));
NOR2X1 g62287(.A (WX3451), .B (_2157_), .Y (n_206));
NOR2X1 g62734(.A (WX2144), .B (_2132_), .Y (n_205));
NOR2X1 g62736(.A (WX9910), .B (_2320_), .Y (n_204));
INVX2 g63273(.A (n_6510), .Y (n_972));
NOR2X1 g62732(.A (WX3477), .B (_2172_), .Y (n_201));
CLKBUFX1 g63401(.A (n_471), .Y (n_823));
NOR2X1 g62730(.A (WX6059), .B (_2210_), .Y (n_200));
NOR2X1 g62268(.A (WX4744), .B (_2189_), .Y (n_199));
NOR2X1 g62728(.A (WX4768), .B (_2177_), .Y (n_198));
NOR2X1 g62722(.A (WX8619), .B (_2287_), .Y (n_197));
NOR2X1 g62716(.A (WX7316), .B (_2260_), .Y (n_195));
NOR2X1 g62713(.A (WX11217), .B (_2345_), .Y (n_194));
NOR2X1 g61756(.A (WX9898), .B (_2326_), .Y (n_193));
NOR2X1 g62249(.A (WX4754), .B (_2184_), .Y (n_192));
NOR2X1 g62708(.A (WX7336), .B (_2250_), .Y (n_191));
NOR2X1 g62706(.A (WX4724), .B (_2199_), .Y (n_190));
NOR2X1 g61557(.A (WX4742), .B (_2190_), .Y (n_189));
NOR2X1 g61993(.A (WX8625), .B (_2300_), .Y (n_188));
NOR2X1 g62235(.A (WX8629), .B (_2282_), .Y (n_187));
NOR2X1 g62694(.A (WX7364), .B (_2268_), .Y (n_186));
NOR2X1 g62228(.A (WX2172), .B (_2118_), .Y (n_185));
NOR2X1 g62696(.A (WX4776), .B (_2173_), .Y (n_184));
NOR2X1 g62697(.A (WX2168), .B (_2120_), .Y (n_183));
NOR2X1 g61738(.A (WX8631), .B (_2281_), .Y (n_181));
NOR2X1 g62692(.A (WX7356), .B (_2268_), .Y (n_180));
NOR2X1 g62688(.A (WX4740), .B (_2191_), .Y (n_179));
NOR2X1 g62666(.A (WX6061), .B (_2209_), .Y (n_178));
NOR2X1 g62220(.A (WX7360), .B (_2238_), .Y (n_177));
NOR2X1 g61734(.A (WX3425), .B (_2170_), .Y (n_176));
NOR2X1 g62276(.A (WX3455), .B (_2155_), .Y (n_175));
NOR2X1 g62213(.A (WX11205), .B (_2351_), .Y (n_174));
NOR2X1 g62683(.A (WX4738), .B (_2192_), .Y (n_173));
NOR2X1 g61779(.A (WX6051), .B (_2214_), .Y (n_172));
NOR2X1 g61723(.A (WX3485), .B (_2172_), .Y (n_171));
NOR2X1 g62673(.A (WX3447), .B (_2159_), .Y (n_170));
NOR2X1 g61718(.A (WX4770), .B (_2204_), .Y (n_169));
NOR2X1 g62199(.A (WX11185), .B (_2361_), .Y (n_168));
NOR2X1 g61715(.A (WX7334), .B (_2251_), .Y (n_167));
NOR2X1 g62668(.A (WX6009), .B (_2235_), .Y (n_166));
NOR2X1 g61652(.A (WX7312), .B (_2262_), .Y (n_165));
NOR2X1 g61999(.A (WX6033), .B (_2223_), .Y (n_164));
NOR2X1 g62724(.A (WX4758), .B (_2182_), .Y (n_163));
NOR2X1 g62174(.A (WX4718), .B (_2202_), .Y (n_162));
NOR2X1 g62652(.A (WX2192), .B (_2140_), .Y (n_161));
NOR2X1 g62648(.A (WX11209), .B (_2349_), .Y (n_160));
NOR2X1 g62171(.A (WX7314), .B (_2261_), .Y (n_159));
NOR2X1 g62645(.A (WX11243), .B (_2364_), .Y (n_158));
NOR2X1 g62639(.A (WX7340), .B (_2248_), .Y (n_157));
NOR2X1 g62163(.A (WX6021), .B (_2229_), .Y (n_156));
NOR2X1 g61692(.A (WX3467), .B (_2149_), .Y (n_155));
NOR2X1 g62546(.A (WX4748), .B (_2187_), .Y (n_154));
NOR2X1 g61685(.A (WX11241), .B (_2333_), .Y (n_153));
NOR2X1 g61677(.A (WX2188), .B (_2110_), .Y (n_152));
NOR2X1 g61678(.A (WX11203), .B (_2352_), .Y (n_151));
NOR2X1 g61665(.A (WX7342), .B (_2268_), .Y (n_150));
NOR2X1 g61660(.A (WX2182), .B (_2113_), .Y (n_149));
NOR2X1 g62142(.A (WX7326), .B (_2255_), .Y (n_148));
NOR2X1 g61657(.A (WX8601), .B (_2296_), .Y (n_147));
INVX2 g63655(.A (n_7480), .Y (n_979));
NOR2X1 g62139(.A (WX8653), .B (_2270_), .Y (n_146));
INVX4 g63656(.A (n_7480), .Y (n_1000));
NOR2X1 g62619(.A (WX4766), .B (_2178_), .Y (n_145));
NOR2X1 g61646(.A (WX11191), .B (_2358_), .Y (n_144));
NOR2X1 g61643(.A (WX11237), .B (_2335_), .Y (n_143));
NOR2X1 g62628(.A (WX4764), .B (_2179_), .Y (n_142));
NOR2X1 g62123(.A (WX4762), .B (_2180_), .Y (n_141));
INVX4 g63238(.A (n_6622), .Y (n_943));
NOR2X1 g61628(.A (WX6019), .B (_2230_), .Y (n_137));
NOR2X1 g61622(.A (WX2138), .B (_2135_), .Y (n_136));
NOR2X1 g61614(.A (WX9900), .B (_2325_), .Y (n_135));
NOR2X1 g62616(.A (WX6013), .B (_2233_), .Y (n_133));
NOR2X1 g61604(.A (WX9940), .B (_2305_), .Y (n_131));
INVX1 g62887(.A (WX1940), .Y (n_1335));
INVX1 g62969(.A (WX821), .Y (n_130));
INVX1 g62946(.A (WX833), .Y (n_129));
INVX1 g63302(.A (WX845), .Y (n_308));
INVX1 g62856(.A (WX691), .Y (n_995));
INVX1 g62982(.A (WX1980), .Y (n_1288));
INVX1 g62817(.A (WX861), .Y (n_244));
INVX1 g62811(.A (WX863), .Y (n_438));
INVX1 g63579(.A (RESET), .Y (n_127));
INVX1 g62797(.A (WX899), .Y (n_480));
INVX1 g62845(.A (WX835), .Y (n_126));
INVX1 g63294(.A (WX677), .Y (n_938));
INVX1 g62824(.A (_2363_), .Y (n_124));
INVX1 g62967(.A (WX671), .Y (n_992));
INVX1 g62828(.A (WX1960), .Y (n_1320));
INVX1 g63297(.A (WX853), .Y (n_264));
INVX1 g62926(.A (WX659), .Y (n_940));
INVX2 g63049(.A (TM0), .Y (n_456));
INVX1 g62980(.A (WX1992), .Y (n_1437));
INVX1 g63002(.A (WX771), .Y (n_120));
INVX1 g62818(.A (WX699), .Y (n_973));
INVX1 g62771(.A (WX1952), .Y (n_1341));
INVX1 g63305(.A (WX807), .Y (n_119));
INVX1 g62833(.A (WX805), .Y (n_118));
INVX1 g63670(.A (WX803), .Y (n_117));
INVX1 g62908(.A (WX855), .Y (n_434));
INVX1 g62772(.A (WX765), .Y (n_113));
INVX1 g62829(.A (WX763), .Y (n_112));
INVX1 g62837(.A (WX759), .Y (n_111));
INVX1 g62800(.A (WX1950), .Y (n_1284));
INVX1 g62939(.A (WX731), .Y (n_109));
INVX1 g62949(.A (_2139_), .Y (n_108));
INVX1 g62985(.A (WX891), .Y (n_448));
INVX1 g63282(.A (WX1958), .Y (n_1419));
INVX1 g62974(.A (WX749), .Y (n_106));
INVX1 g62914(.A (WX723), .Y (n_105));
INVX1 g62891(.A (WX703), .Y (n_956));
INVX1 g62783(.A (WX725), .Y (n_104));
INVX1 g62781(.A (WX2000), .Y (n_2675));
INVX1 g63280(.A (WX729), .Y (n_101));
INVX1 g62954(.A (WX751), .Y (n_100));
INVX1 g63674(.A (WX1968), .Y (n_2825));
INVX1 g62894(.A (WX785), .Y (n_98));
INVX1 g62794(.A (WX839), .Y (n_276));
INVX1 g62857(.A (WX819), .Y (n_96));
INVX1 g60143(.A (WX709), .Y (n_95));
INVX1 g62938(.A (WX679), .Y (n_932));
INVX1 g62995(.A (WX897), .Y (n_443));
INVX1 g62973(.A (WX867), .Y (n_476));
INVX1 g62924(.A (WX705), .Y (n_951));
INVX1 g62879(.A (WX797), .Y (n_89));
INVX1 g63275(.A (WX1998), .Y (n_1451));
INVX1 g63307(.A (WX1944), .Y (n_1339));
INVX1 g62902(.A (WX665), .Y (n_953));
INVX1 g63308(.A (WX675), .Y (n_948));
INVX1 g62779(.A (WX895), .Y (n_278));
INVX1 g62978(.A (WX769), .Y (n_87));
INVX1 g62996(.A (WX767), .Y (n_85));
INVX1 g63298(.A (WX775), .Y (n_83));
INVX1 g62883(.A (WX673), .Y (n_987));
INVX1 g62898(.A (WX777), .Y (n_81));
INVX1 g62776(.A (WX859), .Y (n_280));
INVX1 g62780(.A (WX651), .Y (n_927));
INVX1 g62862(.A (WX663), .Y (n_920));
INVX1 g62847(.A (WX795), .Y (n_79));
INVX1 g62890(.A (WX847), .Y (n_252));
INVX1 g62945(.A (WX875), .Y (n_429));
INVX1 g62803(.A (WX1974), .Y (n_1348));
INVX1 g62988(.A (WX815), .Y (n_73));
INVX1 g62855(.A (WX647), .Y (n_997));
INVX1 g63293(.A (WX881), .Y (n_261));
INVX1 g62918(.A (WX715), .Y (n_71));
INVX1 g63675(.A (WX817), .Y (n_70));
INVX2 g63010(.A (TM0), .Y (n_450));
INVX1 g63279(.A (WX653), .Y (n_990));
INVX1 g62998(.A (WX1984), .Y (n_1282));
INVX1 g62962(.A (WX869), .Y (n_474));
INVX1 g62966(.A (WX1994), .Y (n_1429));
INVX1 g63303(.A (WX823), .Y (n_69));
INVX1 g62941(.A (WX829), .Y (n_68));
INVX1 g62897(.A (WX1982), .Y (n_1309));
INVX1 g62814(.A (WX701), .Y (n_962));
INVX1 g62788(.A (WX757), .Y (n_67));
INVX1 g62948(.A (WX655), .Y (n_905));
INVX1 g63311(.A (WX683), .Y (n_964));
INVX1 g62957(.A (WX1972), .Y (n_1431));
INVX1 g62968(.A (WX1942), .Y (n_1359));
INVX1 g62922(.A (WX711), .Y (n_65));
INVX1 g62808(.A (WX885), .Y (n_482));
INVX1 g63276(.A (WX713), .Y (n_63));
INVX1 g62896(.A (WX649), .Y (n_929));
INVX1 g62905(.A (WX865), .Y (n_462));
INVX1 g62882(.A (WX1964), .Y (n_1323));
INVX1 g62956(.A (WX1986), .Y (n_2691));
INVX1 g62901(.A (WX645), .Y (n_1006));
INVX1 g62839(.A (WX697), .Y (n_970));
INVX1 g62990(.A (WX667), .Y (n_1001));
BUFX3 g63456(.A (RESET), .Y (n_471));
INVX1 g62886(.A (WX873), .Y (n_486));
INVX1 g62892(.A (WX1954), .Y (n_1449));
INVX1 g62936(.A (WX827), .Y (n_58));
INVX1 g62927(.A (WX1966), .Y (n_1427));
CLKBUFX3 g63578(.A (RESET), .Y (n_1297));
INVX1 g62854(.A (WX689), .Y (n_1004));
INVX1 g63001(.A (WX893), .Y (n_451));
INVX1 g62881(.A (WX1988), .Y (n_1442));
INVX1 g62909(.A (WX787), .Y (n_56));
INVX1 g62866(.A (WX687), .Y (n_958));
INVX1 g62931(.A (WX727), .Y (n_52));
INVX1 g62878(.A (WX695), .Y (n_975));
INVX1 g62769(.A (WX733), .Y (n_51));
INVX1 g62925(.A (WX1956), .Y (n_1421));
INVX1 g62953(.A (WX851), .Y (n_454));
INVX1 g63289(.A (WX813), .Y (n_49));
INVX1 g62831(.A (WX737), .Y (n_48));
INVX1 g62798(.A (WX739), .Y (n_46));
INVX1 g62920(.A (WX745), .Y (n_44));
INVX1 g63006(.A (WX747), .Y (n_43));
INVX1 g62930(.A (WX843), .Y (n_436));
INVX1 g62900(.A (blif_reset_net), .Y (n_6171));
INVX1 g62827(.A (WX841), .Y (n_273));
INVX1 g62782(.A (WX1978), .Y (n_1374));
INVX1 g63679(.A (WX779), .Y (n_41));
INVX1 g62801(.A (WX781), .Y (n_40));
INVX1 g62790(.A (WX793), .Y (n_38));
INVX1 g62819(.A (WX799), .Y (n_36));
INVX1 g62785(.A (WX791), .Y (n_35));
INVX1 g62958(.A (WX809), .Y (n_33));
INVX1 g62981(.A (WX661), .Y (n_935));
INVX1 g62852(.A (WX761), .Y (n_32));
INVX1 g62836(.A (WX485), .Y (n_3599));
INVX1 g62844(.A (WX883), .Y (n_484));
INVX1 g63004(.A (WX801), .Y (n_28));
INVX1 g63309(.A (WX789), .Y (n_27));
INVX1 g62863(.A (WX783), .Y (n_24));
INVX1 g62965(.A (WX849), .Y (n_420));
INVX1 g62851(.A (WX877), .Y (n_271));
INVX1 g62787(.A (WX693), .Y (n_985));
INVX1 g62867(.A (WX811), .Y (n_21));
INVX1 g62986(.A (WX741), .Y (n_20));
INVX1 g62935(.A (WX879), .Y (n_431));
INVX1 g62822(.A (WX755), .Y (n_19));
INVX1 g63286(.A (WX753), .Y (n_18));
INVX1 g62917(.A (WX1962), .Y (n_1345));
INVX1 g62976(.A (WX743), .Y (n_16));
INVX1 g62872(.A (WX707), .Y (n_944));
INVX1 g62870(.A (WX735), .Y (n_14));
INVX1 g62950(.A (WX1990), .Y (n_1328));
INVX1 g63278(.A (WX1970), .Y (n_1350));
INVX1 g62821(.A (WX685), .Y (n_913));
INVX1 g62913(.A (WX857), .Y (n_354));
INVX1 g62812(.A (WX721), .Y (n_12));
INVX1 g62869(.A (WX669), .Y (n_981));
INVX1 g58184(.A (WX837), .Y (n_139));
INVX1 g63678(.A (WX657), .Y (n_977));
INVX1 g62873(.A (WX1946), .Y (n_1412));
INVX1 g63288(.A (WX1996), .Y (n_1318));
INVX1 g62877(.A (WX1976), .Y (n_1286));
INVX1 g63285(.A (WX871), .Y (n_283));
INVX1 g62893(.A (WX1948), .Y (n_1357));
INVX1 g62916(.A (WX681), .Y (n_924));
INVX1 g62840(.A (WX831), .Y (n_5));
INVX1 g62804(.A (WX719), .Y (n_4));
INVX1 g62865(.A (WX10989), .Y (n_1315));
INVX1 g62876(.A (WX887), .Y (n_266));
INVX1 g55946(.A (WX489), .Y (n_3685));
INVX1 g63672(.A (WX825), .Y (n_3));
INVX1 g62991(.A (WX717), .Y (n_2));
INVX1 g62861(.A (WX889), .Y (n_268));
INVX1 g63677(.A (WX1938), .Y (n_1337));
INVX1 g58623(.A (WX773), .Y (n_0));
XOR2X1 g24(.A (WX3319), .B (n_6424), .Y (n_6425));
XOR2X1 g25(.A (WX3255), .B (n_6423), .Y (n_6424));
INVX1 g29(.A (n_6422), .Y (n_6423));
INVX2 g30(.A (n_7487), .Y (n_6422));
CLKBUFX1 g26(.A (n_7487), .Y (n_6428));
INVX1 g27(.A (n_7487), .Y (n_6429));
INVX2 g3(.A (n_6430), .Y (n_6431));
INVX2 g4(.A (TM1), .Y (n_6430));
INVX4 g1(.A (n_6430), .Y (n_6432));
INVX2 g2(.A (n_6430), .Y (n_6433));
NOR2X1 g14(.A (n_6438), .B (WX10845), .Y (n_6439));
INVX1 g65498(.A (n_6437), .Y (n_6438));
INVX4 g65499(.A (n_6624), .Y (n_6437));
NOR3X1 g65504(.A (n_6446), .B (n_6449), .C (n_6450), .Y (n_6451));
INVX2 g46(.A (n_6624), .Y (n_6446));
NOR2X1 g65505(.A (n_6447), .B (n_6448), .Y (n_6449));
XOR2X1 g65506(.A (WX7240), .B (WX7304), .Y (n_6447));
XOR2X1 g65507(.A (WX7176), .B (n_3034), .Y (n_6448));
AND2X1 g65508(.A (n_6448), .B (n_6447), .Y (n_6450));
INVX4 g43(.A (n_6446), .Y (n_6452));
OAI21X1 g40(.A0 (n_6458), .A1 (n_3426), .B0 (n_6466), .Y (n_6467));
INVX1 g42(.A (n_6457), .Y (n_6458));
NAND2X1 g65509(.A (n_6455), .B (n_6456), .Y (n_6457));
NAND2X1 g52(.A (n_3222), .B (n_6454), .Y (n_6455));
INVX1 g57(.A (WX10865), .Y (n_6454));
NAND2X1 g46_dup(.A (n_4100), .B (n_3737), .Y (n_6456));
OR2X1 g41(.A (n_5535), .B (n_6465), .Y (n_6466));
AOI22X1 g44(.A0 (_2346_), .A1 (n_3835), .B0 (n_4670), .B1(DATA_0_13), .Y (n_6465));
INVX1 g45(.A (n_6468), .Y (n_6469));
NAND2X1 g65511(.A (n_4100), .B (n_3737), .Y (n_6468));
OAI21X1 g36(.A0 (n_6475), .A1 (n_6480), .B0 (n_6485), .Y (n_6486));
INVX1 g38(.A (n_6474), .Y (n_6475));
NAND2X1 g39(.A (n_6472), .B (n_6473), .Y (n_6474));
NAND2X1 g65512(.A (n_3225), .B (n_6471), .Y (n_6472));
INVX1 g54(.A (WX10875), .Y (n_6471));
NAND2X1 g42_dup(.A (n_4094), .B (n_3894), .Y (n_6473));
INVX1 g65514(.A (n_6479), .Y (n_6480));
CLKBUFX1 g65515(.A (n_6497), .Y (n_6479));
OR2X1 g37(.A (n_5439), .B (n_6484), .Y (n_6485));
CLKBUFX3 g65520(.A (n_7089), .Y (n_6482));
AOI22X1 g65522(.A0 (_2341_), .A1 (n_5873), .B0 (n_3828), .B1(DATA_0_8), .Y (n_6484));
INVX1 g65523(.A (n_6487), .Y (n_6488));
NAND2X1 g65524(.A (n_4094), .B (n_3894), .Y (n_6487));
OAI21X1 g35(.A0 (n_6495), .A1 (n_6480), .B0 (n_6504), .Y (n_6505));
INVX1 g65526(.A (n_6494), .Y (n_6495));
NAND2X1 g65527(.A (n_6492), .B (n_6493), .Y (n_6494));
NAND2X1 g65528(.A (n_3223), .B (n_6491), .Y (n_6492));
INVX1 g65530(.A (WX9542), .Y (n_6491));
NAND2X1 g41_dup(.A (n_4101), .B (n_4000), .Y (n_6493));
CLKBUFX3 g65534(.A (n_7086), .Y (n_6497));
OAI21X1 g65536(.A0 (n_4549), .A1 (n_6501), .B0 (n_6503), .Y (n_6504));
AND2X1 g65537(.A (n_4586), .B (_2329_), .Y (n_6501));
CLKBUFX3 g51(.A (n_7089), .Y (n_6503));
INVX1 g65540(.A (n_6507), .Y (n_6508));
NAND2X1 g65541(.A (n_4101), .B (n_4000), .Y (n_6507));
XOR2X1 g21(.A (WX7216), .B (n_6514), .Y (n_6515));
XOR2X1 g22(.A (WX7152), .B (n_6513), .Y (n_6514));
INVX2 g65543(.A (n_6512), .Y (n_6513));
INVX4 g65544(.A (n_6511), .Y (n_6512));
INVX2 g65545(.A (n_6510), .Y (n_6511));
INVX2 g65546(.A (TM0), .Y (n_6510));
NAND2X2 g19(.A (n_6520), .B (n_6523), .Y (n_6524));
NAND2X2 g20(.A (n_6555), .B (n_6519), .Y (n_6520));
OAI21X1 g65549(.A0 (n_5944), .A1 (n_5889), .B0 (n_5898), .Y (n_6519));
NAND2X1 g65550(.A (n_6521), .B (n_2922), .Y (n_6523));
INVX1 g65551(.A (n_4165), .Y (n_6521));
NAND2X2 g65554(.A (n_6529), .B (n_6532), .Y (n_6533));
NAND2X2 g65555(.A (n_6575), .B (n_6528), .Y (n_6529));
OAI21X1 g65557(.A0 (n_5727), .A1 (n_5889), .B0 (n_5671), .Y (n_6528));
NAND2X2 g65558(.A (n_6530), .B (n_2922), .Y (n_6532));
INVX1 g65559(.A (n_4157), .Y (n_6530));
NAND2X2 g65561(.A (n_6537), .B (n_6540), .Y (n_6541));
NAND2X2 g65562(.A (n_6575), .B (n_6536), .Y (n_6537));
OAI21X1 g65565(.A0 (n_5543), .A1 (n_5889), .B0 (n_5445), .Y (n_6536));
NAND2X2 g65566(.A (n_6538), .B (n_2922), .Y (n_6540));
INVX1 g65567(.A (n_4151), .Y (n_6538));
NAND2X2 g65569(.A (n_6545), .B (n_6548), .Y (n_6549));
NAND2X2 g65570(.A (n_6583), .B (n_6544), .Y (n_6545));
OAI21X1 g65572(.A0 (n_5164), .A1 (n_5889), .B0 (n_5065), .Y (n_6544));
NAND2X2 g65573(.A (n_6546), .B (n_2922), .Y (n_6548));
INVX1 g65574(.A (n_4142), .Y (n_6546));
MX2X1 g65576(.A (n_6551), .B (n_6550), .S0 (n_6552), .Y (n_6553));
INVX1 g65577(.A (n_6550), .Y (n_6551));
NAND2X1 g65578(.A (n_541), .B (n_539), .Y (n_6550));
MX2X1 g65579(.A (n_101), .B (WX729), .S0 (n_2421), .Y (n_6552));
NAND2X2 g65580(.A (n_6557), .B (n_6560), .Y (n_6561));
NAND2X2 g65581(.A (n_6555), .B (n_6556), .Y (n_6557));
CLKBUFX3 g65582(.A (n_6614), .Y (n_6555));
OAI21X1 g65584(.A0 (n_5903), .A1 (n_5889), .B0 (n_5848), .Y (n_6556));
NAND2X1 g65585(.A (n_6558), .B (n_2922), .Y (n_6560));
INVX1 g65586(.A (n_4163), .Y (n_6558));
MX2X1 g65595(.A (n_6571), .B (n_6570), .S0 (n_6572), .Y (n_6573));
INVX1 g65596(.A (n_6570), .Y (n_6571));
NAND2X1 g65597(.A (n_558), .B (n_556), .Y (n_6570));
MX2X1 g65598(.A (n_44), .B (WX745), .S0 (n_2440), .Y (n_6572));
NAND2X2 g65599(.A (n_6577), .B (n_6580), .Y (n_6581));
NAND2X2 g65600(.A (n_6575), .B (n_6576), .Y (n_6577));
CLKBUFX3 g65601(.A (n_6614), .Y (n_6575));
OAI21X1 g65602(.A0 (n_5612), .A1 (n_5889), .B0 (n_5539), .Y (n_6576));
NAND2X1 g65603(.A (n_6578), .B (n_6619), .Y (n_6580));
INVX1 g65604(.A (n_4153), .Y (n_6578));
NAND2X2 g65606(.A (n_6585), .B (n_6588), .Y (n_6589));
NAND2X2 g65607(.A (n_6583), .B (n_6584), .Y (n_6585));
CLKBUFX3 g65608(.A (n_6614), .Y (n_6583));
OAI21X1 g65610(.A0 (n_5450), .A1 (n_5889), .B0 (n_5355), .Y (n_6584));
NAND2X1 g65611(.A (n_6586), .B (n_6619), .Y (n_6588));
INVX1 g65612(.A (n_4148), .Y (n_6586));
MX2X1 g65621(.A (n_6599), .B (n_6598), .S0 (n_6600), .Y (n_6601));
INVX1 g65622(.A (n_6598), .Y (n_6599));
NAND2X1 g65623(.A (n_587), .B (n_595), .Y (n_6598));
MX2X1 g65624(.A (n_111), .B (WX759), .S0 (n_2488), .Y (n_6600));
MX2X1 g65632(.A (n_6611), .B (n_6610), .S0 (n_6612), .Y (n_6613));
INVX1 g65633(.A (n_6610), .Y (n_6611));
NAND2X1 g65634(.A (n_585), .B (n_574), .Y (n_6610));
MX2X1 g65635(.A (n_113), .B (WX765), .S0 (n_2434), .Y (n_6612));
NAND2X2 g65636(.A (n_6617), .B (n_6620), .Y (n_6621));
NAND2X2 g65637(.A (n_6615), .B (n_6616), .Y (n_6617));
CLKBUFX2 g65638(.A (n_6614), .Y (n_6615));
AND2X1 g23(.A (n_3140), .B (RESET), .Y (n_6614));
OAI21X1 g65639(.A0 (n_4863), .A1 (n_5889), .B0 (n_4655), .Y (n_6616));
NAND2X1 g65640(.A (n_6618), .B (n_6619), .Y (n_6620));
INVX1 g65641(.A (n_4136), .Y (n_6618));
INVX1 g65642(.A (n_4697), .Y (n_6619));
NOR3X1 g65643(.A (n_5873), .B (n_6630), .C (n_6631), .Y (n_6632));
INVX4 g65645(.A (n_6437), .Y (n_6626));
CLKBUFX3 g65647(.A (n_6623), .Y (n_6624));
CLKBUFX3 g65648(.A (n_6622), .Y (n_6623));
INVX2 g65649(.A (TM0), .Y (n_6622));
NOR2X1 g65650(.A (n_6628), .B (n_6629), .Y (n_6630));
XOR2X1 g65651(.A (WX4676), .B (WX4740), .Y (n_6628));
XOR2X1 g65652(.A (WX4612), .B (n_3149), .Y (n_6629));
AND2X1 g65653(.A (n_6629), .B (n_6628), .Y (n_6631));
INVX4 g65654(.A (n_5873), .Y (n_6633));
MX2X1 g65663(.A (n_6643), .B (n_6642), .S0 (n_6644), .Y (n_6645));
INVX1 g65664(.A (n_6642), .Y (n_6643));
NAND2X1 g65665(.A (n_589), .B (n_592), .Y (n_6642));
MX2X1 g65666(.A (n_109), .B (WX731), .S0 (n_2508), .Y (n_6644));
AND2X1 g65763(.A (n_4099), .B (n_6884), .Y (n_6885));
AND2X1 g58048_dup(.A (n_4099), .B (n_6884), .Y (n_6886));
MX2X1 g65840(.A (n_7060), .B (n_7059), .S0 (n_7061), .Y (n_7062));
INVX1 g65841(.A (n_7059), .Y (n_7060));
NAND2X1 g65842(.A (n_562), .B (n_560), .Y (n_7059));
MX2X1 g65843(.A (n_104), .B (WX725), .S0 (n_2457), .Y (n_7061));
MX2X1 g65844(.A (n_7064), .B (n_7063), .S0 (n_7065), .Y (n_7066));
INVX1 g65845(.A (n_7063), .Y (n_7064));
NAND2X1 g65846(.A (n_588), .B (n_594), .Y (n_7063));
MX2X1 g65847(.A (n_4), .B (WX719), .S0 (n_2409), .Y (n_7065));
MX2X1 g65848(.A (n_7068), .B (n_7067), .S0 (n_7069), .Y (n_7070));
INVX1 g65849(.A (n_7067), .Y (n_7068));
NAND2X1 g65850(.A (n_554), .B (n_553), .Y (n_7067));
MX2X1 g65851(.A (n_52), .B (WX727), .S0 (n_2439), .Y (n_7069));
MX2X1 g65852(.A (n_7072), .B (n_7071), .S0 (n_7073), .Y (n_7074));
INVX1 g65853(.A (n_7071), .Y (n_7072));
NAND2X1 g65854(.A (n_581), .B (n_524), .Y (n_7071));
MX2X1 g65855(.A (n_14), .B (WX735), .S0 (n_2419), .Y (n_7073));
MX2X1 g65856(.A (n_7076), .B (n_7075), .S0 (n_7077), .Y (n_7078));
INVX1 g65857(.A (n_7075), .Y (n_7076));
NAND2X1 g65858(.A (n_546), .B (n_586), .Y (n_7075));
MX2X1 g65859(.A (n_46), .B (WX739), .S0 (n_2481), .Y (n_7077));
MX2X1 g65860(.A (n_7080), .B (n_7079), .S0 (n_7081), .Y (n_7082));
INVX1 g65861(.A (n_7079), .Y (n_7080));
NAND2X1 g65862(.A (n_575), .B (n_577), .Y (n_7079));
MX2X1 g65863(.A (n_63), .B (WX713), .S0 (n_2431), .Y (n_7081));
OAI21X1 g65864(.A0 (n_7085), .A1 (n_7088), .B0 (n_7093), .Y (n_7094));
NOR2X1 g65865(.A (n_7083), .B (n_7084), .Y (n_7085));
NOR2X1 g65866(.A (WX10861), .B (n_5427), .Y (n_7083));
AND2X1 g65867(.A (n_3741), .B (n_6633), .Y (n_7084));
INVX8 g65868(.A (n_7087), .Y (n_7088));
CLKBUFX3 g65869(.A (n_7086), .Y (n_7087));
AND2X1 g65870(.A (RESET), .B (n_3140), .Y (n_7086));
OR2X1 g65871(.A (n_5841), .B (n_7092), .Y (n_7093));
CLKBUFX3 g49(.A (n_7089), .Y (n_7090));
NOR2X1 g50(.A (n_3140), .B (n_127), .Y (n_7089));
AOI22X1 g65872(.A0 (_2348_), .A1 (n_3835), .B0 (n_5968), .B1(DATA_0_15), .Y (n_7092));
XOR2X1 g66050(.A (WX8467), .B (n_7484), .Y (n_7485));
XOR2X1 g66051(.A (WX8403), .B (n_7483), .Y (n_7484));
INVX2 g66052(.A (n_7482), .Y (n_7483));
INVX4 g66053(.A (n_7481), .Y (n_7482));
INVX2 g66054(.A (n_7480), .Y (n_7481));
INVX4 g33(.A (TM1), .Y (n_7480));
INVX4 g66056(.A (n_7480), .Y (n_7487));
INVX1 g66057(.A (n_7483), .Y (n_7488));
INVX4 g66059(.A (n_7480), .Y (n_7490));
AND2X1 g66953(.A (n_4017), .B (n_8314), .Y (n_9404));
AND2X1 g57917_dup(.A (n_4017), .B (n_8314), .Y (n_9405));
AND2X1 g66954(.A (n_4101), .B (n_8315), .Y (n_9406));
AND2X1 g58144_dup(.A (n_4101), .B (n_8315), .Y (n_9407));
AND2X1 g66955(.A (n_4099), .B (n_8316), .Y (n_9408));
AND2X1 g57947_dup(.A (n_4099), .B (n_8316), .Y (n_9409));
AND2X1 g66956(.A (n_4096), .B (n_8317), .Y (n_9410));
AND2X1 g57919_dup(.A (n_4096), .B (n_8317), .Y (n_9411));
AND2X1 g66957(.A (n_4017), .B (n_8318), .Y (n_9412));
AND2X1 g57941_dup(.A (n_4017), .B (n_8318), .Y (n_9413));
AND2X1 g66958(.A (n_4100), .B (n_8319), .Y (n_9414));
AND2X1 g58090_dup(.A (n_4100), .B (n_8319), .Y (n_9415));
AND2X1 g66959(.A (n_4106), .B (n_8321), .Y (n_9416));
AND2X1 g57967_dup(.A (n_4106), .B (n_8321), .Y (n_15867));
AND2X1 g66960(.A (n_4105), .B (n_8323), .Y (n_9418));
AND2X1 g57911_dup(.A (n_4105), .B (n_8323), .Y (n_9419));
AND2X1 g66961(.A (n_4103), .B (n_8324), .Y (n_9420));
AND2X1 g58008_dup(.A (n_4103), .B (n_8324), .Y (n_9421));
AND2X1 g66962(.A (n_6633), .B (n_8325), .Y (n_9422));
AND2X1 g58077_dup(.A (n_6633), .B (n_8325), .Y (n_9423));
CLKBUFX2 g66963(.A (n_6511), .Y (n_9424));
CLKBUFX1 g65547_dup(.A (n_6511), .Y (n_9425));
AND2X1 g66964(.A (n_4101), .B (n_8326), .Y (n_9426));
AND2X1 g58016_dup(.A (n_4101), .B (n_8326), .Y (n_9427));
AND2X1 g66965(.A (n_4103), .B (n_8327), .Y (n_9428));
AND2X1 g58150_dup(.A (n_4103), .B (n_8327), .Y (n_9429));
MX2X1 g66966(.A (n_9431), .B (n_9430), .S0 (n_9432), .Y (n_9433));
INVX1 g66967(.A (n_9430), .Y (n_9431));
NAND2X1 g66968(.A (n_817), .B (n_830), .Y (n_9430));
MX2X1 g66969(.A (n_95), .B (WX709), .S0 (n_2425), .Y (n_9432));
MX2X1 g66970(.A (n_9435), .B (n_9434), .S0 (n_9436), .Y (n_9437));
INVX1 g66971(.A (n_9434), .Y (n_9435));
NAND2X1 g66972(.A (n_572), .B (n_550), .Y (n_9434));
MX2X1 g66973(.A (n_120), .B (WX771), .S0 (n_2465), .Y (n_9436));
MX2X1 g67130(.A (n_9798), .B (n_9797), .S0 (n_9799), .Y (n_9800));
INVX1 g67131(.A (n_9797), .Y (n_9798));
NAND2X1 g67132(.A (n_591), .B (n_571), .Y (n_9797));
MX2X1 g67133(.A (n_48), .B (WX737), .S0 (n_2503), .Y (n_9799));
AND2X1 g67587(.A (n_4100), .B (n_8350), .Y (n_10712));
AND2X1 g58158_dup(.A (n_4100), .B (n_8350), .Y (n_10713));
AND2X1 g67588(.A (n_4095), .B (n_8351), .Y (n_10714));
AND2X1 g58100_dup(.A (n_4095), .B (n_8351), .Y (n_15863));
AND2X1 g67589(.A (n_4095), .B (n_8352), .Y (n_10716));
AND2X1 g58029_dup(.A (n_4095), .B (n_8352), .Y (n_10717));
AND2X1 g67590(.A (n_4106), .B (n_8353), .Y (n_10718));
AND2X1 g58099_dup(.A (n_4106), .B (n_8353), .Y (n_10719));
AND2X1 g67591(.A (n_6452), .B (n_8354), .Y (n_10720));
AND2X1 g58112_dup(.A (n_6452), .B (n_8354), .Y (n_10721));
AND2X1 g67592(.A (n_4104), .B (n_8355), .Y (n_10722));
AND2X1 g58036_dup(.A (n_4104), .B (n_8355), .Y (n_10723));
MX2X1 g67593(.A (n_10725), .B (n_10724), .S0 (n_10726), .Y (n_10727));
INVX1 g67594(.A (n_10724), .Y (n_10725));
NAND2X1 g67595(.A (n_565), .B (n_542), .Y (n_10724));
MX2X1 g67596(.A (n_105), .B (WX723), .S0 (n_2493), .Y (n_10726));
MX2X1 g67597(.A (n_10729), .B (n_10728), .S0 (n_10730), .Y (n_10731));
INVX1 g67598(.A (n_10728), .Y (n_10729));
NAND2X1 g67599(.A (n_561), .B (n_579), .Y (n_10728));
MX2X1 g67600(.A (n_51), .B (WX733), .S0 (n_2497), .Y (n_10730));
MX2X1 g67601(.A (n_10733), .B (n_10732), .S0 (n_10734), .Y (n_10735));
INVX1 g67602(.A (n_10732), .Y (n_10733));
NAND2X1 g67603(.A (n_552), .B (n_549), .Y (n_10732));
MX2X1 g67604(.A (n_43), .B (WX747), .S0 (n_2428), .Y (n_10734));
MX2X1 g67605(.A (n_10737), .B (n_10736), .S0 (n_10738), .Y (n_10739));
INVX1 g67606(.A (n_10736), .Y (n_10737));
NAND2X1 g67607(.A (n_540), .B (n_543), .Y (n_10736));
MX2X1 g67608(.A (n_100), .B (WX751), .S0 (n_2412), .Y (n_10738));
MX2X1 g67609(.A (n_10741), .B (n_10740), .S0 (n_10742), .Y (n_10743));
INVX1 g67610(.A (n_10740), .Y (n_10741));
NAND2X1 g67611(.A (n_584), .B (n_580), .Y (n_10740));
MX2X1 g67612(.A (n_32), .B (WX761), .S0 (n_2484), .Y (n_10742));
MX2X1 g67613(.A (n_10745), .B (n_10744), .S0 (n_10746), .Y (n_10747));
INVX1 g67614(.A (n_10744), .Y (n_10745));
NAND2X1 g67615(.A (n_523), .B (n_567), .Y (n_10744));
MX2X1 g67616(.A (n_65), .B (WX711), .S0 (n_2505), .Y (n_10746));
AND2X1 g68036(.A (n_4105), .B (n_9384), .Y (n_11595));
AND2X1 g57962_dup(.A (n_4105), .B (n_9384), .Y (n_11596));
AND2X1 g68037(.A (n_4099), .B (n_9385), .Y (n_11597));
AND2X1 g57951_dup(.A (n_4099), .B (n_9385), .Y (n_15865));
AND2X1 g68038(.A (n_4100), .B (n_9386), .Y (n_11599));
AND2X1 g58108_dup(.A (n_4100), .B (n_9386), .Y (n_11600));
AND2X1 g68039(.A (n_4094), .B (n_9387), .Y (n_11601));
AND2X1 g57968_dup(.A (n_4094), .B (n_9387), .Y (n_11602));
AND2X1 g68040(.A (n_4099), .B (n_9388), .Y (n_11603));
AND2X1 g58103_dup(.A (n_4099), .B (n_9388), .Y (n_11604));
AND2X1 g68041(.A (n_4017), .B (n_9389), .Y (n_11605));
AND2X1 g57918_dup(.A (n_4017), .B (n_9389), .Y (n_15855));
AND2X1 g68042(.A (n_6452), .B (n_9390), .Y (n_11607));
AND2X1 g58012_dup(.A (n_6452), .B (n_9390), .Y (n_11608));
AND2X1 g68043(.A (n_4094), .B (n_9391), .Y (n_11609));
AND2X1 g58146_dup(.A (n_4094), .B (n_9391), .Y (n_15857));
AND2X1 g68044(.A (n_6633), .B (n_9392), .Y (n_11611));
AND2X1 g58056_dup(.A (n_6633), .B (n_9392), .Y (n_11612));
AND2X1 g68045(.A (n_6452), .B (n_9393), .Y (n_11613));
AND2X1 g58148_dup(.A (n_6452), .B (n_9393), .Y (n_11614));
AND2X1 g68046(.A (n_4095), .B (n_9394), .Y (n_11615));
AND2X1 g58017_dup(.A (n_4095), .B (n_9394), .Y (n_11616));
AND2X1 g68047(.A (n_4096), .B (n_9395), .Y (n_11617));
AND2X1 g58088_dup(.A (n_4096), .B (n_9395), .Y (n_11618));
AND2X1 g68048(.A (n_4017), .B (n_9396), .Y (n_11619));
AND2X1 g57933_dup(.A (n_4017), .B (n_9396), .Y (n_15851));
AND2X1 g68049(.A (n_4103), .B (n_9397), .Y (n_11621));
AND2X1 g58094_dup(.A (n_4103), .B (n_9397), .Y (n_15859));
AND2X1 g68050(.A (n_4105), .B (n_9398), .Y (n_11623));
AND2X1 g57943_dup(.A (n_4105), .B (n_9398), .Y (n_15861));
AND2X1 g68051(.A (n_4094), .B (n_9399), .Y (n_11625));
AND2X1 g58096_dup(.A (n_4094), .B (n_9399), .Y (n_11626));
endmodule
